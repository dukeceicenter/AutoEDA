../macros/freepdk45_sram_1w1r_12x256/freepdk45_sram_1w1r_12x256.lef