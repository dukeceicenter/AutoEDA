VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_128x32_32
   CLASS BLOCK ;
   SIZE 147.245 BY 134.51 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.075 1.1075 24.21 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.935 1.1075 27.07 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.795 1.1075 29.93 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.655 1.1075 32.79 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.515 1.1075 35.65 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.375 1.1075 38.51 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.235 1.1075 41.37 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.095 1.1075 44.23 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.955 1.1075 47.09 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.815 1.1075 49.95 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.675 1.1075 52.81 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.535 1.1075 55.67 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.395 1.1075 58.53 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.255 1.1075 61.39 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.115 1.1075 64.25 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.975 1.1075 67.11 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.835 1.1075 69.97 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.695 1.1075 72.83 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.555 1.1075 75.69 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.415 1.1075 78.55 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.275 1.1075 81.41 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.135 1.1075 84.27 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.995 1.1075 87.13 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.855 1.1075 89.99 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.715 1.1075 92.85 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.575 1.1075 95.71 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.435 1.1075 98.57 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.295 1.1075 101.43 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.155 1.1075 104.29 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.015 1.1075 107.15 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.875 1.1075 110.01 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.735 1.1075 112.87 1.2425 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.215 1.1075 21.35 1.2425 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 45.6975 15.63 45.8325 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 48.4275 15.63 48.5625 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 50.6375 15.63 50.7725 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 53.3675 15.63 53.5025 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 55.5775 15.63 55.7125 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 58.3075 15.63 58.4425 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.895 132.0025 123.03 132.1375 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 19.5675 131.61 19.7025 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 16.8375 131.61 16.9725 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 14.6275 131.61 14.7625 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 11.8975 131.61 12.0325 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 9.6875 131.61 9.8225 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 6.9575 131.61 7.0925 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.825 133.2675 146.96 133.4025 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.7225 133.1825 140.8575 133.3175 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.8225 129.515 35.9575 129.65 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.1725 129.515 38.3075 129.65 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.5225 129.515 40.6575 129.65 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.8725 129.515 43.0075 129.65 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.2225 129.515 45.3575 129.65 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.5725 129.515 47.7075 129.65 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.9225 129.515 50.0575 129.65 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.2725 129.515 52.4075 129.65 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.6225 129.515 54.7575 129.65 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.9725 129.515 57.1075 129.65 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.3225 129.515 59.4575 129.65 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.6725 129.515 61.8075 129.65 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.0225 129.515 64.1575 129.65 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.3725 129.515 66.5075 129.65 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.7225 129.515 68.8575 129.65 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.0725 129.515 71.2075 129.65 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.4225 129.515 73.5575 129.65 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.7725 129.515 75.9075 129.65 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.1225 129.515 78.2575 129.65 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.4725 129.515 80.6075 129.65 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.8225 129.515 82.9575 129.65 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.1725 129.515 85.3075 129.65 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.5225 129.515 87.6575 129.65 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.8725 129.515 90.0075 129.65 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.2225 129.515 92.3575 129.65 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.5725 129.515 94.7075 129.65 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.9225 129.515 97.0575 129.65 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.2725 129.515 99.4075 129.65 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.6225 129.515 101.7575 129.65 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.9725 129.515 104.1075 129.65 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.3225 129.515 106.4575 129.65 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.6725 129.515 108.8075 129.65 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  125.4625 31.1375 125.5975 31.2725 ;
         LAYER metal3 ;
         RECT  32.6375 120.105 112.2975 120.175 ;
         LAYER metal3 ;
         RECT  21.3125 22.1675 21.4475 22.3025 ;
         LAYER metal3 ;
         RECT  23.7925 2.4725 23.9275 2.6075 ;
         LAYER metal3 ;
         RECT  115.2825 117.8475 115.4175 117.9825 ;
         LAYER metal3 ;
         RECT  25.575 11.9075 25.71 12.0425 ;
         LAYER metal3 ;
         RECT  46.6725 2.4725 46.8075 2.6075 ;
         LAYER metal3 ;
         RECT  119.29 117.06 119.425 117.195 ;
         LAYER metal3 ;
         RECT  125.4625 40.1075 125.5975 40.2425 ;
         LAYER metal3 ;
         RECT  21.3125 43.0975 21.4475 43.2325 ;
         LAYER metal3 ;
         RECT  92.4325 2.4725 92.5675 2.6075 ;
         LAYER metal3 ;
         RECT  103.8725 2.4725 104.0075 2.6075 ;
         LAYER metal3 ;
         RECT  58.1125 2.4725 58.2475 2.6075 ;
         LAYER metal3 ;
         RECT  125.4625 25.1575 125.5975 25.2925 ;
         LAYER metal3 ;
         RECT  121.2 124.9375 121.335 125.0725 ;
         LAYER metal3 ;
         RECT  32.6375 126.9575 109.4775 127.0275 ;
         LAYER metal4 ;
         RECT  17.93 2.47 18.07 17.43 ;
         LAYER metal4 ;
         RECT  114.2 17.5 114.34 119.41 ;
         LAYER metal3 ;
         RECT  21.3125 25.1575 21.4475 25.2925 ;
         LAYER metal4 ;
         RECT  131.755 5.85 131.895 20.81 ;
         LAYER metal3 ;
         RECT  80.9925 2.4725 81.1275 2.6075 ;
         LAYER metal3 ;
         RECT  123.1775 130.6375 123.3125 130.7725 ;
         LAYER metal3 ;
         RECT  125.4625 43.0975 125.5975 43.2325 ;
         LAYER metal4 ;
         RECT  15.21 44.59 15.35 59.55 ;
         LAYER metal3 ;
         RECT  21.3125 40.1075 21.4475 40.2425 ;
         LAYER metal3 ;
         RECT  125.4625 22.1675 125.5975 22.3025 ;
         LAYER metal4 ;
         RECT  119.905 20.67 120.045 116.56 ;
         LAYER metal3 ;
         RECT  35.2325 2.4725 35.3675 2.6075 ;
         LAYER metal3 ;
         RECT  27.485 19.965 27.62 20.1 ;
         LAYER metal4 ;
         RECT  146.4175 102.26 146.5575 124.6625 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal4 ;
         RECT  129.035 122.02 129.175 132.04 ;
         LAYER metal3 ;
         RECT  31.4925 19.1775 31.6275 19.3125 ;
         LAYER metal3 ;
         RECT  21.3125 34.1275 21.4475 34.2625 ;
         LAYER metal3 ;
         RECT  21.3125 31.1375 21.4475 31.2725 ;
         LAYER metal3 ;
         RECT  20.9325 2.4725 21.0675 2.6075 ;
         LAYER metal4 ;
         RECT  32.57 17.5 32.71 119.41 ;
         LAYER metal3 ;
         RECT  125.4625 34.1275 125.5975 34.2625 ;
         LAYER metal3 ;
         RECT  32.6375 16.805 111.1225 16.875 ;
         LAYER metal4 ;
         RECT  26.865 20.67 27.005 116.56 ;
         LAYER metal3 ;
         RECT  144.685 131.9025 144.82 132.0375 ;
         LAYER metal3 ;
         RECT  69.5525 2.4725 69.6875 2.6075 ;
         LAYER metal4 ;
         RECT  115.28 20.67 115.42 116.49 ;
         LAYER metal4 ;
         RECT  31.49 20.67 31.63 116.49 ;
         LAYER metal3 ;
         RECT  32.6375 8.415 109.4775 8.485 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  24.93 20.6375 25.07 116.56 ;
         LAYER metal3 ;
         RECT  19.785 26.6525 19.92 26.7875 ;
         LAYER metal3 ;
         RECT  106.7325 0.0025 106.8675 0.1375 ;
         LAYER metal4 ;
         RECT  140.86 119.55 141.0 134.51 ;
         LAYER metal3 ;
         RECT  19.785 41.6025 19.92 41.7375 ;
         LAYER metal3 ;
         RECT  121.2 127.4075 121.335 127.5425 ;
         LAYER metal3 ;
         RECT  19.785 38.6125 19.92 38.7475 ;
         LAYER metal3 ;
         RECT  83.8525 0.0025 83.9875 0.1375 ;
         LAYER metal3 ;
         RECT  32.6375 10.465 109.4775 10.535 ;
         LAYER metal3 ;
         RECT  32.6375 14.185 111.155 14.255 ;
         LAYER metal4 ;
         RECT  18.07 44.525 18.21 59.615 ;
         LAYER metal4 ;
         RECT  27.425 20.6375 27.565 116.5225 ;
         LAYER metal4 ;
         RECT  113.74 17.5 113.88 119.41 ;
         LAYER metal3 ;
         RECT  126.99 26.6525 127.125 26.7875 ;
         LAYER metal4 ;
         RECT  33.03 17.5 33.17 119.41 ;
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal3 ;
         RECT  19.785 20.6725 19.92 20.8075 ;
         LAYER metal3 ;
         RECT  144.685 134.3725 144.82 134.5075 ;
         LAYER metal3 ;
         RECT  120.3175 133.1075 120.4525 133.2425 ;
         LAYER metal3 ;
         RECT  49.5325 0.0025 49.6675 0.1375 ;
         LAYER metal4 ;
         RECT  128.895 5.785 129.035 20.875 ;
         LAYER metal4 ;
         RECT  121.84 20.6375 121.98 116.56 ;
         LAYER metal3 ;
         RECT  126.99 29.6425 127.125 29.7775 ;
         LAYER metal3 ;
         RECT  126.99 44.5925 127.125 44.7275 ;
         LAYER metal3 ;
         RECT  121.2 122.4675 121.335 122.6025 ;
         LAYER metal3 ;
         RECT  32.6375 122.725 111.155 122.795 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal3 ;
         RECT  23.7925 0.0025 23.9275 0.1375 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal3 ;
         RECT  19.785 32.6325 19.92 32.7675 ;
         LAYER metal3 ;
         RECT  126.99 23.6625 127.125 23.7975 ;
         LAYER metal3 ;
         RECT  25.575 14.3775 25.71 14.5125 ;
         LAYER metal4 ;
         RECT  144.355 102.2275 144.495 124.63 ;
         LAYER metal3 ;
         RECT  19.785 29.6425 19.92 29.7775 ;
         LAYER metal3 ;
         RECT  72.4125 0.0025 72.5475 0.1375 ;
         LAYER metal3 ;
         RECT  95.2925 0.0025 95.4275 0.1375 ;
         LAYER metal3 ;
         RECT  25.575 9.4375 25.71 9.5725 ;
         LAYER metal3 ;
         RECT  126.99 41.6025 127.125 41.7375 ;
         LAYER metal3 ;
         RECT  38.0925 0.0025 38.2275 0.1375 ;
         LAYER metal3 ;
         RECT  60.9725 0.0025 61.1075 0.1375 ;
         LAYER metal3 ;
         RECT  126.99 20.6725 127.125 20.8075 ;
         LAYER metal3 ;
         RECT  32.6375 125.065 109.5125 125.135 ;
         LAYER metal3 ;
         RECT  126.99 35.6225 127.125 35.7575 ;
         LAYER metal3 ;
         RECT  19.785 23.6625 19.92 23.7975 ;
         LAYER metal3 ;
         RECT  26.6525 0.0025 26.7875 0.1375 ;
         LAYER metal3 ;
         RECT  19.785 44.5925 19.92 44.7275 ;
         LAYER metal4 ;
         RECT  119.345 20.6375 119.485 116.5225 ;
         LAYER metal3 ;
         RECT  19.785 35.6225 19.92 35.7575 ;
         LAYER metal3 ;
         RECT  126.99 32.6325 127.125 32.7675 ;
         LAYER metal3 ;
         RECT  126.99 38.6125 127.125 38.7475 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 147.105 134.37 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 147.105 134.37 ;
   LAYER  metal3 ;
      RECT  24.35 0.9675 26.795 1.3825 ;
      RECT  27.21 0.9675 29.655 1.3825 ;
      RECT  30.07 0.9675 32.515 1.3825 ;
      RECT  32.93 0.9675 35.375 1.3825 ;
      RECT  35.79 0.9675 38.235 1.3825 ;
      RECT  38.65 0.9675 41.095 1.3825 ;
      RECT  41.51 0.9675 43.955 1.3825 ;
      RECT  44.37 0.9675 46.815 1.3825 ;
      RECT  47.23 0.9675 49.675 1.3825 ;
      RECT  50.09 0.9675 52.535 1.3825 ;
      RECT  52.95 0.9675 55.395 1.3825 ;
      RECT  55.81 0.9675 58.255 1.3825 ;
      RECT  58.67 0.9675 61.115 1.3825 ;
      RECT  61.53 0.9675 63.975 1.3825 ;
      RECT  64.39 0.9675 66.835 1.3825 ;
      RECT  67.25 0.9675 69.695 1.3825 ;
      RECT  70.11 0.9675 72.555 1.3825 ;
      RECT  72.97 0.9675 75.415 1.3825 ;
      RECT  75.83 0.9675 78.275 1.3825 ;
      RECT  78.69 0.9675 81.135 1.3825 ;
      RECT  81.55 0.9675 83.995 1.3825 ;
      RECT  84.41 0.9675 86.855 1.3825 ;
      RECT  87.27 0.9675 89.715 1.3825 ;
      RECT  90.13 0.9675 92.575 1.3825 ;
      RECT  92.99 0.9675 95.435 1.3825 ;
      RECT  95.85 0.9675 98.295 1.3825 ;
      RECT  98.71 0.9675 101.155 1.3825 ;
      RECT  101.57 0.9675 104.015 1.3825 ;
      RECT  104.43 0.9675 106.875 1.3825 ;
      RECT  107.29 0.9675 109.735 1.3825 ;
      RECT  110.15 0.9675 112.595 1.3825 ;
      RECT  113.01 0.9675 147.105 1.3825 ;
      RECT  21.49 0.9675 23.935 1.3825 ;
      RECT  0.14 45.5575 15.355 45.9725 ;
      RECT  0.14 45.9725 15.355 134.37 ;
      RECT  15.355 1.3825 15.77 45.5575 ;
      RECT  15.77 45.5575 23.935 45.9725 ;
      RECT  15.77 45.9725 23.935 134.37 ;
      RECT  15.355 45.9725 15.77 48.2875 ;
      RECT  15.355 48.7025 15.77 50.4975 ;
      RECT  15.355 50.9125 15.77 53.2275 ;
      RECT  15.355 53.6425 15.77 55.4375 ;
      RECT  15.355 55.8525 15.77 58.1675 ;
      RECT  15.355 58.5825 15.77 134.37 ;
      RECT  24.35 131.8625 122.755 132.2775 ;
      RECT  122.755 132.2775 123.17 134.37 ;
      RECT  123.17 1.3825 131.335 19.4275 ;
      RECT  123.17 19.4275 131.335 19.8425 ;
      RECT  131.335 19.8425 131.75 131.8625 ;
      RECT  131.75 1.3825 147.105 19.4275 ;
      RECT  131.75 19.4275 147.105 19.8425 ;
      RECT  131.335 17.1125 131.75 19.4275 ;
      RECT  131.335 14.9025 131.75 16.6975 ;
      RECT  131.335 12.1725 131.75 14.4875 ;
      RECT  131.335 9.9625 131.75 11.7575 ;
      RECT  131.335 1.3825 131.75 6.8175 ;
      RECT  131.335 7.2325 131.75 9.5475 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  146.685 132.2775 147.1 133.1275 ;
      RECT  146.685 133.5425 147.1 134.37 ;
      RECT  147.1 132.2775 147.105 133.1275 ;
      RECT  147.1 133.1275 147.105 133.5425 ;
      RECT  147.1 133.5425 147.105 134.37 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 45.5575 ;
      RECT  6.5225 1.3825 15.355 1.4675 ;
      RECT  6.5225 1.4675 15.355 45.5575 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 21.075 1.0525 ;
      RECT  6.5225 1.0525 21.075 1.3825 ;
      RECT  123.17 132.2775 140.5825 133.0425 ;
      RECT  123.17 133.0425 140.5825 133.1275 ;
      RECT  140.5825 132.2775 140.9975 133.0425 ;
      RECT  140.9975 132.2775 146.685 133.0425 ;
      RECT  140.9975 133.0425 146.685 133.1275 ;
      RECT  123.17 133.1275 140.5825 133.4575 ;
      RECT  123.17 133.4575 140.5825 133.5425 ;
      RECT  140.5825 133.4575 140.9975 133.5425 ;
      RECT  140.9975 133.1275 146.685 133.4575 ;
      RECT  140.9975 133.4575 146.685 133.5425 ;
      RECT  24.35 129.375 35.6825 129.79 ;
      RECT  24.35 129.79 35.6825 131.8625 ;
      RECT  35.6825 129.79 36.0975 131.8625 ;
      RECT  36.0975 129.79 122.755 131.8625 ;
      RECT  36.0975 129.375 38.0325 129.79 ;
      RECT  38.4475 129.375 40.3825 129.79 ;
      RECT  40.7975 129.375 42.7325 129.79 ;
      RECT  43.1475 129.375 45.0825 129.79 ;
      RECT  45.4975 129.375 47.4325 129.79 ;
      RECT  47.8475 129.375 49.7825 129.79 ;
      RECT  50.1975 129.375 52.1325 129.79 ;
      RECT  52.5475 129.375 54.4825 129.79 ;
      RECT  54.8975 129.375 56.8325 129.79 ;
      RECT  57.2475 129.375 59.1825 129.79 ;
      RECT  59.5975 129.375 61.5325 129.79 ;
      RECT  61.9475 129.375 63.8825 129.79 ;
      RECT  64.2975 129.375 66.2325 129.79 ;
      RECT  66.6475 129.375 68.5825 129.79 ;
      RECT  68.9975 129.375 70.9325 129.79 ;
      RECT  71.3475 129.375 73.2825 129.79 ;
      RECT  73.6975 129.375 75.6325 129.79 ;
      RECT  76.0475 129.375 77.9825 129.79 ;
      RECT  78.3975 129.375 80.3325 129.79 ;
      RECT  80.7475 129.375 82.6825 129.79 ;
      RECT  83.0975 129.375 85.0325 129.79 ;
      RECT  85.4475 129.375 87.3825 129.79 ;
      RECT  87.7975 129.375 89.7325 129.79 ;
      RECT  90.1475 129.375 92.0825 129.79 ;
      RECT  92.4975 129.375 94.4325 129.79 ;
      RECT  94.8475 129.375 96.7825 129.79 ;
      RECT  97.1975 129.375 99.1325 129.79 ;
      RECT  99.5475 129.375 101.4825 129.79 ;
      RECT  101.8975 129.375 103.8325 129.79 ;
      RECT  104.2475 129.375 106.1825 129.79 ;
      RECT  106.5975 129.375 108.5325 129.79 ;
      RECT  108.9475 129.375 122.755 129.79 ;
      RECT  123.17 19.8425 125.3225 30.9975 ;
      RECT  123.17 30.9975 125.3225 31.4125 ;
      RECT  125.7375 30.9975 131.335 31.4125 ;
      RECT  24.35 119.965 32.4975 120.315 ;
      RECT  24.35 120.315 32.4975 129.375 ;
      RECT  112.4375 119.965 122.755 120.315 ;
      RECT  15.77 22.0275 21.1725 22.4425 ;
      RECT  21.5875 22.0275 23.935 22.4425 ;
      RECT  21.5875 22.4425 23.935 45.5575 ;
      RECT  23.935 1.3825 24.0675 2.3325 ;
      RECT  23.935 2.7475 24.0675 134.37 ;
      RECT  24.0675 1.3825 24.35 2.3325 ;
      RECT  24.0675 2.3325 24.35 2.7475 ;
      RECT  24.0675 2.7475 24.35 134.37 ;
      RECT  21.5875 1.3825 23.6525 2.3325 ;
      RECT  21.5875 2.3325 23.6525 2.7475 ;
      RECT  21.5875 2.7475 23.6525 22.0275 ;
      RECT  23.6525 1.3825 23.935 2.3325 ;
      RECT  23.6525 2.7475 23.935 22.0275 ;
      RECT  112.4375 1.3825 115.1425 117.7075 ;
      RECT  112.4375 117.7075 115.1425 118.1225 ;
      RECT  112.4375 118.1225 115.1425 119.965 ;
      RECT  115.1425 1.3825 115.5575 117.7075 ;
      RECT  115.1425 118.1225 115.5575 119.965 ;
      RECT  115.5575 117.7075 122.755 118.1225 ;
      RECT  115.5575 118.1225 122.755 119.965 ;
      RECT  24.35 1.3825 25.435 11.7675 ;
      RECT  24.35 11.7675 25.435 12.1825 ;
      RECT  24.35 12.1825 25.435 119.965 ;
      RECT  25.85 1.3825 32.4975 11.7675 ;
      RECT  25.85 11.7675 32.4975 12.1825 ;
      RECT  36.0975 1.3825 46.5325 2.3325 ;
      RECT  36.0975 2.3325 46.5325 2.7475 ;
      RECT  46.5325 1.3825 46.9475 2.3325 ;
      RECT  46.9475 1.3825 112.4375 2.3325 ;
      RECT  115.5575 1.3825 119.15 116.92 ;
      RECT  115.5575 116.92 119.15 117.335 ;
      RECT  115.5575 117.335 119.15 117.7075 ;
      RECT  119.15 1.3825 119.565 116.92 ;
      RECT  119.15 117.335 119.565 117.7075 ;
      RECT  119.565 1.3825 122.755 116.92 ;
      RECT  119.565 116.92 122.755 117.335 ;
      RECT  119.565 117.335 122.755 117.7075 ;
      RECT  21.1725 43.3725 21.5875 45.5575 ;
      RECT  92.7075 2.3325 103.7325 2.7475 ;
      RECT  104.1475 2.3325 112.4375 2.7475 ;
      RECT  46.9475 2.3325 57.9725 2.7475 ;
      RECT  125.3225 25.4325 125.7375 30.9975 ;
      RECT  112.4375 120.315 121.06 124.7975 ;
      RECT  112.4375 124.7975 121.06 125.2125 ;
      RECT  112.4375 125.2125 121.06 129.375 ;
      RECT  121.475 120.315 122.755 124.7975 ;
      RECT  121.475 124.7975 122.755 125.2125 ;
      RECT  121.475 125.2125 122.755 129.375 ;
      RECT  32.4975 127.1675 35.6825 129.375 ;
      RECT  35.6825 127.1675 36.0975 129.375 ;
      RECT  36.0975 127.1675 109.6175 129.375 ;
      RECT  109.6175 126.8175 112.4375 127.1675 ;
      RECT  109.6175 127.1675 112.4375 129.375 ;
      RECT  21.1725 22.4425 21.5875 25.0175 ;
      RECT  81.2675 2.3325 92.2925 2.7475 ;
      RECT  122.755 1.3825 123.0375 130.4975 ;
      RECT  122.755 130.4975 123.0375 130.9125 ;
      RECT  122.755 130.9125 123.0375 131.8625 ;
      RECT  123.0375 1.3825 123.17 130.4975 ;
      RECT  123.0375 130.9125 123.17 131.8625 ;
      RECT  123.17 31.4125 123.4525 130.4975 ;
      RECT  123.17 130.9125 123.4525 131.8625 ;
      RECT  123.4525 31.4125 125.3225 130.4975 ;
      RECT  123.4525 130.4975 125.3225 130.9125 ;
      RECT  123.4525 130.9125 125.3225 131.8625 ;
      RECT  125.3225 40.3825 125.7375 42.9575 ;
      RECT  125.3225 43.3725 125.7375 131.8625 ;
      RECT  21.1725 40.3825 21.5875 42.9575 ;
      RECT  125.3225 19.8425 125.7375 22.0275 ;
      RECT  125.3225 22.4425 125.7375 25.0175 ;
      RECT  32.4975 1.3825 35.0925 2.3325 ;
      RECT  32.4975 2.3325 35.0925 2.7475 ;
      RECT  35.0925 1.3825 35.5075 2.3325 ;
      RECT  35.5075 1.3825 35.6825 2.3325 ;
      RECT  35.5075 2.3325 35.6825 2.7475 ;
      RECT  25.85 12.1825 27.345 19.825 ;
      RECT  25.85 19.825 27.345 20.24 ;
      RECT  25.85 20.24 27.345 119.965 ;
      RECT  27.345 12.1825 27.76 19.825 ;
      RECT  27.345 20.24 27.76 119.965 ;
      RECT  27.76 19.825 32.4975 20.24 ;
      RECT  27.76 20.24 32.4975 119.965 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 45.5575 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 45.5575 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 45.5575 ;
      RECT  27.76 12.1825 31.3525 19.0375 ;
      RECT  27.76 19.0375 31.3525 19.4525 ;
      RECT  27.76 19.4525 31.3525 19.825 ;
      RECT  31.3525 12.1825 31.7675 19.0375 ;
      RECT  31.3525 19.4525 31.7675 19.825 ;
      RECT  31.7675 12.1825 32.4975 19.0375 ;
      RECT  31.7675 19.0375 32.4975 19.4525 ;
      RECT  31.7675 19.4525 32.4975 19.825 ;
      RECT  21.1725 34.4025 21.5875 39.9675 ;
      RECT  21.1725 25.4325 21.5875 30.9975 ;
      RECT  21.1725 31.4125 21.5875 33.9875 ;
      RECT  15.77 1.3825 20.7925 2.3325 ;
      RECT  15.77 2.3325 20.7925 2.7475 ;
      RECT  20.7925 1.3825 21.1725 2.3325 ;
      RECT  20.7925 2.7475 21.1725 22.0275 ;
      RECT  21.1725 1.3825 21.2075 2.3325 ;
      RECT  21.1725 2.7475 21.2075 22.0275 ;
      RECT  21.2075 1.3825 21.5875 2.3325 ;
      RECT  21.2075 2.3325 21.5875 2.7475 ;
      RECT  21.2075 2.7475 21.5875 22.0275 ;
      RECT  125.3225 31.4125 125.7375 33.9875 ;
      RECT  125.3225 34.4025 125.7375 39.9675 ;
      RECT  35.6825 17.015 36.0975 119.965 ;
      RECT  36.0975 17.015 46.5325 119.965 ;
      RECT  46.5325 17.015 46.9475 119.965 ;
      RECT  46.9475 17.015 111.2625 119.965 ;
      RECT  111.2625 16.665 112.4375 17.015 ;
      RECT  111.2625 17.015 112.4375 119.965 ;
      RECT  32.4975 17.015 35.0925 119.965 ;
      RECT  35.0925 17.015 35.5075 119.965 ;
      RECT  35.5075 17.015 35.6825 119.965 ;
      RECT  123.17 131.8625 144.545 132.1775 ;
      RECT  123.17 132.1775 144.545 132.2775 ;
      RECT  144.545 132.1775 144.96 132.2775 ;
      RECT  144.96 131.8625 147.105 132.1775 ;
      RECT  144.96 132.1775 147.105 132.2775 ;
      RECT  131.75 19.8425 144.545 131.7625 ;
      RECT  131.75 131.7625 144.545 131.8625 ;
      RECT  144.545 19.8425 144.96 131.7625 ;
      RECT  144.96 19.8425 147.105 131.7625 ;
      RECT  144.96 131.7625 147.105 131.8625 ;
      RECT  58.3875 2.3325 69.4125 2.7475 ;
      RECT  69.8275 2.3325 80.8525 2.7475 ;
      RECT  35.6825 1.3825 36.0975 8.275 ;
      RECT  36.0975 2.7475 46.5325 8.275 ;
      RECT  46.5325 2.7475 46.9475 8.275 ;
      RECT  46.9475 2.7475 109.6175 8.275 ;
      RECT  109.6175 2.7475 111.2625 8.275 ;
      RECT  109.6175 8.275 111.2625 8.625 ;
      RECT  32.4975 2.7475 35.0925 8.275 ;
      RECT  35.0925 2.7475 35.5075 8.275 ;
      RECT  35.5075 2.7475 35.6825 8.275 ;
      RECT  15.77 22.4425 19.645 26.5125 ;
      RECT  15.77 26.5125 19.645 26.9275 ;
      RECT  15.77 26.9275 19.645 45.5575 ;
      RECT  20.06 22.4425 21.1725 26.5125 ;
      RECT  20.06 26.5125 21.1725 26.9275 ;
      RECT  20.06 26.9275 21.1725 45.5575 ;
      RECT  24.35 0.2775 106.5925 0.9675 ;
      RECT  106.5925 0.2775 107.0075 0.9675 ;
      RECT  107.0075 0.14 147.105 0.2775 ;
      RECT  107.0075 0.2775 147.105 0.9675 ;
      RECT  121.06 125.2125 121.475 127.2675 ;
      RECT  121.06 127.6825 121.475 129.375 ;
      RECT  19.645 38.8875 20.06 41.4625 ;
      RECT  35.6825 8.625 36.0975 10.325 ;
      RECT  36.0975 8.625 46.5325 10.325 ;
      RECT  46.5325 8.625 46.9475 10.325 ;
      RECT  46.9475 8.625 109.6175 10.325 ;
      RECT  32.4975 8.625 35.0925 10.325 ;
      RECT  35.0925 8.625 35.5075 10.325 ;
      RECT  35.5075 8.625 35.6825 10.325 ;
      RECT  111.2625 2.7475 111.295 14.045 ;
      RECT  111.2625 14.395 111.295 16.665 ;
      RECT  111.295 2.7475 112.4375 14.045 ;
      RECT  111.295 14.045 112.4375 14.395 ;
      RECT  111.295 14.395 112.4375 16.665 ;
      RECT  109.6175 8.625 111.2625 14.045 ;
      RECT  109.6175 14.395 111.2625 16.665 ;
      RECT  35.6825 10.675 36.0975 14.045 ;
      RECT  35.6825 14.395 36.0975 16.665 ;
      RECT  36.0975 10.675 46.5325 14.045 ;
      RECT  36.0975 14.395 46.5325 16.665 ;
      RECT  46.5325 10.675 46.9475 14.045 ;
      RECT  46.5325 14.395 46.9475 16.665 ;
      RECT  46.9475 10.675 109.6175 14.045 ;
      RECT  46.9475 14.395 109.6175 16.665 ;
      RECT  32.4975 10.675 35.0925 14.045 ;
      RECT  32.4975 14.395 35.0925 16.665 ;
      RECT  35.0925 10.675 35.5075 14.045 ;
      RECT  35.0925 14.395 35.5075 16.665 ;
      RECT  35.5075 10.675 35.6825 14.045 ;
      RECT  35.5075 14.395 35.6825 16.665 ;
      RECT  125.7375 19.8425 126.85 26.5125 ;
      RECT  125.7375 26.5125 126.85 26.9275 ;
      RECT  125.7375 26.9275 126.85 30.9975 ;
      RECT  127.265 19.8425 131.335 26.5125 ;
      RECT  127.265 26.5125 131.335 26.9275 ;
      RECT  127.265 26.9275 131.335 30.9975 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  0.14 0.2775 2.285 0.9675 ;
      RECT  2.285 0.2775 2.7 0.9675 ;
      RECT  2.7 0.2775 23.935 0.9675 ;
      RECT  15.77 2.7475 19.645 20.5325 ;
      RECT  15.77 20.5325 19.645 20.9475 ;
      RECT  15.77 20.9475 19.645 22.0275 ;
      RECT  19.645 2.7475 20.06 20.5325 ;
      RECT  19.645 20.9475 20.06 22.0275 ;
      RECT  20.06 2.7475 20.7925 20.5325 ;
      RECT  20.06 20.5325 20.7925 20.9475 ;
      RECT  20.06 20.9475 20.7925 22.0275 ;
      RECT  123.17 133.5425 144.545 134.2325 ;
      RECT  123.17 134.2325 144.545 134.37 ;
      RECT  144.545 133.5425 144.96 134.2325 ;
      RECT  144.96 133.5425 146.685 134.2325 ;
      RECT  144.96 134.2325 146.685 134.37 ;
      RECT  24.35 132.2775 120.1775 132.9675 ;
      RECT  24.35 132.9675 120.1775 133.3825 ;
      RECT  24.35 133.3825 120.1775 134.37 ;
      RECT  120.1775 132.2775 120.5925 132.9675 ;
      RECT  120.1775 133.3825 120.5925 134.37 ;
      RECT  120.5925 132.2775 122.755 132.9675 ;
      RECT  120.5925 132.9675 122.755 133.3825 ;
      RECT  120.5925 133.3825 122.755 134.37 ;
      RECT  126.85 26.9275 127.265 29.5025 ;
      RECT  126.85 29.9175 127.265 30.9975 ;
      RECT  125.7375 31.4125 126.85 44.4525 ;
      RECT  125.7375 44.4525 126.85 44.8675 ;
      RECT  125.7375 44.8675 126.85 131.8625 ;
      RECT  126.85 44.8675 127.265 131.8625 ;
      RECT  127.265 31.4125 131.335 44.4525 ;
      RECT  127.265 44.4525 131.335 44.8675 ;
      RECT  127.265 44.8675 131.335 131.8625 ;
      RECT  121.06 120.315 121.475 122.3275 ;
      RECT  121.06 122.7425 121.475 124.7975 ;
      RECT  32.4975 120.315 35.6825 122.585 ;
      RECT  35.6825 120.315 36.0975 122.585 ;
      RECT  36.0975 120.315 109.6175 122.585 ;
      RECT  109.6175 120.315 111.295 122.585 ;
      RECT  111.295 120.315 112.4375 122.585 ;
      RECT  111.295 122.585 112.4375 122.935 ;
      RECT  111.295 122.935 112.4375 126.8175 ;
      RECT  23.935 0.2775 24.0675 0.9675 ;
      RECT  24.0675 0.14 24.35 0.2775 ;
      RECT  24.0675 0.2775 24.35 0.9675 ;
      RECT  2.7 0.14 23.6525 0.2775 ;
      RECT  126.85 23.9375 127.265 26.5125 ;
      RECT  25.435 12.1825 25.85 14.2375 ;
      RECT  25.435 14.6525 25.85 119.965 ;
      RECT  19.645 26.9275 20.06 29.5025 ;
      RECT  19.645 29.9175 20.06 32.4925 ;
      RECT  72.6875 0.14 83.7125 0.2775 ;
      RECT  84.1275 0.14 95.1525 0.2775 ;
      RECT  95.5675 0.14 106.5925 0.2775 ;
      RECT  25.435 1.3825 25.85 9.2975 ;
      RECT  25.435 9.7125 25.85 11.7675 ;
      RECT  126.85 41.8775 127.265 44.4525 ;
      RECT  38.3675 0.14 49.3925 0.2775 ;
      RECT  49.8075 0.14 60.8325 0.2775 ;
      RECT  61.2475 0.14 72.2725 0.2775 ;
      RECT  126.85 19.8425 127.265 20.5325 ;
      RECT  126.85 20.9475 127.265 23.5225 ;
      RECT  32.4975 122.935 35.6825 124.925 ;
      RECT  32.4975 125.275 35.6825 126.8175 ;
      RECT  35.6825 122.935 36.0975 124.925 ;
      RECT  35.6825 125.275 36.0975 126.8175 ;
      RECT  36.0975 122.935 109.6175 124.925 ;
      RECT  36.0975 125.275 109.6175 126.8175 ;
      RECT  109.6175 122.935 109.6525 124.925 ;
      RECT  109.6175 125.275 109.6525 126.8175 ;
      RECT  109.6525 122.935 111.295 124.925 ;
      RECT  109.6525 124.925 111.295 125.275 ;
      RECT  109.6525 125.275 111.295 126.8175 ;
      RECT  19.645 22.4425 20.06 23.5225 ;
      RECT  19.645 23.9375 20.06 26.5125 ;
      RECT  24.35 0.14 26.5125 0.2775 ;
      RECT  26.9275 0.14 37.9525 0.2775 ;
      RECT  19.645 41.8775 20.06 44.4525 ;
      RECT  19.645 44.8675 20.06 45.5575 ;
      RECT  19.645 32.9075 20.06 35.4825 ;
      RECT  19.645 35.8975 20.06 38.4725 ;
      RECT  126.85 31.4125 127.265 32.4925 ;
      RECT  126.85 32.9075 127.265 35.4825 ;
      RECT  126.85 35.8975 127.265 38.4725 ;
      RECT  126.85 38.8875 127.265 41.4625 ;
   LAYER  metal4 ;
      RECT  17.65 0.14 18.35 2.19 ;
      RECT  18.35 0.14 147.105 2.19 ;
      RECT  18.35 2.19 113.92 17.22 ;
      RECT  113.92 2.19 114.62 17.22 ;
      RECT  18.35 119.69 113.92 134.37 ;
      RECT  113.92 119.69 114.62 134.37 ;
      RECT  131.475 2.19 132.175 5.57 ;
      RECT  132.175 2.19 147.105 5.57 ;
      RECT  132.175 5.57 147.105 17.22 ;
      RECT  132.175 17.22 147.105 17.71 ;
      RECT  131.475 21.09 132.175 119.69 ;
      RECT  132.175 17.71 147.105 21.09 ;
      RECT  0.14 44.31 14.93 59.83 ;
      RECT  0.14 59.83 14.93 134.37 ;
      RECT  14.93 17.71 15.63 44.31 ;
      RECT  14.93 59.83 15.63 134.37 ;
      RECT  15.63 17.71 17.65 44.31 ;
      RECT  15.63 44.31 17.65 59.83 ;
      RECT  15.63 59.83 17.65 134.37 ;
      RECT  114.62 116.84 119.625 119.69 ;
      RECT  119.625 116.84 120.325 119.69 ;
      RECT  120.325 116.84 131.475 119.69 ;
      RECT  146.1375 124.9425 146.8375 134.37 ;
      RECT  146.8375 119.69 147.105 124.9425 ;
      RECT  146.8375 124.9425 147.105 134.37 ;
      RECT  146.1375 21.09 146.8375 101.98 ;
      RECT  146.8375 21.09 147.105 101.98 ;
      RECT  146.8375 101.98 147.105 119.69 ;
      RECT  114.62 119.69 128.755 121.74 ;
      RECT  114.62 121.74 128.755 124.9425 ;
      RECT  128.755 119.69 129.455 121.74 ;
      RECT  114.62 124.9425 128.755 132.32 ;
      RECT  114.62 132.32 128.755 134.37 ;
      RECT  128.755 132.32 129.455 134.37 ;
      RECT  18.35 17.22 32.29 17.71 ;
      RECT  18.35 116.84 26.585 119.69 ;
      RECT  26.585 116.84 27.285 119.69 ;
      RECT  27.285 116.84 32.29 119.69 ;
      RECT  114.62 20.39 115.0 21.09 ;
      RECT  114.62 21.09 115.0 116.77 ;
      RECT  114.62 116.77 115.0 116.84 ;
      RECT  115.0 116.77 115.7 116.84 ;
      RECT  31.21 116.77 31.91 116.84 ;
      RECT  31.91 20.39 32.29 116.77 ;
      RECT  31.91 116.77 32.29 116.84 ;
      RECT  0.14 2.19 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 17.71 ;
      RECT  0.4075 2.19 1.1075 9.5675 ;
      RECT  0.14 17.71 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 44.31 ;
      RECT  0.4075 32.53 1.1075 44.31 ;
      RECT  18.35 17.71 24.65 20.3575 ;
      RECT  18.35 20.3575 24.65 20.39 ;
      RECT  24.65 17.71 25.35 20.3575 ;
      RECT  25.35 17.71 26.585 20.3575 ;
      RECT  25.35 20.3575 26.585 20.39 ;
      RECT  25.35 20.39 26.585 116.84 ;
      RECT  132.175 101.98 140.58 119.27 ;
      RECT  132.175 119.27 140.58 119.69 ;
      RECT  140.58 101.98 141.28 119.27 ;
      RECT  129.455 119.69 140.58 121.74 ;
      RECT  129.455 121.74 140.58 124.9425 ;
      RECT  129.455 124.9425 140.58 132.32 ;
      RECT  141.28 124.9425 146.1375 132.32 ;
      RECT  129.455 132.32 140.58 134.37 ;
      RECT  141.28 132.32 146.1375 134.37 ;
      RECT  17.65 17.71 17.79 44.245 ;
      RECT  17.65 44.245 17.79 59.895 ;
      RECT  17.65 59.895 17.79 134.37 ;
      RECT  17.79 17.71 18.35 44.245 ;
      RECT  17.79 59.895 18.35 134.37 ;
      RECT  18.35 20.39 18.49 44.245 ;
      RECT  18.35 59.895 18.49 116.84 ;
      RECT  18.49 20.39 24.65 44.245 ;
      RECT  18.49 44.245 24.65 59.895 ;
      RECT  18.49 59.895 24.65 116.84 ;
      RECT  26.585 17.71 27.145 20.3575 ;
      RECT  26.585 20.3575 27.145 20.39 ;
      RECT  27.145 17.71 27.285 20.3575 ;
      RECT  27.285 17.71 27.845 20.3575 ;
      RECT  27.845 17.71 32.29 20.3575 ;
      RECT  27.845 20.3575 32.29 20.39 ;
      RECT  27.845 20.39 31.21 116.77 ;
      RECT  27.285 116.8025 27.845 116.84 ;
      RECT  27.845 116.77 31.21 116.8025 ;
      RECT  27.845 116.8025 31.21 116.84 ;
      RECT  33.45 17.22 113.46 17.71 ;
      RECT  33.45 17.71 113.46 119.69 ;
      RECT  114.62 2.19 128.615 5.505 ;
      RECT  114.62 5.505 128.615 5.57 ;
      RECT  128.615 2.19 129.315 5.505 ;
      RECT  129.315 2.19 131.475 5.505 ;
      RECT  129.315 5.505 131.475 5.57 ;
      RECT  114.62 5.57 128.615 17.22 ;
      RECT  129.315 5.57 131.475 17.22 ;
      RECT  114.62 17.22 128.615 17.71 ;
      RECT  129.315 17.22 131.475 17.71 ;
      RECT  129.315 17.71 131.475 20.39 ;
      RECT  129.315 20.39 131.475 21.09 ;
      RECT  128.615 21.155 129.315 116.84 ;
      RECT  129.315 21.09 131.475 21.155 ;
      RECT  129.315 21.155 131.475 116.84 ;
      RECT  120.325 17.71 121.56 20.3575 ;
      RECT  120.325 20.3575 121.56 20.39 ;
      RECT  121.56 17.71 122.26 20.3575 ;
      RECT  122.26 17.71 128.615 20.3575 ;
      RECT  122.26 20.3575 128.615 20.39 ;
      RECT  120.325 20.39 121.56 21.09 ;
      RECT  122.26 20.39 128.615 21.09 ;
      RECT  120.325 21.09 121.56 21.155 ;
      RECT  122.26 21.09 128.615 21.155 ;
      RECT  120.325 21.155 121.56 116.84 ;
      RECT  122.26 21.155 128.615 116.84 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 17.71 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  1.1075 17.71 2.47 32.53 ;
      RECT  3.17 17.71 14.93 32.53 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 44.31 ;
      RECT  2.47 32.5625 3.17 44.31 ;
      RECT  3.17 32.53 14.93 32.5625 ;
      RECT  3.17 32.5625 14.93 44.31 ;
      RECT  0.14 0.14 5.825 2.19 ;
      RECT  6.525 0.14 17.65 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 17.65 9.5675 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  6.525 9.5675 17.65 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  3.17 15.24 5.825 17.71 ;
      RECT  5.825 15.24 6.525 17.71 ;
      RECT  6.525 9.6 17.65 15.24 ;
      RECT  6.525 15.24 17.65 17.71 ;
      RECT  132.175 21.09 144.075 101.9475 ;
      RECT  132.175 101.9475 144.075 101.98 ;
      RECT  144.075 21.09 144.775 101.9475 ;
      RECT  144.775 21.09 146.1375 101.9475 ;
      RECT  144.775 101.9475 146.1375 101.98 ;
      RECT  141.28 101.98 144.075 119.27 ;
      RECT  144.775 101.98 146.1375 119.27 ;
      RECT  141.28 119.27 144.075 119.69 ;
      RECT  144.775 119.27 146.1375 119.69 ;
      RECT  141.28 119.69 144.075 121.74 ;
      RECT  144.775 119.69 146.1375 121.74 ;
      RECT  141.28 121.74 144.075 124.91 ;
      RECT  141.28 124.91 144.075 124.9425 ;
      RECT  144.075 124.91 144.775 124.9425 ;
      RECT  144.775 121.74 146.1375 124.91 ;
      RECT  144.775 124.91 146.1375 124.9425 ;
      RECT  114.62 17.71 119.065 20.3575 ;
      RECT  114.62 20.3575 119.065 20.39 ;
      RECT  119.065 17.71 119.625 20.3575 ;
      RECT  119.625 17.71 119.765 20.3575 ;
      RECT  119.765 17.71 120.325 20.3575 ;
      RECT  119.765 20.3575 120.325 20.39 ;
      RECT  115.7 20.39 119.065 21.09 ;
      RECT  115.7 21.09 119.065 116.77 ;
      RECT  115.7 116.77 119.065 116.8025 ;
      RECT  115.7 116.8025 119.065 116.84 ;
      RECT  119.065 116.8025 119.625 116.84 ;
   END
END    freepdk45_sram_1w1r_128x32_32
END    LIBRARY
