VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_11x128
   CLASS BLOCK ;
   SIZE 114.955 BY 88.425 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.085 1.105 23.22 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  25.945 1.105 26.08 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.805 1.105 28.94 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.665 1.105 31.8 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.525 1.105 34.66 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.385 1.105 37.52 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.245 1.105 40.38 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.105 1.105 43.24 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.965 1.105 46.1 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.825 1.105 48.96 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.685 1.105 51.82 1.24 ;
      END
   END din0[10]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.365 1.105 17.5 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.225 1.105 20.36 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.645 43.09 11.78 43.225 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.645 45.82 11.78 45.955 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.645 48.03 11.78 48.165 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.645 50.76 11.78 50.895 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.645 52.97 11.78 53.105 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.455 87.185 94.59 87.32 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.595 87.185 91.73 87.32 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.035 19.95 103.17 20.085 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.035 17.22 103.17 17.355 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.035 15.01 103.17 15.145 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.035 12.28 103.17 12.415 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.035 10.07 103.17 10.205 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.49 0.42 1.625 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.535 85.81 114.67 85.945 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.575 6.3825 1.71 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.4325 85.725 108.5675 85.86 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.4275 82.3175 31.5625 82.4525 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.1275 82.3175 36.2625 82.4525 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.8275 82.3175 40.9625 82.4525 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.5275 82.3175 45.6625 82.4525 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.2275 82.3175 50.3625 82.4525 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.9275 82.3175 55.0625 82.4525 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.6275 82.3175 59.7625 82.4525 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.3275 82.3175 64.4625 82.4525 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.0275 82.3175 69.1625 82.4525 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.7275 82.3175 73.8625 82.4525 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.4275 82.3175 78.5625 82.4525 ;
      END
   END dout1[10]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  14.08 2.8525 14.22 17.8125 ;
         LAYER metal3 ;
         RECT  28.2425 79.76 79.2325 79.83 ;
         LAYER metal4 ;
         RECT  11.36 41.9825 11.5 54.5375 ;
         LAYER metal3 ;
         RECT  27.0975 19.56 27.2325 19.695 ;
         LAYER metal3 ;
         RECT  96.7425 40.49 96.8775 40.625 ;
         LAYER metal3 ;
         RECT  45.6825 2.47 45.8175 2.605 ;
         LAYER metal4 ;
         RECT  21.45 4.845 21.59 14.865 ;
         LAYER metal3 ;
         RECT  90.57 69.6025 90.705 69.7375 ;
         LAYER metal4 ;
         RECT  27.095 21.0525 27.235 69.0325 ;
         LAYER metal4 ;
         RECT  0.6875 10.23 0.8275 32.6325 ;
         LAYER metal4 ;
         RECT  93.03 75.04 93.17 85.06 ;
         LAYER metal3 ;
         RECT  96.7425 31.52 96.8775 31.655 ;
         LAYER metal3 ;
         RECT  17.7425 31.52 17.8775 31.655 ;
         LAYER metal4 ;
         RECT  86.305 17.8825 86.445 71.9525 ;
         LAYER metal3 ;
         RECT  96.3975 22.55 96.5325 22.685 ;
         LAYER metal4 ;
         RECT  100.595 74.5625 100.735 84.5825 ;
         LAYER metal3 ;
         RECT  28.2425 17.1875 83.2275 17.2575 ;
         LAYER metal3 ;
         RECT  96.7425 34.51 96.8775 34.645 ;
         LAYER metal3 ;
         RECT  87.3875 70.39 87.5225 70.525 ;
         LAYER metal3 ;
         RECT  17.7425 34.51 17.8775 34.645 ;
         LAYER metal4 ;
         RECT  23.295 21.0525 23.435 69.1025 ;
         LAYER metal3 ;
         RECT  34.2425 2.47 34.3775 2.605 ;
         LAYER metal3 ;
         RECT  2.425 2.855 2.56 2.99 ;
         LAYER metal3 ;
         RECT  28.2425 72.6475 84.4025 72.7175 ;
         LAYER metal4 ;
         RECT  28.175 17.8825 28.315 71.9525 ;
         LAYER metal3 ;
         RECT  112.395 84.445 112.53 84.58 ;
         LAYER metal3 ;
         RECT  28.2425 8.5375 79.2325 8.6075 ;
         LAYER metal3 ;
         RECT  96.3975 25.54 96.5325 25.675 ;
         LAYER metal3 ;
         RECT  22.8025 2.47 22.9375 2.605 ;
         LAYER metal3 ;
         RECT  18.0875 22.55 18.2225 22.685 ;
         LAYER metal3 ;
         RECT  17.7425 37.5 17.8775 37.635 ;
         LAYER metal3 ;
         RECT  17.7425 40.49 17.8775 40.625 ;
         LAYER metal4 ;
         RECT  114.1275 54.8025 114.2675 77.205 ;
         LAYER metal4 ;
         RECT  103.315 8.6375 103.455 21.1925 ;
         LAYER metal3 ;
         RECT  17.0825 2.47 17.2175 2.605 ;
         LAYER metal4 ;
         RECT  91.185 21.0525 91.325 69.1025 ;
         LAYER metal3 ;
         RECT  18.0875 25.54 18.2225 25.675 ;
         LAYER metal3 ;
         RECT  94.7375 85.82 94.8725 85.955 ;
         LAYER metal4 ;
         RECT  87.385 21.0525 87.525 69.0325 ;
         LAYER metal3 ;
         RECT  23.915 20.3475 24.05 20.4825 ;
         LAYER metal3 ;
         RECT  96.7425 37.5 96.8775 37.635 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  28.2425 75.2675 83.26 75.3375 ;
         LAYER metal3 ;
         RECT  37.1025 0.0 37.2375 0.135 ;
         LAYER metal3 ;
         RECT  15.935 33.015 16.07 33.15 ;
         LAYER metal3 ;
         RECT  48.5425 0.0 48.6775 0.135 ;
         LAYER metal3 ;
         RECT  97.925 27.035 98.06 27.17 ;
         LAYER metal4 ;
         RECT  21.705 21.02 21.845 69.1025 ;
         LAYER metal4 ;
         RECT  94.6925 74.9725 94.8325 85.1275 ;
         LAYER metal3 ;
         RECT  28.2425 14.5675 83.26 14.6375 ;
         LAYER metal3 ;
         RECT  2.425 0.385 2.56 0.52 ;
         LAYER metal3 ;
         RECT  28.2425 10.5875 79.2325 10.6575 ;
         LAYER metal4 ;
         RECT  85.845 17.8825 85.985 71.9525 ;
         LAYER metal3 ;
         RECT  15.935 30.025 16.07 30.16 ;
         LAYER metal4 ;
         RECT  14.22 41.9175 14.36 54.4725 ;
         LAYER metal3 ;
         RECT  16.56 24.045 16.695 24.18 ;
         LAYER metal3 ;
         RECT  28.2425 77.8675 79.2675 77.9375 ;
         LAYER metal3 ;
         RECT  25.6625 0.0 25.7975 0.135 ;
         LAYER metal3 ;
         RECT  16.56 21.055 16.695 21.19 ;
         LAYER metal3 ;
         RECT  112.395 86.915 112.53 87.05 ;
         LAYER metal4 ;
         RECT  92.775 21.02 92.915 69.1025 ;
         LAYER metal4 ;
         RECT  2.75 10.2625 2.89 32.665 ;
         LAYER metal4 ;
         RECT  112.065 54.77 112.205 77.1725 ;
         LAYER metal3 ;
         RECT  98.55 41.985 98.685 42.12 ;
         LAYER metal3 ;
         RECT  98.55 36.005 98.685 36.14 ;
         LAYER metal3 ;
         RECT  19.9425 0.0 20.0775 0.135 ;
         LAYER metal4 ;
         RECT  100.455 8.7025 100.595 21.2575 ;
         LAYER metal4 ;
         RECT  23.855 21.02 23.995 69.065 ;
         LAYER metal3 ;
         RECT  15.935 38.995 16.07 39.13 ;
         LAYER metal4 ;
         RECT  108.57 72.0925 108.71 87.0525 ;
         LAYER metal3 ;
         RECT  98.55 38.995 98.685 39.13 ;
         LAYER metal3 ;
         RECT  97.925 21.055 98.06 21.19 ;
         LAYER metal4 ;
         RECT  19.7875 4.7775 19.9275 14.9325 ;
         LAYER metal3 ;
         RECT  15.935 36.005 16.07 36.14 ;
         LAYER metal4 ;
         RECT  90.625 21.02 90.765 69.065 ;
         LAYER metal3 ;
         RECT  16.56 27.035 16.695 27.17 ;
         LAYER metal3 ;
         RECT  91.8775 88.29 92.0125 88.425 ;
         LAYER metal3 ;
         RECT  15.935 41.985 16.07 42.12 ;
         LAYER metal3 ;
         RECT  98.55 30.025 98.685 30.16 ;
         LAYER metal3 ;
         RECT  97.925 24.045 98.06 24.18 ;
         LAYER metal3 ;
         RECT  98.55 33.015 98.685 33.15 ;
         LAYER metal4 ;
         RECT  28.635 17.8825 28.775 71.9525 ;
         LAYER metal4 ;
         RECT  6.105 0.3825 6.245 15.3425 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 114.815 88.285 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 114.815 88.285 ;
   LAYER  metal3 ;
      RECT  22.945 0.14 23.36 0.965 ;
      RECT  23.36 0.965 25.805 1.38 ;
      RECT  26.22 0.965 28.665 1.38 ;
      RECT  29.08 0.965 31.525 1.38 ;
      RECT  31.94 0.965 34.385 1.38 ;
      RECT  34.8 0.965 37.245 1.38 ;
      RECT  37.66 0.965 40.105 1.38 ;
      RECT  40.52 0.965 42.965 1.38 ;
      RECT  43.38 0.965 45.825 1.38 ;
      RECT  46.24 0.965 48.685 1.38 ;
      RECT  49.1 0.965 51.545 1.38 ;
      RECT  51.96 0.965 114.815 1.38 ;
      RECT  17.64 0.965 20.085 1.38 ;
      RECT  20.5 0.965 22.945 1.38 ;
      RECT  0.14 42.95 11.505 43.365 ;
      RECT  0.14 43.365 11.505 88.285 ;
      RECT  11.505 1.38 11.92 42.95 ;
      RECT  11.92 42.95 22.945 43.365 ;
      RECT  11.92 43.365 22.945 88.285 ;
      RECT  11.505 43.365 11.92 45.68 ;
      RECT  11.505 46.095 11.92 47.89 ;
      RECT  11.505 48.305 11.92 50.62 ;
      RECT  11.505 51.035 11.92 52.83 ;
      RECT  11.505 53.245 11.92 88.285 ;
      RECT  94.315 87.46 94.73 88.285 ;
      RECT  94.73 87.46 114.815 88.285 ;
      RECT  23.36 87.045 91.455 87.46 ;
      RECT  91.87 87.045 94.315 87.46 ;
      RECT  94.73 1.38 102.895 19.81 ;
      RECT  94.73 19.81 102.895 20.225 ;
      RECT  102.895 20.225 103.31 87.045 ;
      RECT  103.31 1.38 114.815 19.81 ;
      RECT  103.31 19.81 114.815 20.225 ;
      RECT  102.895 17.495 103.31 19.81 ;
      RECT  102.895 15.285 103.31 17.08 ;
      RECT  102.895 12.555 103.31 14.87 ;
      RECT  102.895 1.38 103.31 9.93 ;
      RECT  102.895 10.345 103.31 12.14 ;
      RECT  0.14 0.965 0.145 1.35 ;
      RECT  0.14 1.35 0.145 1.38 ;
      RECT  0.145 0.965 0.56 1.35 ;
      RECT  0.56 0.965 17.225 1.35 ;
      RECT  0.56 1.35 17.225 1.38 ;
      RECT  0.14 1.38 0.145 1.765 ;
      RECT  0.14 1.765 0.145 42.95 ;
      RECT  0.145 1.765 0.56 42.95 ;
      RECT  114.395 20.225 114.81 85.67 ;
      RECT  114.395 86.085 114.81 87.045 ;
      RECT  114.81 20.225 114.815 85.67 ;
      RECT  114.81 85.67 114.815 86.085 ;
      RECT  114.81 86.085 114.815 87.045 ;
      RECT  0.56 1.38 6.1075 1.435 ;
      RECT  0.56 1.435 6.1075 1.765 ;
      RECT  6.1075 1.38 6.5225 1.435 ;
      RECT  6.5225 1.38 11.505 1.435 ;
      RECT  6.5225 1.435 11.505 1.765 ;
      RECT  0.56 1.765 6.1075 1.85 ;
      RECT  6.1075 1.85 6.5225 42.95 ;
      RECT  6.5225 1.765 11.505 1.85 ;
      RECT  6.5225 1.85 11.505 42.95 ;
      RECT  103.31 20.225 108.2925 85.585 ;
      RECT  103.31 85.585 108.2925 85.67 ;
      RECT  108.2925 20.225 108.7075 85.585 ;
      RECT  108.7075 85.585 114.395 85.67 ;
      RECT  103.31 85.67 108.2925 86.0 ;
      RECT  103.31 86.0 108.2925 86.085 ;
      RECT  108.2925 86.0 108.7075 86.085 ;
      RECT  108.7075 85.67 114.395 86.0 ;
      RECT  108.7075 86.0 114.395 86.085 ;
      RECT  23.36 82.1775 31.2875 82.5925 ;
      RECT  23.36 82.5925 31.2875 87.045 ;
      RECT  31.2875 82.5925 31.7025 87.045 ;
      RECT  31.7025 82.5925 94.315 87.045 ;
      RECT  31.7025 82.1775 35.9875 82.5925 ;
      RECT  36.4025 82.1775 40.6875 82.5925 ;
      RECT  41.1025 82.1775 45.3875 82.5925 ;
      RECT  45.8025 82.1775 50.0875 82.5925 ;
      RECT  50.5025 82.1775 54.7875 82.5925 ;
      RECT  55.2025 82.1775 59.4875 82.5925 ;
      RECT  59.9025 82.1775 64.1875 82.5925 ;
      RECT  64.6025 82.1775 68.8875 82.5925 ;
      RECT  69.3025 82.1775 73.5875 82.5925 ;
      RECT  74.0025 82.1775 78.2875 82.5925 ;
      RECT  78.7025 82.1775 94.315 82.5925 ;
      RECT  23.36 79.62 28.1025 79.97 ;
      RECT  23.36 79.97 28.1025 82.1775 ;
      RECT  28.1025 79.97 31.2875 82.1775 ;
      RECT  31.2875 79.97 31.7025 82.1775 ;
      RECT  31.7025 79.97 79.3725 82.1775 ;
      RECT  79.3725 79.62 94.315 79.97 ;
      RECT  79.3725 79.97 94.315 82.1775 ;
      RECT  23.36 1.38 26.9575 19.42 ;
      RECT  23.36 19.42 26.9575 19.835 ;
      RECT  26.9575 1.38 27.3725 19.42 ;
      RECT  26.9575 19.835 27.3725 79.62 ;
      RECT  27.3725 1.38 28.1025 19.42 ;
      RECT  27.3725 19.42 28.1025 19.835 ;
      RECT  27.3725 19.835 28.1025 79.62 ;
      RECT  94.73 40.35 96.6025 40.765 ;
      RECT  96.6025 40.765 97.0175 87.045 ;
      RECT  97.0175 40.35 102.895 40.765 ;
      RECT  31.7025 1.38 45.5425 2.33 ;
      RECT  45.5425 1.38 45.9575 2.33 ;
      RECT  45.9575 1.38 79.3725 2.33 ;
      RECT  45.9575 2.33 79.3725 2.745 ;
      RECT  79.3725 69.4625 90.43 69.8775 ;
      RECT  90.43 1.38 90.845 69.4625 ;
      RECT  90.43 69.8775 90.845 79.62 ;
      RECT  90.845 1.38 94.315 69.4625 ;
      RECT  90.845 69.4625 94.315 69.8775 ;
      RECT  90.845 69.8775 94.315 79.62 ;
      RECT  11.92 31.38 17.6025 31.795 ;
      RECT  18.0175 31.38 22.945 31.795 ;
      RECT  18.0175 31.795 22.945 42.95 ;
      RECT  94.73 20.225 96.2575 22.41 ;
      RECT  94.73 22.41 96.2575 22.825 ;
      RECT  94.73 22.825 96.2575 40.35 ;
      RECT  96.2575 20.225 96.6025 22.41 ;
      RECT  96.6025 20.225 96.6725 22.41 ;
      RECT  96.6725 20.225 97.0175 22.41 ;
      RECT  96.6725 22.41 97.0175 22.825 ;
      RECT  96.6725 22.825 97.0175 31.38 ;
      RECT  79.3725 17.3975 83.3675 69.4625 ;
      RECT  83.3675 17.0475 90.43 17.3975 ;
      RECT  83.3675 17.3975 90.43 69.4625 ;
      RECT  96.6025 31.795 97.0175 34.37 ;
      RECT  79.3725 69.8775 87.2475 70.25 ;
      RECT  79.3725 70.25 87.2475 70.665 ;
      RECT  87.2475 69.8775 87.6625 70.25 ;
      RECT  87.2475 70.665 87.6625 79.62 ;
      RECT  87.6625 69.8775 90.43 70.25 ;
      RECT  87.6625 70.25 90.43 70.665 ;
      RECT  87.6625 70.665 90.43 79.62 ;
      RECT  17.6025 31.795 18.0175 34.37 ;
      RECT  31.7025 2.33 34.1025 2.745 ;
      RECT  34.5175 2.33 45.5425 2.745 ;
      RECT  0.56 1.85 2.285 2.715 ;
      RECT  0.56 2.715 2.285 3.13 ;
      RECT  0.56 3.13 2.285 42.95 ;
      RECT  2.285 1.85 2.7 2.715 ;
      RECT  2.285 3.13 2.7 42.95 ;
      RECT  2.7 1.85 6.1075 2.715 ;
      RECT  2.7 2.715 6.1075 3.13 ;
      RECT  2.7 3.13 6.1075 42.95 ;
      RECT  28.1025 17.3975 31.2875 72.5075 ;
      RECT  31.2875 17.3975 31.7025 72.5075 ;
      RECT  31.7025 17.3975 45.5425 72.5075 ;
      RECT  45.5425 17.3975 45.9575 72.5075 ;
      RECT  45.9575 17.3975 79.3725 72.5075 ;
      RECT  79.3725 70.665 84.5425 72.5075 ;
      RECT  84.5425 70.665 87.2475 72.5075 ;
      RECT  84.5425 72.5075 87.2475 72.8575 ;
      RECT  84.5425 72.8575 87.2475 79.62 ;
      RECT  108.7075 20.225 112.255 84.305 ;
      RECT  108.7075 84.305 112.255 84.72 ;
      RECT  108.7075 84.72 112.255 85.585 ;
      RECT  112.255 20.225 112.67 84.305 ;
      RECT  112.255 84.72 112.67 85.585 ;
      RECT  112.67 20.225 114.395 84.305 ;
      RECT  112.67 84.305 114.395 84.72 ;
      RECT  112.67 84.72 114.395 85.585 ;
      RECT  28.1025 1.38 31.2875 8.3975 ;
      RECT  31.2875 1.38 31.7025 8.3975 ;
      RECT  31.7025 2.745 45.5425 8.3975 ;
      RECT  45.5425 2.745 45.9575 8.3975 ;
      RECT  45.9575 2.745 79.3725 8.3975 ;
      RECT  96.2575 22.825 96.6025 25.4 ;
      RECT  96.2575 25.815 96.6025 40.35 ;
      RECT  96.6025 22.825 96.6725 25.4 ;
      RECT  96.6025 25.815 96.6725 31.38 ;
      RECT  22.945 1.38 23.0775 2.33 ;
      RECT  22.945 2.745 23.0775 88.285 ;
      RECT  23.0775 1.38 23.36 2.33 ;
      RECT  23.0775 2.33 23.36 2.745 ;
      RECT  23.0775 2.745 23.36 88.285 ;
      RECT  18.0175 1.38 22.6625 2.33 ;
      RECT  18.0175 2.33 22.6625 2.745 ;
      RECT  22.6625 1.38 22.945 2.33 ;
      RECT  22.6625 2.745 22.945 31.38 ;
      RECT  17.6025 1.38 17.9475 22.41 ;
      RECT  17.6025 22.41 17.9475 22.825 ;
      RECT  17.6025 22.825 17.9475 31.38 ;
      RECT  17.9475 1.38 18.0175 22.41 ;
      RECT  18.0175 2.745 18.3625 22.41 ;
      RECT  18.3625 2.745 22.6625 22.41 ;
      RECT  18.3625 22.41 22.6625 22.825 ;
      RECT  18.3625 22.825 22.6625 31.38 ;
      RECT  17.6025 34.785 18.0175 37.36 ;
      RECT  17.6025 37.775 18.0175 40.35 ;
      RECT  17.6025 40.765 18.0175 42.95 ;
      RECT  11.92 1.38 16.9425 2.33 ;
      RECT  11.92 2.33 16.9425 2.745 ;
      RECT  16.9425 1.38 17.3575 2.33 ;
      RECT  16.9425 2.745 17.3575 31.38 ;
      RECT  17.3575 1.38 17.6025 2.33 ;
      RECT  17.3575 2.33 17.6025 2.745 ;
      RECT  17.3575 2.745 17.6025 31.38 ;
      RECT  17.9475 22.825 18.0175 25.4 ;
      RECT  17.9475 25.815 18.0175 31.38 ;
      RECT  18.0175 22.825 18.3625 25.4 ;
      RECT  18.0175 25.815 18.3625 31.38 ;
      RECT  94.315 1.38 94.5975 85.68 ;
      RECT  94.315 85.68 94.5975 86.095 ;
      RECT  94.315 86.095 94.5975 87.045 ;
      RECT  94.5975 1.38 94.73 85.68 ;
      RECT  94.5975 86.095 94.73 87.045 ;
      RECT  94.73 40.765 95.0125 85.68 ;
      RECT  94.73 86.095 95.0125 87.045 ;
      RECT  95.0125 40.765 96.6025 85.68 ;
      RECT  95.0125 85.68 96.6025 86.095 ;
      RECT  95.0125 86.095 96.6025 87.045 ;
      RECT  23.36 19.835 23.775 20.2075 ;
      RECT  23.36 20.2075 23.775 20.6225 ;
      RECT  23.36 20.6225 23.775 79.62 ;
      RECT  23.775 19.835 24.19 20.2075 ;
      RECT  23.775 20.6225 24.19 79.62 ;
      RECT  24.19 19.835 26.9575 20.2075 ;
      RECT  24.19 20.2075 26.9575 20.6225 ;
      RECT  24.19 20.6225 26.9575 79.62 ;
      RECT  96.6025 34.785 97.0175 37.36 ;
      RECT  96.6025 37.775 97.0175 40.35 ;
      RECT  28.1025 72.8575 31.2875 75.1275 ;
      RECT  31.2875 72.8575 31.7025 75.1275 ;
      RECT  31.7025 72.8575 45.5425 75.1275 ;
      RECT  45.5425 72.8575 45.9575 75.1275 ;
      RECT  45.9575 72.8575 79.3725 75.1275 ;
      RECT  79.3725 72.8575 83.4 75.1275 ;
      RECT  83.4 72.8575 84.5425 75.1275 ;
      RECT  83.4 75.1275 84.5425 75.4775 ;
      RECT  83.4 75.4775 84.5425 79.62 ;
      RECT  23.36 0.275 36.9625 0.965 ;
      RECT  36.9625 0.275 37.3775 0.965 ;
      RECT  37.3775 0.275 114.815 0.965 ;
      RECT  11.92 31.795 15.795 32.875 ;
      RECT  11.92 32.875 15.795 33.29 ;
      RECT  11.92 33.29 15.795 42.95 ;
      RECT  15.795 31.795 16.21 32.875 ;
      RECT  16.21 31.795 17.6025 32.875 ;
      RECT  16.21 32.875 17.6025 33.29 ;
      RECT  16.21 33.29 17.6025 42.95 ;
      RECT  37.3775 0.14 48.4025 0.275 ;
      RECT  48.8175 0.14 114.815 0.275 ;
      RECT  97.0175 20.225 97.785 26.895 ;
      RECT  97.0175 26.895 97.785 27.31 ;
      RECT  97.0175 27.31 97.785 40.35 ;
      RECT  97.785 27.31 98.2 40.35 ;
      RECT  98.2 20.225 102.895 26.895 ;
      RECT  98.2 26.895 102.895 27.31 ;
      RECT  79.3725 1.38 83.3675 14.4275 ;
      RECT  79.3725 14.7775 83.3675 17.0475 ;
      RECT  83.3675 1.38 83.4 14.4275 ;
      RECT  83.3675 14.7775 83.4 17.0475 ;
      RECT  83.4 1.38 90.43 14.4275 ;
      RECT  83.4 14.4275 90.43 14.7775 ;
      RECT  83.4 14.7775 90.43 17.0475 ;
      RECT  28.1025 14.7775 31.2875 17.0475 ;
      RECT  31.2875 14.7775 31.7025 17.0475 ;
      RECT  31.7025 14.7775 45.5425 17.0475 ;
      RECT  45.5425 14.7775 45.9575 17.0475 ;
      RECT  45.9575 14.7775 79.3725 17.0475 ;
      RECT  0.14 0.14 2.285 0.245 ;
      RECT  0.14 0.245 2.285 0.66 ;
      RECT  0.14 0.66 2.285 0.965 ;
      RECT  2.285 0.14 2.7 0.245 ;
      RECT  2.285 0.66 2.7 0.965 ;
      RECT  2.7 0.66 22.945 0.965 ;
      RECT  28.1025 8.7475 31.2875 10.4475 ;
      RECT  28.1025 10.7975 31.2875 14.4275 ;
      RECT  31.2875 8.7475 31.7025 10.4475 ;
      RECT  31.2875 10.7975 31.7025 14.4275 ;
      RECT  31.7025 8.7475 45.5425 10.4475 ;
      RECT  31.7025 10.7975 45.5425 14.4275 ;
      RECT  45.5425 8.7475 45.9575 10.4475 ;
      RECT  45.5425 10.7975 45.9575 14.4275 ;
      RECT  45.9575 8.7475 79.3725 10.4475 ;
      RECT  45.9575 10.7975 79.3725 14.4275 ;
      RECT  11.92 2.745 15.795 29.885 ;
      RECT  11.92 29.885 15.795 30.3 ;
      RECT  11.92 30.3 15.795 31.38 ;
      RECT  15.795 2.745 16.21 29.885 ;
      RECT  15.795 30.3 16.21 31.38 ;
      RECT  16.21 29.885 16.9425 30.3 ;
      RECT  16.21 30.3 16.9425 31.38 ;
      RECT  16.21 2.745 16.42 23.905 ;
      RECT  16.21 23.905 16.42 24.32 ;
      RECT  16.21 24.32 16.42 29.885 ;
      RECT  16.835 2.745 16.9425 23.905 ;
      RECT  16.835 23.905 16.9425 24.32 ;
      RECT  16.835 24.32 16.9425 29.885 ;
      RECT  28.1025 75.4775 31.2875 77.7275 ;
      RECT  28.1025 78.0775 31.2875 79.62 ;
      RECT  31.2875 75.4775 31.7025 77.7275 ;
      RECT  31.2875 78.0775 31.7025 79.62 ;
      RECT  31.7025 75.4775 45.5425 77.7275 ;
      RECT  31.7025 78.0775 45.5425 79.62 ;
      RECT  45.5425 75.4775 45.9575 77.7275 ;
      RECT  45.5425 78.0775 45.9575 79.62 ;
      RECT  45.9575 75.4775 79.3725 77.7275 ;
      RECT  45.9575 78.0775 79.3725 79.62 ;
      RECT  79.3725 75.4775 79.4075 77.7275 ;
      RECT  79.3725 78.0775 79.4075 79.62 ;
      RECT  79.4075 75.4775 83.4 77.7275 ;
      RECT  79.4075 77.7275 83.4 78.0775 ;
      RECT  79.4075 78.0775 83.4 79.62 ;
      RECT  23.36 0.14 25.5225 0.275 ;
      RECT  25.9375 0.14 36.9625 0.275 ;
      RECT  16.42 2.745 16.835 20.915 ;
      RECT  16.42 21.33 16.835 23.905 ;
      RECT  94.73 87.045 112.255 87.19 ;
      RECT  94.73 87.19 112.255 87.46 ;
      RECT  112.255 87.19 112.67 87.46 ;
      RECT  112.67 87.045 114.815 87.19 ;
      RECT  112.67 87.19 114.815 87.46 ;
      RECT  103.31 86.085 112.255 86.775 ;
      RECT  103.31 86.775 112.255 87.045 ;
      RECT  112.255 86.085 112.67 86.775 ;
      RECT  112.67 86.085 114.395 86.775 ;
      RECT  112.67 86.775 114.395 87.045 ;
      RECT  97.0175 40.765 98.41 41.845 ;
      RECT  97.0175 41.845 98.41 42.26 ;
      RECT  97.0175 42.26 98.41 87.045 ;
      RECT  98.41 40.765 98.825 41.845 ;
      RECT  98.41 42.26 98.825 87.045 ;
      RECT  98.825 40.765 102.895 41.845 ;
      RECT  98.825 41.845 102.895 42.26 ;
      RECT  98.825 42.26 102.895 87.045 ;
      RECT  98.2 27.31 98.41 35.865 ;
      RECT  98.2 35.865 98.41 36.28 ;
      RECT  98.2 36.28 98.41 40.35 ;
      RECT  98.825 27.31 102.895 35.865 ;
      RECT  98.825 35.865 102.895 36.28 ;
      RECT  98.825 36.28 102.895 40.35 ;
      RECT  2.7 0.14 19.8025 0.245 ;
      RECT  20.2175 0.14 22.945 0.245 ;
      RECT  2.7 0.245 19.8025 0.275 ;
      RECT  2.7 0.275 19.8025 0.66 ;
      RECT  19.8025 0.275 20.2175 0.66 ;
      RECT  20.2175 0.245 22.945 0.275 ;
      RECT  20.2175 0.275 22.945 0.66 ;
      RECT  98.41 36.28 98.825 38.855 ;
      RECT  98.41 39.27 98.825 40.35 ;
      RECT  97.785 20.225 98.2 20.915 ;
      RECT  15.795 33.29 16.21 35.865 ;
      RECT  15.795 36.28 16.21 38.855 ;
      RECT  16.42 24.32 16.835 26.895 ;
      RECT  16.42 27.31 16.835 29.885 ;
      RECT  23.36 87.46 91.7375 88.15 ;
      RECT  23.36 88.15 91.7375 88.285 ;
      RECT  91.7375 87.46 92.1525 88.15 ;
      RECT  92.1525 87.46 94.315 88.15 ;
      RECT  92.1525 88.15 94.315 88.285 ;
      RECT  15.795 39.27 16.21 41.845 ;
      RECT  15.795 42.26 16.21 42.95 ;
      RECT  98.41 27.31 98.825 29.885 ;
      RECT  97.785 21.33 98.2 23.905 ;
      RECT  97.785 24.32 98.2 26.895 ;
      RECT  98.41 30.3 98.825 32.875 ;
      RECT  98.41 33.29 98.825 35.865 ;
   LAYER  metal4 ;
      RECT  13.8 0.14 14.5 2.5725 ;
      RECT  14.5 0.14 114.815 2.5725 ;
      RECT  0.14 41.7025 11.08 54.8175 ;
      RECT  0.14 54.8175 11.08 88.285 ;
      RECT  11.08 18.0925 11.78 41.7025 ;
      RECT  11.08 54.8175 11.78 88.285 ;
      RECT  11.78 18.0925 13.8 41.7025 ;
      RECT  11.78 41.7025 13.8 54.8175 ;
      RECT  11.78 54.8175 13.8 88.285 ;
      RECT  21.17 2.5725 21.87 4.565 ;
      RECT  21.17 15.145 21.87 18.0925 ;
      RECT  21.87 2.5725 114.815 4.565 ;
      RECT  26.815 18.0925 27.515 20.7725 ;
      RECT  26.815 69.3125 27.515 88.285 ;
      RECT  0.14 2.5725 0.4075 9.95 ;
      RECT  0.14 9.95 0.4075 18.0925 ;
      RECT  0.4075 2.5725 1.1075 9.95 ;
      RECT  0.14 18.0925 0.4075 32.9125 ;
      RECT  0.14 32.9125 0.4075 41.7025 ;
      RECT  0.4075 32.9125 1.1075 41.7025 ;
      RECT  27.515 74.76 92.75 85.34 ;
      RECT  27.515 85.34 92.75 88.285 ;
      RECT  92.75 85.34 93.45 88.285 ;
      RECT  21.87 15.145 86.025 17.6025 ;
      RECT  86.025 15.145 86.725 17.6025 ;
      RECT  27.515 72.2325 86.025 74.76 ;
      RECT  86.025 72.2325 86.725 74.76 ;
      RECT  86.725 72.2325 92.75 74.76 ;
      RECT  93.45 69.3125 100.315 74.2825 ;
      RECT  100.315 69.3125 101.015 74.2825 ;
      RECT  100.315 84.8625 101.015 85.34 ;
      RECT  14.5 69.3825 23.015 88.285 ;
      RECT  23.015 69.3825 23.715 88.285 ;
      RECT  23.715 69.3825 26.815 88.285 ;
      RECT  21.87 17.6025 27.895 18.0925 ;
      RECT  27.515 18.0925 27.895 20.7725 ;
      RECT  27.515 20.7725 27.895 69.3125 ;
      RECT  27.515 69.3125 27.895 72.2325 ;
      RECT  113.8475 20.7725 114.5475 54.5225 ;
      RECT  114.5475 20.7725 114.815 54.5225 ;
      RECT  114.5475 54.5225 114.815 69.3125 ;
      RECT  114.5475 69.3125 114.815 74.2825 ;
      RECT  114.5475 74.2825 114.815 74.76 ;
      RECT  113.8475 77.485 114.5475 84.8625 ;
      RECT  114.5475 74.76 114.815 77.485 ;
      RECT  114.5475 77.485 114.815 84.8625 ;
      RECT  21.87 4.565 103.035 8.3575 ;
      RECT  103.035 4.565 103.735 8.3575 ;
      RECT  103.735 4.565 114.815 8.3575 ;
      RECT  103.735 8.3575 114.815 15.145 ;
      RECT  103.735 15.145 114.815 17.6025 ;
      RECT  103.735 17.6025 114.815 18.0925 ;
      RECT  103.735 18.0925 114.815 20.7725 ;
      RECT  103.035 21.4725 103.735 54.5225 ;
      RECT  103.735 20.7725 113.8475 21.4725 ;
      RECT  86.725 69.3825 90.905 72.2325 ;
      RECT  90.905 69.3825 91.605 72.2325 ;
      RECT  91.605 69.3825 92.75 72.2325 ;
      RECT  86.725 54.5225 87.105 69.3125 ;
      RECT  86.725 20.7725 87.105 21.4725 ;
      RECT  86.725 21.4725 87.105 54.5225 ;
      RECT  14.5 18.0925 21.425 20.74 ;
      RECT  14.5 20.74 21.425 20.7725 ;
      RECT  21.425 18.0925 22.125 20.74 ;
      RECT  22.125 18.0925 26.815 20.74 ;
      RECT  22.125 20.7725 23.015 69.3125 ;
      RECT  14.5 69.3125 21.425 69.3825 ;
      RECT  22.125 69.3125 23.015 69.3825 ;
      RECT  93.45 85.34 94.4125 85.4075 ;
      RECT  93.45 85.4075 94.4125 88.285 ;
      RECT  94.4125 85.4075 95.1125 88.285 ;
      RECT  93.45 74.2825 94.4125 74.6925 ;
      RECT  93.45 74.6925 94.4125 74.76 ;
      RECT  94.4125 74.2825 95.1125 74.6925 ;
      RECT  95.1125 74.2825 100.315 74.6925 ;
      RECT  95.1125 74.6925 100.315 74.76 ;
      RECT  93.45 74.76 94.4125 84.8625 ;
      RECT  95.1125 74.76 100.315 84.8625 ;
      RECT  93.45 84.8625 94.4125 85.34 ;
      RECT  95.1125 84.8625 100.315 85.34 ;
      RECT  13.8 18.0925 13.94 41.6375 ;
      RECT  13.8 41.6375 13.94 54.7525 ;
      RECT  13.8 54.7525 13.94 88.285 ;
      RECT  13.94 18.0925 14.5 41.6375 ;
      RECT  13.94 54.7525 14.5 88.285 ;
      RECT  14.5 20.7725 14.64 41.6375 ;
      RECT  14.5 54.7525 14.64 69.3125 ;
      RECT  14.64 20.7725 21.425 41.6375 ;
      RECT  14.64 41.6375 21.425 54.7525 ;
      RECT  14.64 54.7525 21.425 69.3125 ;
      RECT  92.75 69.3825 93.195 74.76 ;
      RECT  93.195 69.3125 93.45 69.3825 ;
      RECT  93.195 69.3825 93.45 74.76 ;
      RECT  86.725 18.0925 92.495 20.74 ;
      RECT  92.495 18.0925 93.195 20.74 ;
      RECT  91.605 69.3125 92.495 69.3825 ;
      RECT  91.605 54.5225 92.495 69.3125 ;
      RECT  91.605 20.7725 92.495 21.4725 ;
      RECT  91.605 21.4725 92.495 54.5225 ;
      RECT  1.1075 9.95 2.47 9.9825 ;
      RECT  1.1075 9.9825 2.47 18.0925 ;
      RECT  2.47 9.95 3.17 9.9825 ;
      RECT  1.1075 18.0925 2.47 32.9125 ;
      RECT  3.17 18.0925 11.08 32.9125 ;
      RECT  1.1075 32.9125 2.47 32.945 ;
      RECT  1.1075 32.945 2.47 41.7025 ;
      RECT  2.47 32.945 3.17 41.7025 ;
      RECT  3.17 32.9125 11.08 32.945 ;
      RECT  3.17 32.945 11.08 41.7025 ;
      RECT  112.485 69.3125 113.8475 74.2825 ;
      RECT  112.485 74.2825 113.8475 74.76 ;
      RECT  111.785 77.4525 112.485 77.485 ;
      RECT  112.485 74.76 113.8475 77.4525 ;
      RECT  112.485 77.4525 113.8475 77.485 ;
      RECT  103.735 21.4725 111.785 54.49 ;
      RECT  103.735 54.49 111.785 54.5225 ;
      RECT  111.785 21.4725 112.485 54.49 ;
      RECT  112.485 21.4725 113.8475 54.49 ;
      RECT  112.485 54.49 113.8475 54.5225 ;
      RECT  93.195 54.5225 111.785 69.3125 ;
      RECT  112.485 54.5225 113.8475 69.3125 ;
      RECT  21.87 8.3575 100.175 8.4225 ;
      RECT  21.87 8.4225 100.175 15.145 ;
      RECT  100.175 8.3575 100.875 8.4225 ;
      RECT  100.875 8.3575 103.035 8.4225 ;
      RECT  100.875 8.4225 103.035 15.145 ;
      RECT  86.725 15.145 100.175 17.6025 ;
      RECT  100.875 15.145 103.035 17.6025 ;
      RECT  86.725 17.6025 100.175 18.0925 ;
      RECT  100.875 17.6025 103.035 18.0925 ;
      RECT  93.195 18.0925 100.175 20.74 ;
      RECT  100.875 18.0925 103.035 20.74 ;
      RECT  93.195 20.74 100.175 20.7725 ;
      RECT  100.875 20.74 103.035 20.7725 ;
      RECT  93.195 20.7725 100.175 21.4725 ;
      RECT  100.875 20.7725 103.035 21.4725 ;
      RECT  93.195 21.4725 100.175 21.5375 ;
      RECT  93.195 21.5375 100.175 54.5225 ;
      RECT  100.175 21.5375 100.875 54.5225 ;
      RECT  100.875 21.4725 103.035 21.5375 ;
      RECT  100.875 21.5375 103.035 54.5225 ;
      RECT  24.275 20.7725 26.815 69.3125 ;
      RECT  23.715 69.345 24.275 69.3825 ;
      RECT  24.275 69.3125 26.815 69.345 ;
      RECT  24.275 69.345 26.815 69.3825 ;
      RECT  22.125 20.74 23.575 20.7725 ;
      RECT  24.275 20.74 26.815 20.7725 ;
      RECT  101.015 84.8625 108.29 85.34 ;
      RECT  108.99 84.8625 114.815 85.34 ;
      RECT  101.015 77.485 108.29 84.8625 ;
      RECT  108.99 77.485 113.8475 84.8625 ;
      RECT  95.1125 85.34 108.29 85.4075 ;
      RECT  108.99 85.34 114.815 85.4075 ;
      RECT  95.1125 85.4075 108.29 87.3325 ;
      RECT  95.1125 87.3325 108.29 88.285 ;
      RECT  108.29 87.3325 108.99 88.285 ;
      RECT  108.99 85.4075 114.815 87.3325 ;
      RECT  108.99 87.3325 114.815 88.285 ;
      RECT  101.015 69.3125 108.29 71.8125 ;
      RECT  101.015 71.8125 108.29 74.2825 ;
      RECT  108.29 69.3125 108.99 71.8125 ;
      RECT  108.99 69.3125 111.785 71.8125 ;
      RECT  108.99 71.8125 111.785 74.2825 ;
      RECT  101.015 74.2825 108.29 74.76 ;
      RECT  108.99 74.2825 111.785 74.76 ;
      RECT  101.015 74.76 108.29 77.4525 ;
      RECT  108.99 74.76 111.785 77.4525 ;
      RECT  101.015 77.4525 108.29 77.485 ;
      RECT  108.99 77.4525 111.785 77.485 ;
      RECT  14.5 2.5725 19.5075 4.4975 ;
      RECT  14.5 4.4975 19.5075 4.565 ;
      RECT  19.5075 2.5725 20.2075 4.4975 ;
      RECT  20.2075 2.5725 21.17 4.4975 ;
      RECT  20.2075 4.4975 21.17 4.565 ;
      RECT  14.5 4.565 19.5075 15.145 ;
      RECT  20.2075 4.565 21.17 15.145 ;
      RECT  14.5 15.145 19.5075 15.2125 ;
      RECT  14.5 15.2125 19.5075 18.0925 ;
      RECT  19.5075 15.2125 20.2075 18.0925 ;
      RECT  20.2075 15.145 21.17 15.2125 ;
      RECT  20.2075 15.2125 21.17 18.0925 ;
      RECT  86.725 69.3125 90.345 69.345 ;
      RECT  86.725 69.345 90.345 69.3825 ;
      RECT  90.345 69.345 90.905 69.3825 ;
      RECT  87.805 54.5225 90.345 69.3125 ;
      RECT  87.805 20.7725 90.345 21.4725 ;
      RECT  87.805 21.4725 90.345 54.5225 ;
      RECT  86.725 20.74 90.345 20.7725 ;
      RECT  91.045 20.74 92.495 20.7725 ;
      RECT  29.055 17.6025 85.565 18.0925 ;
      RECT  29.055 18.0925 85.565 20.7725 ;
      RECT  29.055 20.7725 85.565 69.3125 ;
      RECT  29.055 69.3125 85.565 72.2325 ;
      RECT  0.14 0.14 5.825 2.5725 ;
      RECT  6.525 0.14 13.8 2.5725 ;
      RECT  1.1075 2.5725 5.825 9.95 ;
      RECT  6.525 2.5725 13.8 9.95 ;
      RECT  3.17 9.95 5.825 9.9825 ;
      RECT  6.525 9.95 13.8 9.9825 ;
      RECT  3.17 9.9825 5.825 15.6225 ;
      RECT  3.17 15.6225 5.825 18.0925 ;
      RECT  5.825 15.6225 6.525 18.0925 ;
      RECT  6.525 9.9825 13.8 15.6225 ;
      RECT  6.525 15.6225 13.8 18.0925 ;
   END
END    freepdk45_sram_1w1r_11x128
END    LIBRARY
