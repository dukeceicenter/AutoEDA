../macros/freepdk45_sram_1rw0r_64x88_22/freepdk45_sram_1rw0r_64x88_22.lef