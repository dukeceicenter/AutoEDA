**************************************************
* OpenRAM generated memory.
* Words: 45
* Data bits: 512
* Banks: 1
* Column mux: 1:1
* Trimmed: False
* LVS: False
**************************************************
* File: DFFPOSX1.pex.netlist
* Created: Wed Jan  2 18:36:24 2008
* Program "Calibre xRC"
* Version "v2007.2_34.24"
*
.subckt dff D Q clk vdd gnd
*
MM21 Q a_66_6# gnd gnd NMOS_VTG L=5e-08 W=5e-07
MM19 a_76_6# a_2_6# a_66_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM20 gnd Q a_76_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM18 a_66_6# clk a_61_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM17 a_61_6# a_34_4# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM10 gnd clk a_2_6# gnd NMOS_VTG L=5e-08 W=5e-07
MM16 a_34_4# a_22_6# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM15 gnd a_34_4# a_31_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM14 a_31_6# clk a_22_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM13 a_22_6# a_2_6# a_17_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM12 a_17_6# D gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM11 Q a_66_6# vdd vdd PMOS_VTG L=5e-08 W=1e-06
MM9 vdd Q a_76_84# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM8 a_76_84# clk a_66_6# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM7 a_66_6# a_2_6# a_61_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM6 a_61_74# a_34_4# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM0 vdd clk a_2_6# vdd PMOS_VTG L=5e-08 W=1e-06
MM5 a_34_4# a_22_6# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM4 vdd a_34_4# a_31_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM3 a_31_74# a_2_6# a_22_6# vdd PMOS_VTG L=5e-08 W=5e-07
MM2 a_22_6# clk a_17_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM1 a_17_74# D vdd vdd PMOS_VTG L=5e-08 W=5e-07
* c_9 a_66_6# 0 0.271997f
* c_20 clk 0 0.350944f
* c_27 Q 0 0.202617f
* c_32 a_76_84# 0 0.0210573f
* c_38 a_76_6# 0 0.0204911f
* c_45 a_34_4# 0 0.172306f
* c_55 a_2_6# 0 0.283119f
* c_59 a_22_6# 0 0.157312f
* c_64 D 0 0.0816386f
* c_73 gnd 0 0.254131f
* c_81 vdd 0 0.23624f
*
*.include "dff.pex.netlist.dff.pxi"
*
.ends
*
*

.SUBCKT freepdk45_sram_1rw0r_45x512_row_addr_dff
+ din_0 din_1 din_2 din_3 din_4 din_5 dout_0 dout_1 dout_2 dout_3 dout_4
+ dout_5 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 6 cols: 1
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r1_c0
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r2_c0
+ din_2 dout_2 clk vdd gnd
+ dff
Xdff_r3_c0
+ din_3 dout_3 clk vdd gnd
+ dff
Xdff_r4_c0
+ din_4 dout_4 clk vdd gnd
+ dff
Xdff_r5_c0
+ din_5 dout_5 clk vdd gnd
+ dff
.ENDS freepdk45_sram_1rw0r_45x512_row_addr_dff

.SUBCKT freepdk45_sram_1rw0r_45x512_data_dff
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10
+ din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20
+ din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30
+ din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40
+ din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50
+ din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60
+ din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70
+ din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80
+ din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90
+ din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100
+ din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108
+ din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116
+ din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124
+ din_125 din_126 din_127 din_128 din_129 din_130 din_131 din_132
+ din_133 din_134 din_135 din_136 din_137 din_138 din_139 din_140
+ din_141 din_142 din_143 din_144 din_145 din_146 din_147 din_148
+ din_149 din_150 din_151 din_152 din_153 din_154 din_155 din_156
+ din_157 din_158 din_159 din_160 din_161 din_162 din_163 din_164
+ din_165 din_166 din_167 din_168 din_169 din_170 din_171 din_172
+ din_173 din_174 din_175 din_176 din_177 din_178 din_179 din_180
+ din_181 din_182 din_183 din_184 din_185 din_186 din_187 din_188
+ din_189 din_190 din_191 din_192 din_193 din_194 din_195 din_196
+ din_197 din_198 din_199 din_200 din_201 din_202 din_203 din_204
+ din_205 din_206 din_207 din_208 din_209 din_210 din_211 din_212
+ din_213 din_214 din_215 din_216 din_217 din_218 din_219 din_220
+ din_221 din_222 din_223 din_224 din_225 din_226 din_227 din_228
+ din_229 din_230 din_231 din_232 din_233 din_234 din_235 din_236
+ din_237 din_238 din_239 din_240 din_241 din_242 din_243 din_244
+ din_245 din_246 din_247 din_248 din_249 din_250 din_251 din_252
+ din_253 din_254 din_255 din_256 din_257 din_258 din_259 din_260
+ din_261 din_262 din_263 din_264 din_265 din_266 din_267 din_268
+ din_269 din_270 din_271 din_272 din_273 din_274 din_275 din_276
+ din_277 din_278 din_279 din_280 din_281 din_282 din_283 din_284
+ din_285 din_286 din_287 din_288 din_289 din_290 din_291 din_292
+ din_293 din_294 din_295 din_296 din_297 din_298 din_299 din_300
+ din_301 din_302 din_303 din_304 din_305 din_306 din_307 din_308
+ din_309 din_310 din_311 din_312 din_313 din_314 din_315 din_316
+ din_317 din_318 din_319 din_320 din_321 din_322 din_323 din_324
+ din_325 din_326 din_327 din_328 din_329 din_330 din_331 din_332
+ din_333 din_334 din_335 din_336 din_337 din_338 din_339 din_340
+ din_341 din_342 din_343 din_344 din_345 din_346 din_347 din_348
+ din_349 din_350 din_351 din_352 din_353 din_354 din_355 din_356
+ din_357 din_358 din_359 din_360 din_361 din_362 din_363 din_364
+ din_365 din_366 din_367 din_368 din_369 din_370 din_371 din_372
+ din_373 din_374 din_375 din_376 din_377 din_378 din_379 din_380
+ din_381 din_382 din_383 din_384 din_385 din_386 din_387 din_388
+ din_389 din_390 din_391 din_392 din_393 din_394 din_395 din_396
+ din_397 din_398 din_399 din_400 din_401 din_402 din_403 din_404
+ din_405 din_406 din_407 din_408 din_409 din_410 din_411 din_412
+ din_413 din_414 din_415 din_416 din_417 din_418 din_419 din_420
+ din_421 din_422 din_423 din_424 din_425 din_426 din_427 din_428
+ din_429 din_430 din_431 din_432 din_433 din_434 din_435 din_436
+ din_437 din_438 din_439 din_440 din_441 din_442 din_443 din_444
+ din_445 din_446 din_447 din_448 din_449 din_450 din_451 din_452
+ din_453 din_454 din_455 din_456 din_457 din_458 din_459 din_460
+ din_461 din_462 din_463 din_464 din_465 din_466 din_467 din_468
+ din_469 din_470 din_471 din_472 din_473 din_474 din_475 din_476
+ din_477 din_478 din_479 din_480 din_481 din_482 din_483 din_484
+ din_485 din_486 din_487 din_488 din_489 din_490 din_491 din_492
+ din_493 din_494 din_495 din_496 din_497 din_498 din_499 din_500
+ din_501 din_502 din_503 din_504 din_505 din_506 din_507 din_508
+ din_509 din_510 din_511 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5
+ dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14
+ dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22
+ dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30
+ dout_31 dout_32 dout_33 dout_34 dout_35 dout_36 dout_37 dout_38
+ dout_39 dout_40 dout_41 dout_42 dout_43 dout_44 dout_45 dout_46
+ dout_47 dout_48 dout_49 dout_50 dout_51 dout_52 dout_53 dout_54
+ dout_55 dout_56 dout_57 dout_58 dout_59 dout_60 dout_61 dout_62
+ dout_63 dout_64 dout_65 dout_66 dout_67 dout_68 dout_69 dout_70
+ dout_71 dout_72 dout_73 dout_74 dout_75 dout_76 dout_77 dout_78
+ dout_79 dout_80 dout_81 dout_82 dout_83 dout_84 dout_85 dout_86
+ dout_87 dout_88 dout_89 dout_90 dout_91 dout_92 dout_93 dout_94
+ dout_95 dout_96 dout_97 dout_98 dout_99 dout_100 dout_101 dout_102
+ dout_103 dout_104 dout_105 dout_106 dout_107 dout_108 dout_109
+ dout_110 dout_111 dout_112 dout_113 dout_114 dout_115 dout_116
+ dout_117 dout_118 dout_119 dout_120 dout_121 dout_122 dout_123
+ dout_124 dout_125 dout_126 dout_127 dout_128 dout_129 dout_130
+ dout_131 dout_132 dout_133 dout_134 dout_135 dout_136 dout_137
+ dout_138 dout_139 dout_140 dout_141 dout_142 dout_143 dout_144
+ dout_145 dout_146 dout_147 dout_148 dout_149 dout_150 dout_151
+ dout_152 dout_153 dout_154 dout_155 dout_156 dout_157 dout_158
+ dout_159 dout_160 dout_161 dout_162 dout_163 dout_164 dout_165
+ dout_166 dout_167 dout_168 dout_169 dout_170 dout_171 dout_172
+ dout_173 dout_174 dout_175 dout_176 dout_177 dout_178 dout_179
+ dout_180 dout_181 dout_182 dout_183 dout_184 dout_185 dout_186
+ dout_187 dout_188 dout_189 dout_190 dout_191 dout_192 dout_193
+ dout_194 dout_195 dout_196 dout_197 dout_198 dout_199 dout_200
+ dout_201 dout_202 dout_203 dout_204 dout_205 dout_206 dout_207
+ dout_208 dout_209 dout_210 dout_211 dout_212 dout_213 dout_214
+ dout_215 dout_216 dout_217 dout_218 dout_219 dout_220 dout_221
+ dout_222 dout_223 dout_224 dout_225 dout_226 dout_227 dout_228
+ dout_229 dout_230 dout_231 dout_232 dout_233 dout_234 dout_235
+ dout_236 dout_237 dout_238 dout_239 dout_240 dout_241 dout_242
+ dout_243 dout_244 dout_245 dout_246 dout_247 dout_248 dout_249
+ dout_250 dout_251 dout_252 dout_253 dout_254 dout_255 dout_256
+ dout_257 dout_258 dout_259 dout_260 dout_261 dout_262 dout_263
+ dout_264 dout_265 dout_266 dout_267 dout_268 dout_269 dout_270
+ dout_271 dout_272 dout_273 dout_274 dout_275 dout_276 dout_277
+ dout_278 dout_279 dout_280 dout_281 dout_282 dout_283 dout_284
+ dout_285 dout_286 dout_287 dout_288 dout_289 dout_290 dout_291
+ dout_292 dout_293 dout_294 dout_295 dout_296 dout_297 dout_298
+ dout_299 dout_300 dout_301 dout_302 dout_303 dout_304 dout_305
+ dout_306 dout_307 dout_308 dout_309 dout_310 dout_311 dout_312
+ dout_313 dout_314 dout_315 dout_316 dout_317 dout_318 dout_319
+ dout_320 dout_321 dout_322 dout_323 dout_324 dout_325 dout_326
+ dout_327 dout_328 dout_329 dout_330 dout_331 dout_332 dout_333
+ dout_334 dout_335 dout_336 dout_337 dout_338 dout_339 dout_340
+ dout_341 dout_342 dout_343 dout_344 dout_345 dout_346 dout_347
+ dout_348 dout_349 dout_350 dout_351 dout_352 dout_353 dout_354
+ dout_355 dout_356 dout_357 dout_358 dout_359 dout_360 dout_361
+ dout_362 dout_363 dout_364 dout_365 dout_366 dout_367 dout_368
+ dout_369 dout_370 dout_371 dout_372 dout_373 dout_374 dout_375
+ dout_376 dout_377 dout_378 dout_379 dout_380 dout_381 dout_382
+ dout_383 dout_384 dout_385 dout_386 dout_387 dout_388 dout_389
+ dout_390 dout_391 dout_392 dout_393 dout_394 dout_395 dout_396
+ dout_397 dout_398 dout_399 dout_400 dout_401 dout_402 dout_403
+ dout_404 dout_405 dout_406 dout_407 dout_408 dout_409 dout_410
+ dout_411 dout_412 dout_413 dout_414 dout_415 dout_416 dout_417
+ dout_418 dout_419 dout_420 dout_421 dout_422 dout_423 dout_424
+ dout_425 dout_426 dout_427 dout_428 dout_429 dout_430 dout_431
+ dout_432 dout_433 dout_434 dout_435 dout_436 dout_437 dout_438
+ dout_439 dout_440 dout_441 dout_442 dout_443 dout_444 dout_445
+ dout_446 dout_447 dout_448 dout_449 dout_450 dout_451 dout_452
+ dout_453 dout_454 dout_455 dout_456 dout_457 dout_458 dout_459
+ dout_460 dout_461 dout_462 dout_463 dout_464 dout_465 dout_466
+ dout_467 dout_468 dout_469 dout_470 dout_471 dout_472 dout_473
+ dout_474 dout_475 dout_476 dout_477 dout_478 dout_479 dout_480
+ dout_481 dout_482 dout_483 dout_484 dout_485 dout_486 dout_487
+ dout_488 dout_489 dout_490 dout_491 dout_492 dout_493 dout_494
+ dout_495 dout_496 dout_497 dout_498 dout_499 dout_500 dout_501
+ dout_502 dout_503 dout_504 dout_505 dout_506 dout_507 dout_508
+ dout_509 dout_510 dout_511 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : din_33 
* INPUT : din_34 
* INPUT : din_35 
* INPUT : din_36 
* INPUT : din_37 
* INPUT : din_38 
* INPUT : din_39 
* INPUT : din_40 
* INPUT : din_41 
* INPUT : din_42 
* INPUT : din_43 
* INPUT : din_44 
* INPUT : din_45 
* INPUT : din_46 
* INPUT : din_47 
* INPUT : din_48 
* INPUT : din_49 
* INPUT : din_50 
* INPUT : din_51 
* INPUT : din_52 
* INPUT : din_53 
* INPUT : din_54 
* INPUT : din_55 
* INPUT : din_56 
* INPUT : din_57 
* INPUT : din_58 
* INPUT : din_59 
* INPUT : din_60 
* INPUT : din_61 
* INPUT : din_62 
* INPUT : din_63 
* INPUT : din_64 
* INPUT : din_65 
* INPUT : din_66 
* INPUT : din_67 
* INPUT : din_68 
* INPUT : din_69 
* INPUT : din_70 
* INPUT : din_71 
* INPUT : din_72 
* INPUT : din_73 
* INPUT : din_74 
* INPUT : din_75 
* INPUT : din_76 
* INPUT : din_77 
* INPUT : din_78 
* INPUT : din_79 
* INPUT : din_80 
* INPUT : din_81 
* INPUT : din_82 
* INPUT : din_83 
* INPUT : din_84 
* INPUT : din_85 
* INPUT : din_86 
* INPUT : din_87 
* INPUT : din_88 
* INPUT : din_89 
* INPUT : din_90 
* INPUT : din_91 
* INPUT : din_92 
* INPUT : din_93 
* INPUT : din_94 
* INPUT : din_95 
* INPUT : din_96 
* INPUT : din_97 
* INPUT : din_98 
* INPUT : din_99 
* INPUT : din_100 
* INPUT : din_101 
* INPUT : din_102 
* INPUT : din_103 
* INPUT : din_104 
* INPUT : din_105 
* INPUT : din_106 
* INPUT : din_107 
* INPUT : din_108 
* INPUT : din_109 
* INPUT : din_110 
* INPUT : din_111 
* INPUT : din_112 
* INPUT : din_113 
* INPUT : din_114 
* INPUT : din_115 
* INPUT : din_116 
* INPUT : din_117 
* INPUT : din_118 
* INPUT : din_119 
* INPUT : din_120 
* INPUT : din_121 
* INPUT : din_122 
* INPUT : din_123 
* INPUT : din_124 
* INPUT : din_125 
* INPUT : din_126 
* INPUT : din_127 
* INPUT : din_128 
* INPUT : din_129 
* INPUT : din_130 
* INPUT : din_131 
* INPUT : din_132 
* INPUT : din_133 
* INPUT : din_134 
* INPUT : din_135 
* INPUT : din_136 
* INPUT : din_137 
* INPUT : din_138 
* INPUT : din_139 
* INPUT : din_140 
* INPUT : din_141 
* INPUT : din_142 
* INPUT : din_143 
* INPUT : din_144 
* INPUT : din_145 
* INPUT : din_146 
* INPUT : din_147 
* INPUT : din_148 
* INPUT : din_149 
* INPUT : din_150 
* INPUT : din_151 
* INPUT : din_152 
* INPUT : din_153 
* INPUT : din_154 
* INPUT : din_155 
* INPUT : din_156 
* INPUT : din_157 
* INPUT : din_158 
* INPUT : din_159 
* INPUT : din_160 
* INPUT : din_161 
* INPUT : din_162 
* INPUT : din_163 
* INPUT : din_164 
* INPUT : din_165 
* INPUT : din_166 
* INPUT : din_167 
* INPUT : din_168 
* INPUT : din_169 
* INPUT : din_170 
* INPUT : din_171 
* INPUT : din_172 
* INPUT : din_173 
* INPUT : din_174 
* INPUT : din_175 
* INPUT : din_176 
* INPUT : din_177 
* INPUT : din_178 
* INPUT : din_179 
* INPUT : din_180 
* INPUT : din_181 
* INPUT : din_182 
* INPUT : din_183 
* INPUT : din_184 
* INPUT : din_185 
* INPUT : din_186 
* INPUT : din_187 
* INPUT : din_188 
* INPUT : din_189 
* INPUT : din_190 
* INPUT : din_191 
* INPUT : din_192 
* INPUT : din_193 
* INPUT : din_194 
* INPUT : din_195 
* INPUT : din_196 
* INPUT : din_197 
* INPUT : din_198 
* INPUT : din_199 
* INPUT : din_200 
* INPUT : din_201 
* INPUT : din_202 
* INPUT : din_203 
* INPUT : din_204 
* INPUT : din_205 
* INPUT : din_206 
* INPUT : din_207 
* INPUT : din_208 
* INPUT : din_209 
* INPUT : din_210 
* INPUT : din_211 
* INPUT : din_212 
* INPUT : din_213 
* INPUT : din_214 
* INPUT : din_215 
* INPUT : din_216 
* INPUT : din_217 
* INPUT : din_218 
* INPUT : din_219 
* INPUT : din_220 
* INPUT : din_221 
* INPUT : din_222 
* INPUT : din_223 
* INPUT : din_224 
* INPUT : din_225 
* INPUT : din_226 
* INPUT : din_227 
* INPUT : din_228 
* INPUT : din_229 
* INPUT : din_230 
* INPUT : din_231 
* INPUT : din_232 
* INPUT : din_233 
* INPUT : din_234 
* INPUT : din_235 
* INPUT : din_236 
* INPUT : din_237 
* INPUT : din_238 
* INPUT : din_239 
* INPUT : din_240 
* INPUT : din_241 
* INPUT : din_242 
* INPUT : din_243 
* INPUT : din_244 
* INPUT : din_245 
* INPUT : din_246 
* INPUT : din_247 
* INPUT : din_248 
* INPUT : din_249 
* INPUT : din_250 
* INPUT : din_251 
* INPUT : din_252 
* INPUT : din_253 
* INPUT : din_254 
* INPUT : din_255 
* INPUT : din_256 
* INPUT : din_257 
* INPUT : din_258 
* INPUT : din_259 
* INPUT : din_260 
* INPUT : din_261 
* INPUT : din_262 
* INPUT : din_263 
* INPUT : din_264 
* INPUT : din_265 
* INPUT : din_266 
* INPUT : din_267 
* INPUT : din_268 
* INPUT : din_269 
* INPUT : din_270 
* INPUT : din_271 
* INPUT : din_272 
* INPUT : din_273 
* INPUT : din_274 
* INPUT : din_275 
* INPUT : din_276 
* INPUT : din_277 
* INPUT : din_278 
* INPUT : din_279 
* INPUT : din_280 
* INPUT : din_281 
* INPUT : din_282 
* INPUT : din_283 
* INPUT : din_284 
* INPUT : din_285 
* INPUT : din_286 
* INPUT : din_287 
* INPUT : din_288 
* INPUT : din_289 
* INPUT : din_290 
* INPUT : din_291 
* INPUT : din_292 
* INPUT : din_293 
* INPUT : din_294 
* INPUT : din_295 
* INPUT : din_296 
* INPUT : din_297 
* INPUT : din_298 
* INPUT : din_299 
* INPUT : din_300 
* INPUT : din_301 
* INPUT : din_302 
* INPUT : din_303 
* INPUT : din_304 
* INPUT : din_305 
* INPUT : din_306 
* INPUT : din_307 
* INPUT : din_308 
* INPUT : din_309 
* INPUT : din_310 
* INPUT : din_311 
* INPUT : din_312 
* INPUT : din_313 
* INPUT : din_314 
* INPUT : din_315 
* INPUT : din_316 
* INPUT : din_317 
* INPUT : din_318 
* INPUT : din_319 
* INPUT : din_320 
* INPUT : din_321 
* INPUT : din_322 
* INPUT : din_323 
* INPUT : din_324 
* INPUT : din_325 
* INPUT : din_326 
* INPUT : din_327 
* INPUT : din_328 
* INPUT : din_329 
* INPUT : din_330 
* INPUT : din_331 
* INPUT : din_332 
* INPUT : din_333 
* INPUT : din_334 
* INPUT : din_335 
* INPUT : din_336 
* INPUT : din_337 
* INPUT : din_338 
* INPUT : din_339 
* INPUT : din_340 
* INPUT : din_341 
* INPUT : din_342 
* INPUT : din_343 
* INPUT : din_344 
* INPUT : din_345 
* INPUT : din_346 
* INPUT : din_347 
* INPUT : din_348 
* INPUT : din_349 
* INPUT : din_350 
* INPUT : din_351 
* INPUT : din_352 
* INPUT : din_353 
* INPUT : din_354 
* INPUT : din_355 
* INPUT : din_356 
* INPUT : din_357 
* INPUT : din_358 
* INPUT : din_359 
* INPUT : din_360 
* INPUT : din_361 
* INPUT : din_362 
* INPUT : din_363 
* INPUT : din_364 
* INPUT : din_365 
* INPUT : din_366 
* INPUT : din_367 
* INPUT : din_368 
* INPUT : din_369 
* INPUT : din_370 
* INPUT : din_371 
* INPUT : din_372 
* INPUT : din_373 
* INPUT : din_374 
* INPUT : din_375 
* INPUT : din_376 
* INPUT : din_377 
* INPUT : din_378 
* INPUT : din_379 
* INPUT : din_380 
* INPUT : din_381 
* INPUT : din_382 
* INPUT : din_383 
* INPUT : din_384 
* INPUT : din_385 
* INPUT : din_386 
* INPUT : din_387 
* INPUT : din_388 
* INPUT : din_389 
* INPUT : din_390 
* INPUT : din_391 
* INPUT : din_392 
* INPUT : din_393 
* INPUT : din_394 
* INPUT : din_395 
* INPUT : din_396 
* INPUT : din_397 
* INPUT : din_398 
* INPUT : din_399 
* INPUT : din_400 
* INPUT : din_401 
* INPUT : din_402 
* INPUT : din_403 
* INPUT : din_404 
* INPUT : din_405 
* INPUT : din_406 
* INPUT : din_407 
* INPUT : din_408 
* INPUT : din_409 
* INPUT : din_410 
* INPUT : din_411 
* INPUT : din_412 
* INPUT : din_413 
* INPUT : din_414 
* INPUT : din_415 
* INPUT : din_416 
* INPUT : din_417 
* INPUT : din_418 
* INPUT : din_419 
* INPUT : din_420 
* INPUT : din_421 
* INPUT : din_422 
* INPUT : din_423 
* INPUT : din_424 
* INPUT : din_425 
* INPUT : din_426 
* INPUT : din_427 
* INPUT : din_428 
* INPUT : din_429 
* INPUT : din_430 
* INPUT : din_431 
* INPUT : din_432 
* INPUT : din_433 
* INPUT : din_434 
* INPUT : din_435 
* INPUT : din_436 
* INPUT : din_437 
* INPUT : din_438 
* INPUT : din_439 
* INPUT : din_440 
* INPUT : din_441 
* INPUT : din_442 
* INPUT : din_443 
* INPUT : din_444 
* INPUT : din_445 
* INPUT : din_446 
* INPUT : din_447 
* INPUT : din_448 
* INPUT : din_449 
* INPUT : din_450 
* INPUT : din_451 
* INPUT : din_452 
* INPUT : din_453 
* INPUT : din_454 
* INPUT : din_455 
* INPUT : din_456 
* INPUT : din_457 
* INPUT : din_458 
* INPUT : din_459 
* INPUT : din_460 
* INPUT : din_461 
* INPUT : din_462 
* INPUT : din_463 
* INPUT : din_464 
* INPUT : din_465 
* INPUT : din_466 
* INPUT : din_467 
* INPUT : din_468 
* INPUT : din_469 
* INPUT : din_470 
* INPUT : din_471 
* INPUT : din_472 
* INPUT : din_473 
* INPUT : din_474 
* INPUT : din_475 
* INPUT : din_476 
* INPUT : din_477 
* INPUT : din_478 
* INPUT : din_479 
* INPUT : din_480 
* INPUT : din_481 
* INPUT : din_482 
* INPUT : din_483 
* INPUT : din_484 
* INPUT : din_485 
* INPUT : din_486 
* INPUT : din_487 
* INPUT : din_488 
* INPUT : din_489 
* INPUT : din_490 
* INPUT : din_491 
* INPUT : din_492 
* INPUT : din_493 
* INPUT : din_494 
* INPUT : din_495 
* INPUT : din_496 
* INPUT : din_497 
* INPUT : din_498 
* INPUT : din_499 
* INPUT : din_500 
* INPUT : din_501 
* INPUT : din_502 
* INPUT : din_503 
* INPUT : din_504 
* INPUT : din_505 
* INPUT : din_506 
* INPUT : din_507 
* INPUT : din_508 
* INPUT : din_509 
* INPUT : din_510 
* INPUT : din_511 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* OUTPUT: dout_33 
* OUTPUT: dout_34 
* OUTPUT: dout_35 
* OUTPUT: dout_36 
* OUTPUT: dout_37 
* OUTPUT: dout_38 
* OUTPUT: dout_39 
* OUTPUT: dout_40 
* OUTPUT: dout_41 
* OUTPUT: dout_42 
* OUTPUT: dout_43 
* OUTPUT: dout_44 
* OUTPUT: dout_45 
* OUTPUT: dout_46 
* OUTPUT: dout_47 
* OUTPUT: dout_48 
* OUTPUT: dout_49 
* OUTPUT: dout_50 
* OUTPUT: dout_51 
* OUTPUT: dout_52 
* OUTPUT: dout_53 
* OUTPUT: dout_54 
* OUTPUT: dout_55 
* OUTPUT: dout_56 
* OUTPUT: dout_57 
* OUTPUT: dout_58 
* OUTPUT: dout_59 
* OUTPUT: dout_60 
* OUTPUT: dout_61 
* OUTPUT: dout_62 
* OUTPUT: dout_63 
* OUTPUT: dout_64 
* OUTPUT: dout_65 
* OUTPUT: dout_66 
* OUTPUT: dout_67 
* OUTPUT: dout_68 
* OUTPUT: dout_69 
* OUTPUT: dout_70 
* OUTPUT: dout_71 
* OUTPUT: dout_72 
* OUTPUT: dout_73 
* OUTPUT: dout_74 
* OUTPUT: dout_75 
* OUTPUT: dout_76 
* OUTPUT: dout_77 
* OUTPUT: dout_78 
* OUTPUT: dout_79 
* OUTPUT: dout_80 
* OUTPUT: dout_81 
* OUTPUT: dout_82 
* OUTPUT: dout_83 
* OUTPUT: dout_84 
* OUTPUT: dout_85 
* OUTPUT: dout_86 
* OUTPUT: dout_87 
* OUTPUT: dout_88 
* OUTPUT: dout_89 
* OUTPUT: dout_90 
* OUTPUT: dout_91 
* OUTPUT: dout_92 
* OUTPUT: dout_93 
* OUTPUT: dout_94 
* OUTPUT: dout_95 
* OUTPUT: dout_96 
* OUTPUT: dout_97 
* OUTPUT: dout_98 
* OUTPUT: dout_99 
* OUTPUT: dout_100 
* OUTPUT: dout_101 
* OUTPUT: dout_102 
* OUTPUT: dout_103 
* OUTPUT: dout_104 
* OUTPUT: dout_105 
* OUTPUT: dout_106 
* OUTPUT: dout_107 
* OUTPUT: dout_108 
* OUTPUT: dout_109 
* OUTPUT: dout_110 
* OUTPUT: dout_111 
* OUTPUT: dout_112 
* OUTPUT: dout_113 
* OUTPUT: dout_114 
* OUTPUT: dout_115 
* OUTPUT: dout_116 
* OUTPUT: dout_117 
* OUTPUT: dout_118 
* OUTPUT: dout_119 
* OUTPUT: dout_120 
* OUTPUT: dout_121 
* OUTPUT: dout_122 
* OUTPUT: dout_123 
* OUTPUT: dout_124 
* OUTPUT: dout_125 
* OUTPUT: dout_126 
* OUTPUT: dout_127 
* OUTPUT: dout_128 
* OUTPUT: dout_129 
* OUTPUT: dout_130 
* OUTPUT: dout_131 
* OUTPUT: dout_132 
* OUTPUT: dout_133 
* OUTPUT: dout_134 
* OUTPUT: dout_135 
* OUTPUT: dout_136 
* OUTPUT: dout_137 
* OUTPUT: dout_138 
* OUTPUT: dout_139 
* OUTPUT: dout_140 
* OUTPUT: dout_141 
* OUTPUT: dout_142 
* OUTPUT: dout_143 
* OUTPUT: dout_144 
* OUTPUT: dout_145 
* OUTPUT: dout_146 
* OUTPUT: dout_147 
* OUTPUT: dout_148 
* OUTPUT: dout_149 
* OUTPUT: dout_150 
* OUTPUT: dout_151 
* OUTPUT: dout_152 
* OUTPUT: dout_153 
* OUTPUT: dout_154 
* OUTPUT: dout_155 
* OUTPUT: dout_156 
* OUTPUT: dout_157 
* OUTPUT: dout_158 
* OUTPUT: dout_159 
* OUTPUT: dout_160 
* OUTPUT: dout_161 
* OUTPUT: dout_162 
* OUTPUT: dout_163 
* OUTPUT: dout_164 
* OUTPUT: dout_165 
* OUTPUT: dout_166 
* OUTPUT: dout_167 
* OUTPUT: dout_168 
* OUTPUT: dout_169 
* OUTPUT: dout_170 
* OUTPUT: dout_171 
* OUTPUT: dout_172 
* OUTPUT: dout_173 
* OUTPUT: dout_174 
* OUTPUT: dout_175 
* OUTPUT: dout_176 
* OUTPUT: dout_177 
* OUTPUT: dout_178 
* OUTPUT: dout_179 
* OUTPUT: dout_180 
* OUTPUT: dout_181 
* OUTPUT: dout_182 
* OUTPUT: dout_183 
* OUTPUT: dout_184 
* OUTPUT: dout_185 
* OUTPUT: dout_186 
* OUTPUT: dout_187 
* OUTPUT: dout_188 
* OUTPUT: dout_189 
* OUTPUT: dout_190 
* OUTPUT: dout_191 
* OUTPUT: dout_192 
* OUTPUT: dout_193 
* OUTPUT: dout_194 
* OUTPUT: dout_195 
* OUTPUT: dout_196 
* OUTPUT: dout_197 
* OUTPUT: dout_198 
* OUTPUT: dout_199 
* OUTPUT: dout_200 
* OUTPUT: dout_201 
* OUTPUT: dout_202 
* OUTPUT: dout_203 
* OUTPUT: dout_204 
* OUTPUT: dout_205 
* OUTPUT: dout_206 
* OUTPUT: dout_207 
* OUTPUT: dout_208 
* OUTPUT: dout_209 
* OUTPUT: dout_210 
* OUTPUT: dout_211 
* OUTPUT: dout_212 
* OUTPUT: dout_213 
* OUTPUT: dout_214 
* OUTPUT: dout_215 
* OUTPUT: dout_216 
* OUTPUT: dout_217 
* OUTPUT: dout_218 
* OUTPUT: dout_219 
* OUTPUT: dout_220 
* OUTPUT: dout_221 
* OUTPUT: dout_222 
* OUTPUT: dout_223 
* OUTPUT: dout_224 
* OUTPUT: dout_225 
* OUTPUT: dout_226 
* OUTPUT: dout_227 
* OUTPUT: dout_228 
* OUTPUT: dout_229 
* OUTPUT: dout_230 
* OUTPUT: dout_231 
* OUTPUT: dout_232 
* OUTPUT: dout_233 
* OUTPUT: dout_234 
* OUTPUT: dout_235 
* OUTPUT: dout_236 
* OUTPUT: dout_237 
* OUTPUT: dout_238 
* OUTPUT: dout_239 
* OUTPUT: dout_240 
* OUTPUT: dout_241 
* OUTPUT: dout_242 
* OUTPUT: dout_243 
* OUTPUT: dout_244 
* OUTPUT: dout_245 
* OUTPUT: dout_246 
* OUTPUT: dout_247 
* OUTPUT: dout_248 
* OUTPUT: dout_249 
* OUTPUT: dout_250 
* OUTPUT: dout_251 
* OUTPUT: dout_252 
* OUTPUT: dout_253 
* OUTPUT: dout_254 
* OUTPUT: dout_255 
* OUTPUT: dout_256 
* OUTPUT: dout_257 
* OUTPUT: dout_258 
* OUTPUT: dout_259 
* OUTPUT: dout_260 
* OUTPUT: dout_261 
* OUTPUT: dout_262 
* OUTPUT: dout_263 
* OUTPUT: dout_264 
* OUTPUT: dout_265 
* OUTPUT: dout_266 
* OUTPUT: dout_267 
* OUTPUT: dout_268 
* OUTPUT: dout_269 
* OUTPUT: dout_270 
* OUTPUT: dout_271 
* OUTPUT: dout_272 
* OUTPUT: dout_273 
* OUTPUT: dout_274 
* OUTPUT: dout_275 
* OUTPUT: dout_276 
* OUTPUT: dout_277 
* OUTPUT: dout_278 
* OUTPUT: dout_279 
* OUTPUT: dout_280 
* OUTPUT: dout_281 
* OUTPUT: dout_282 
* OUTPUT: dout_283 
* OUTPUT: dout_284 
* OUTPUT: dout_285 
* OUTPUT: dout_286 
* OUTPUT: dout_287 
* OUTPUT: dout_288 
* OUTPUT: dout_289 
* OUTPUT: dout_290 
* OUTPUT: dout_291 
* OUTPUT: dout_292 
* OUTPUT: dout_293 
* OUTPUT: dout_294 
* OUTPUT: dout_295 
* OUTPUT: dout_296 
* OUTPUT: dout_297 
* OUTPUT: dout_298 
* OUTPUT: dout_299 
* OUTPUT: dout_300 
* OUTPUT: dout_301 
* OUTPUT: dout_302 
* OUTPUT: dout_303 
* OUTPUT: dout_304 
* OUTPUT: dout_305 
* OUTPUT: dout_306 
* OUTPUT: dout_307 
* OUTPUT: dout_308 
* OUTPUT: dout_309 
* OUTPUT: dout_310 
* OUTPUT: dout_311 
* OUTPUT: dout_312 
* OUTPUT: dout_313 
* OUTPUT: dout_314 
* OUTPUT: dout_315 
* OUTPUT: dout_316 
* OUTPUT: dout_317 
* OUTPUT: dout_318 
* OUTPUT: dout_319 
* OUTPUT: dout_320 
* OUTPUT: dout_321 
* OUTPUT: dout_322 
* OUTPUT: dout_323 
* OUTPUT: dout_324 
* OUTPUT: dout_325 
* OUTPUT: dout_326 
* OUTPUT: dout_327 
* OUTPUT: dout_328 
* OUTPUT: dout_329 
* OUTPUT: dout_330 
* OUTPUT: dout_331 
* OUTPUT: dout_332 
* OUTPUT: dout_333 
* OUTPUT: dout_334 
* OUTPUT: dout_335 
* OUTPUT: dout_336 
* OUTPUT: dout_337 
* OUTPUT: dout_338 
* OUTPUT: dout_339 
* OUTPUT: dout_340 
* OUTPUT: dout_341 
* OUTPUT: dout_342 
* OUTPUT: dout_343 
* OUTPUT: dout_344 
* OUTPUT: dout_345 
* OUTPUT: dout_346 
* OUTPUT: dout_347 
* OUTPUT: dout_348 
* OUTPUT: dout_349 
* OUTPUT: dout_350 
* OUTPUT: dout_351 
* OUTPUT: dout_352 
* OUTPUT: dout_353 
* OUTPUT: dout_354 
* OUTPUT: dout_355 
* OUTPUT: dout_356 
* OUTPUT: dout_357 
* OUTPUT: dout_358 
* OUTPUT: dout_359 
* OUTPUT: dout_360 
* OUTPUT: dout_361 
* OUTPUT: dout_362 
* OUTPUT: dout_363 
* OUTPUT: dout_364 
* OUTPUT: dout_365 
* OUTPUT: dout_366 
* OUTPUT: dout_367 
* OUTPUT: dout_368 
* OUTPUT: dout_369 
* OUTPUT: dout_370 
* OUTPUT: dout_371 
* OUTPUT: dout_372 
* OUTPUT: dout_373 
* OUTPUT: dout_374 
* OUTPUT: dout_375 
* OUTPUT: dout_376 
* OUTPUT: dout_377 
* OUTPUT: dout_378 
* OUTPUT: dout_379 
* OUTPUT: dout_380 
* OUTPUT: dout_381 
* OUTPUT: dout_382 
* OUTPUT: dout_383 
* OUTPUT: dout_384 
* OUTPUT: dout_385 
* OUTPUT: dout_386 
* OUTPUT: dout_387 
* OUTPUT: dout_388 
* OUTPUT: dout_389 
* OUTPUT: dout_390 
* OUTPUT: dout_391 
* OUTPUT: dout_392 
* OUTPUT: dout_393 
* OUTPUT: dout_394 
* OUTPUT: dout_395 
* OUTPUT: dout_396 
* OUTPUT: dout_397 
* OUTPUT: dout_398 
* OUTPUT: dout_399 
* OUTPUT: dout_400 
* OUTPUT: dout_401 
* OUTPUT: dout_402 
* OUTPUT: dout_403 
* OUTPUT: dout_404 
* OUTPUT: dout_405 
* OUTPUT: dout_406 
* OUTPUT: dout_407 
* OUTPUT: dout_408 
* OUTPUT: dout_409 
* OUTPUT: dout_410 
* OUTPUT: dout_411 
* OUTPUT: dout_412 
* OUTPUT: dout_413 
* OUTPUT: dout_414 
* OUTPUT: dout_415 
* OUTPUT: dout_416 
* OUTPUT: dout_417 
* OUTPUT: dout_418 
* OUTPUT: dout_419 
* OUTPUT: dout_420 
* OUTPUT: dout_421 
* OUTPUT: dout_422 
* OUTPUT: dout_423 
* OUTPUT: dout_424 
* OUTPUT: dout_425 
* OUTPUT: dout_426 
* OUTPUT: dout_427 
* OUTPUT: dout_428 
* OUTPUT: dout_429 
* OUTPUT: dout_430 
* OUTPUT: dout_431 
* OUTPUT: dout_432 
* OUTPUT: dout_433 
* OUTPUT: dout_434 
* OUTPUT: dout_435 
* OUTPUT: dout_436 
* OUTPUT: dout_437 
* OUTPUT: dout_438 
* OUTPUT: dout_439 
* OUTPUT: dout_440 
* OUTPUT: dout_441 
* OUTPUT: dout_442 
* OUTPUT: dout_443 
* OUTPUT: dout_444 
* OUTPUT: dout_445 
* OUTPUT: dout_446 
* OUTPUT: dout_447 
* OUTPUT: dout_448 
* OUTPUT: dout_449 
* OUTPUT: dout_450 
* OUTPUT: dout_451 
* OUTPUT: dout_452 
* OUTPUT: dout_453 
* OUTPUT: dout_454 
* OUTPUT: dout_455 
* OUTPUT: dout_456 
* OUTPUT: dout_457 
* OUTPUT: dout_458 
* OUTPUT: dout_459 
* OUTPUT: dout_460 
* OUTPUT: dout_461 
* OUTPUT: dout_462 
* OUTPUT: dout_463 
* OUTPUT: dout_464 
* OUTPUT: dout_465 
* OUTPUT: dout_466 
* OUTPUT: dout_467 
* OUTPUT: dout_468 
* OUTPUT: dout_469 
* OUTPUT: dout_470 
* OUTPUT: dout_471 
* OUTPUT: dout_472 
* OUTPUT: dout_473 
* OUTPUT: dout_474 
* OUTPUT: dout_475 
* OUTPUT: dout_476 
* OUTPUT: dout_477 
* OUTPUT: dout_478 
* OUTPUT: dout_479 
* OUTPUT: dout_480 
* OUTPUT: dout_481 
* OUTPUT: dout_482 
* OUTPUT: dout_483 
* OUTPUT: dout_484 
* OUTPUT: dout_485 
* OUTPUT: dout_486 
* OUTPUT: dout_487 
* OUTPUT: dout_488 
* OUTPUT: dout_489 
* OUTPUT: dout_490 
* OUTPUT: dout_491 
* OUTPUT: dout_492 
* OUTPUT: dout_493 
* OUTPUT: dout_494 
* OUTPUT: dout_495 
* OUTPUT: dout_496 
* OUTPUT: dout_497 
* OUTPUT: dout_498 
* OUTPUT: dout_499 
* OUTPUT: dout_500 
* OUTPUT: dout_501 
* OUTPUT: dout_502 
* OUTPUT: dout_503 
* OUTPUT: dout_504 
* OUTPUT: dout_505 
* OUTPUT: dout_506 
* OUTPUT: dout_507 
* OUTPUT: dout_508 
* OUTPUT: dout_509 
* OUTPUT: dout_510 
* OUTPUT: dout_511 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 512
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r0_c1
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r0_c2
+ din_2 dout_2 clk vdd gnd
+ dff
Xdff_r0_c3
+ din_3 dout_3 clk vdd gnd
+ dff
Xdff_r0_c4
+ din_4 dout_4 clk vdd gnd
+ dff
Xdff_r0_c5
+ din_5 dout_5 clk vdd gnd
+ dff
Xdff_r0_c6
+ din_6 dout_6 clk vdd gnd
+ dff
Xdff_r0_c7
+ din_7 dout_7 clk vdd gnd
+ dff
Xdff_r0_c8
+ din_8 dout_8 clk vdd gnd
+ dff
Xdff_r0_c9
+ din_9 dout_9 clk vdd gnd
+ dff
Xdff_r0_c10
+ din_10 dout_10 clk vdd gnd
+ dff
Xdff_r0_c11
+ din_11 dout_11 clk vdd gnd
+ dff
Xdff_r0_c12
+ din_12 dout_12 clk vdd gnd
+ dff
Xdff_r0_c13
+ din_13 dout_13 clk vdd gnd
+ dff
Xdff_r0_c14
+ din_14 dout_14 clk vdd gnd
+ dff
Xdff_r0_c15
+ din_15 dout_15 clk vdd gnd
+ dff
Xdff_r0_c16
+ din_16 dout_16 clk vdd gnd
+ dff
Xdff_r0_c17
+ din_17 dout_17 clk vdd gnd
+ dff
Xdff_r0_c18
+ din_18 dout_18 clk vdd gnd
+ dff
Xdff_r0_c19
+ din_19 dout_19 clk vdd gnd
+ dff
Xdff_r0_c20
+ din_20 dout_20 clk vdd gnd
+ dff
Xdff_r0_c21
+ din_21 dout_21 clk vdd gnd
+ dff
Xdff_r0_c22
+ din_22 dout_22 clk vdd gnd
+ dff
Xdff_r0_c23
+ din_23 dout_23 clk vdd gnd
+ dff
Xdff_r0_c24
+ din_24 dout_24 clk vdd gnd
+ dff
Xdff_r0_c25
+ din_25 dout_25 clk vdd gnd
+ dff
Xdff_r0_c26
+ din_26 dout_26 clk vdd gnd
+ dff
Xdff_r0_c27
+ din_27 dout_27 clk vdd gnd
+ dff
Xdff_r0_c28
+ din_28 dout_28 clk vdd gnd
+ dff
Xdff_r0_c29
+ din_29 dout_29 clk vdd gnd
+ dff
Xdff_r0_c30
+ din_30 dout_30 clk vdd gnd
+ dff
Xdff_r0_c31
+ din_31 dout_31 clk vdd gnd
+ dff
Xdff_r0_c32
+ din_32 dout_32 clk vdd gnd
+ dff
Xdff_r0_c33
+ din_33 dout_33 clk vdd gnd
+ dff
Xdff_r0_c34
+ din_34 dout_34 clk vdd gnd
+ dff
Xdff_r0_c35
+ din_35 dout_35 clk vdd gnd
+ dff
Xdff_r0_c36
+ din_36 dout_36 clk vdd gnd
+ dff
Xdff_r0_c37
+ din_37 dout_37 clk vdd gnd
+ dff
Xdff_r0_c38
+ din_38 dout_38 clk vdd gnd
+ dff
Xdff_r0_c39
+ din_39 dout_39 clk vdd gnd
+ dff
Xdff_r0_c40
+ din_40 dout_40 clk vdd gnd
+ dff
Xdff_r0_c41
+ din_41 dout_41 clk vdd gnd
+ dff
Xdff_r0_c42
+ din_42 dout_42 clk vdd gnd
+ dff
Xdff_r0_c43
+ din_43 dout_43 clk vdd gnd
+ dff
Xdff_r0_c44
+ din_44 dout_44 clk vdd gnd
+ dff
Xdff_r0_c45
+ din_45 dout_45 clk vdd gnd
+ dff
Xdff_r0_c46
+ din_46 dout_46 clk vdd gnd
+ dff
Xdff_r0_c47
+ din_47 dout_47 clk vdd gnd
+ dff
Xdff_r0_c48
+ din_48 dout_48 clk vdd gnd
+ dff
Xdff_r0_c49
+ din_49 dout_49 clk vdd gnd
+ dff
Xdff_r0_c50
+ din_50 dout_50 clk vdd gnd
+ dff
Xdff_r0_c51
+ din_51 dout_51 clk vdd gnd
+ dff
Xdff_r0_c52
+ din_52 dout_52 clk vdd gnd
+ dff
Xdff_r0_c53
+ din_53 dout_53 clk vdd gnd
+ dff
Xdff_r0_c54
+ din_54 dout_54 clk vdd gnd
+ dff
Xdff_r0_c55
+ din_55 dout_55 clk vdd gnd
+ dff
Xdff_r0_c56
+ din_56 dout_56 clk vdd gnd
+ dff
Xdff_r0_c57
+ din_57 dout_57 clk vdd gnd
+ dff
Xdff_r0_c58
+ din_58 dout_58 clk vdd gnd
+ dff
Xdff_r0_c59
+ din_59 dout_59 clk vdd gnd
+ dff
Xdff_r0_c60
+ din_60 dout_60 clk vdd gnd
+ dff
Xdff_r0_c61
+ din_61 dout_61 clk vdd gnd
+ dff
Xdff_r0_c62
+ din_62 dout_62 clk vdd gnd
+ dff
Xdff_r0_c63
+ din_63 dout_63 clk vdd gnd
+ dff
Xdff_r0_c64
+ din_64 dout_64 clk vdd gnd
+ dff
Xdff_r0_c65
+ din_65 dout_65 clk vdd gnd
+ dff
Xdff_r0_c66
+ din_66 dout_66 clk vdd gnd
+ dff
Xdff_r0_c67
+ din_67 dout_67 clk vdd gnd
+ dff
Xdff_r0_c68
+ din_68 dout_68 clk vdd gnd
+ dff
Xdff_r0_c69
+ din_69 dout_69 clk vdd gnd
+ dff
Xdff_r0_c70
+ din_70 dout_70 clk vdd gnd
+ dff
Xdff_r0_c71
+ din_71 dout_71 clk vdd gnd
+ dff
Xdff_r0_c72
+ din_72 dout_72 clk vdd gnd
+ dff
Xdff_r0_c73
+ din_73 dout_73 clk vdd gnd
+ dff
Xdff_r0_c74
+ din_74 dout_74 clk vdd gnd
+ dff
Xdff_r0_c75
+ din_75 dout_75 clk vdd gnd
+ dff
Xdff_r0_c76
+ din_76 dout_76 clk vdd gnd
+ dff
Xdff_r0_c77
+ din_77 dout_77 clk vdd gnd
+ dff
Xdff_r0_c78
+ din_78 dout_78 clk vdd gnd
+ dff
Xdff_r0_c79
+ din_79 dout_79 clk vdd gnd
+ dff
Xdff_r0_c80
+ din_80 dout_80 clk vdd gnd
+ dff
Xdff_r0_c81
+ din_81 dout_81 clk vdd gnd
+ dff
Xdff_r0_c82
+ din_82 dout_82 clk vdd gnd
+ dff
Xdff_r0_c83
+ din_83 dout_83 clk vdd gnd
+ dff
Xdff_r0_c84
+ din_84 dout_84 clk vdd gnd
+ dff
Xdff_r0_c85
+ din_85 dout_85 clk vdd gnd
+ dff
Xdff_r0_c86
+ din_86 dout_86 clk vdd gnd
+ dff
Xdff_r0_c87
+ din_87 dout_87 clk vdd gnd
+ dff
Xdff_r0_c88
+ din_88 dout_88 clk vdd gnd
+ dff
Xdff_r0_c89
+ din_89 dout_89 clk vdd gnd
+ dff
Xdff_r0_c90
+ din_90 dout_90 clk vdd gnd
+ dff
Xdff_r0_c91
+ din_91 dout_91 clk vdd gnd
+ dff
Xdff_r0_c92
+ din_92 dout_92 clk vdd gnd
+ dff
Xdff_r0_c93
+ din_93 dout_93 clk vdd gnd
+ dff
Xdff_r0_c94
+ din_94 dout_94 clk vdd gnd
+ dff
Xdff_r0_c95
+ din_95 dout_95 clk vdd gnd
+ dff
Xdff_r0_c96
+ din_96 dout_96 clk vdd gnd
+ dff
Xdff_r0_c97
+ din_97 dout_97 clk vdd gnd
+ dff
Xdff_r0_c98
+ din_98 dout_98 clk vdd gnd
+ dff
Xdff_r0_c99
+ din_99 dout_99 clk vdd gnd
+ dff
Xdff_r0_c100
+ din_100 dout_100 clk vdd gnd
+ dff
Xdff_r0_c101
+ din_101 dout_101 clk vdd gnd
+ dff
Xdff_r0_c102
+ din_102 dout_102 clk vdd gnd
+ dff
Xdff_r0_c103
+ din_103 dout_103 clk vdd gnd
+ dff
Xdff_r0_c104
+ din_104 dout_104 clk vdd gnd
+ dff
Xdff_r0_c105
+ din_105 dout_105 clk vdd gnd
+ dff
Xdff_r0_c106
+ din_106 dout_106 clk vdd gnd
+ dff
Xdff_r0_c107
+ din_107 dout_107 clk vdd gnd
+ dff
Xdff_r0_c108
+ din_108 dout_108 clk vdd gnd
+ dff
Xdff_r0_c109
+ din_109 dout_109 clk vdd gnd
+ dff
Xdff_r0_c110
+ din_110 dout_110 clk vdd gnd
+ dff
Xdff_r0_c111
+ din_111 dout_111 clk vdd gnd
+ dff
Xdff_r0_c112
+ din_112 dout_112 clk vdd gnd
+ dff
Xdff_r0_c113
+ din_113 dout_113 clk vdd gnd
+ dff
Xdff_r0_c114
+ din_114 dout_114 clk vdd gnd
+ dff
Xdff_r0_c115
+ din_115 dout_115 clk vdd gnd
+ dff
Xdff_r0_c116
+ din_116 dout_116 clk vdd gnd
+ dff
Xdff_r0_c117
+ din_117 dout_117 clk vdd gnd
+ dff
Xdff_r0_c118
+ din_118 dout_118 clk vdd gnd
+ dff
Xdff_r0_c119
+ din_119 dout_119 clk vdd gnd
+ dff
Xdff_r0_c120
+ din_120 dout_120 clk vdd gnd
+ dff
Xdff_r0_c121
+ din_121 dout_121 clk vdd gnd
+ dff
Xdff_r0_c122
+ din_122 dout_122 clk vdd gnd
+ dff
Xdff_r0_c123
+ din_123 dout_123 clk vdd gnd
+ dff
Xdff_r0_c124
+ din_124 dout_124 clk vdd gnd
+ dff
Xdff_r0_c125
+ din_125 dout_125 clk vdd gnd
+ dff
Xdff_r0_c126
+ din_126 dout_126 clk vdd gnd
+ dff
Xdff_r0_c127
+ din_127 dout_127 clk vdd gnd
+ dff
Xdff_r0_c128
+ din_128 dout_128 clk vdd gnd
+ dff
Xdff_r0_c129
+ din_129 dout_129 clk vdd gnd
+ dff
Xdff_r0_c130
+ din_130 dout_130 clk vdd gnd
+ dff
Xdff_r0_c131
+ din_131 dout_131 clk vdd gnd
+ dff
Xdff_r0_c132
+ din_132 dout_132 clk vdd gnd
+ dff
Xdff_r0_c133
+ din_133 dout_133 clk vdd gnd
+ dff
Xdff_r0_c134
+ din_134 dout_134 clk vdd gnd
+ dff
Xdff_r0_c135
+ din_135 dout_135 clk vdd gnd
+ dff
Xdff_r0_c136
+ din_136 dout_136 clk vdd gnd
+ dff
Xdff_r0_c137
+ din_137 dout_137 clk vdd gnd
+ dff
Xdff_r0_c138
+ din_138 dout_138 clk vdd gnd
+ dff
Xdff_r0_c139
+ din_139 dout_139 clk vdd gnd
+ dff
Xdff_r0_c140
+ din_140 dout_140 clk vdd gnd
+ dff
Xdff_r0_c141
+ din_141 dout_141 clk vdd gnd
+ dff
Xdff_r0_c142
+ din_142 dout_142 clk vdd gnd
+ dff
Xdff_r0_c143
+ din_143 dout_143 clk vdd gnd
+ dff
Xdff_r0_c144
+ din_144 dout_144 clk vdd gnd
+ dff
Xdff_r0_c145
+ din_145 dout_145 clk vdd gnd
+ dff
Xdff_r0_c146
+ din_146 dout_146 clk vdd gnd
+ dff
Xdff_r0_c147
+ din_147 dout_147 clk vdd gnd
+ dff
Xdff_r0_c148
+ din_148 dout_148 clk vdd gnd
+ dff
Xdff_r0_c149
+ din_149 dout_149 clk vdd gnd
+ dff
Xdff_r0_c150
+ din_150 dout_150 clk vdd gnd
+ dff
Xdff_r0_c151
+ din_151 dout_151 clk vdd gnd
+ dff
Xdff_r0_c152
+ din_152 dout_152 clk vdd gnd
+ dff
Xdff_r0_c153
+ din_153 dout_153 clk vdd gnd
+ dff
Xdff_r0_c154
+ din_154 dout_154 clk vdd gnd
+ dff
Xdff_r0_c155
+ din_155 dout_155 clk vdd gnd
+ dff
Xdff_r0_c156
+ din_156 dout_156 clk vdd gnd
+ dff
Xdff_r0_c157
+ din_157 dout_157 clk vdd gnd
+ dff
Xdff_r0_c158
+ din_158 dout_158 clk vdd gnd
+ dff
Xdff_r0_c159
+ din_159 dout_159 clk vdd gnd
+ dff
Xdff_r0_c160
+ din_160 dout_160 clk vdd gnd
+ dff
Xdff_r0_c161
+ din_161 dout_161 clk vdd gnd
+ dff
Xdff_r0_c162
+ din_162 dout_162 clk vdd gnd
+ dff
Xdff_r0_c163
+ din_163 dout_163 clk vdd gnd
+ dff
Xdff_r0_c164
+ din_164 dout_164 clk vdd gnd
+ dff
Xdff_r0_c165
+ din_165 dout_165 clk vdd gnd
+ dff
Xdff_r0_c166
+ din_166 dout_166 clk vdd gnd
+ dff
Xdff_r0_c167
+ din_167 dout_167 clk vdd gnd
+ dff
Xdff_r0_c168
+ din_168 dout_168 clk vdd gnd
+ dff
Xdff_r0_c169
+ din_169 dout_169 clk vdd gnd
+ dff
Xdff_r0_c170
+ din_170 dout_170 clk vdd gnd
+ dff
Xdff_r0_c171
+ din_171 dout_171 clk vdd gnd
+ dff
Xdff_r0_c172
+ din_172 dout_172 clk vdd gnd
+ dff
Xdff_r0_c173
+ din_173 dout_173 clk vdd gnd
+ dff
Xdff_r0_c174
+ din_174 dout_174 clk vdd gnd
+ dff
Xdff_r0_c175
+ din_175 dout_175 clk vdd gnd
+ dff
Xdff_r0_c176
+ din_176 dout_176 clk vdd gnd
+ dff
Xdff_r0_c177
+ din_177 dout_177 clk vdd gnd
+ dff
Xdff_r0_c178
+ din_178 dout_178 clk vdd gnd
+ dff
Xdff_r0_c179
+ din_179 dout_179 clk vdd gnd
+ dff
Xdff_r0_c180
+ din_180 dout_180 clk vdd gnd
+ dff
Xdff_r0_c181
+ din_181 dout_181 clk vdd gnd
+ dff
Xdff_r0_c182
+ din_182 dout_182 clk vdd gnd
+ dff
Xdff_r0_c183
+ din_183 dout_183 clk vdd gnd
+ dff
Xdff_r0_c184
+ din_184 dout_184 clk vdd gnd
+ dff
Xdff_r0_c185
+ din_185 dout_185 clk vdd gnd
+ dff
Xdff_r0_c186
+ din_186 dout_186 clk vdd gnd
+ dff
Xdff_r0_c187
+ din_187 dout_187 clk vdd gnd
+ dff
Xdff_r0_c188
+ din_188 dout_188 clk vdd gnd
+ dff
Xdff_r0_c189
+ din_189 dout_189 clk vdd gnd
+ dff
Xdff_r0_c190
+ din_190 dout_190 clk vdd gnd
+ dff
Xdff_r0_c191
+ din_191 dout_191 clk vdd gnd
+ dff
Xdff_r0_c192
+ din_192 dout_192 clk vdd gnd
+ dff
Xdff_r0_c193
+ din_193 dout_193 clk vdd gnd
+ dff
Xdff_r0_c194
+ din_194 dout_194 clk vdd gnd
+ dff
Xdff_r0_c195
+ din_195 dout_195 clk vdd gnd
+ dff
Xdff_r0_c196
+ din_196 dout_196 clk vdd gnd
+ dff
Xdff_r0_c197
+ din_197 dout_197 clk vdd gnd
+ dff
Xdff_r0_c198
+ din_198 dout_198 clk vdd gnd
+ dff
Xdff_r0_c199
+ din_199 dout_199 clk vdd gnd
+ dff
Xdff_r0_c200
+ din_200 dout_200 clk vdd gnd
+ dff
Xdff_r0_c201
+ din_201 dout_201 clk vdd gnd
+ dff
Xdff_r0_c202
+ din_202 dout_202 clk vdd gnd
+ dff
Xdff_r0_c203
+ din_203 dout_203 clk vdd gnd
+ dff
Xdff_r0_c204
+ din_204 dout_204 clk vdd gnd
+ dff
Xdff_r0_c205
+ din_205 dout_205 clk vdd gnd
+ dff
Xdff_r0_c206
+ din_206 dout_206 clk vdd gnd
+ dff
Xdff_r0_c207
+ din_207 dout_207 clk vdd gnd
+ dff
Xdff_r0_c208
+ din_208 dout_208 clk vdd gnd
+ dff
Xdff_r0_c209
+ din_209 dout_209 clk vdd gnd
+ dff
Xdff_r0_c210
+ din_210 dout_210 clk vdd gnd
+ dff
Xdff_r0_c211
+ din_211 dout_211 clk vdd gnd
+ dff
Xdff_r0_c212
+ din_212 dout_212 clk vdd gnd
+ dff
Xdff_r0_c213
+ din_213 dout_213 clk vdd gnd
+ dff
Xdff_r0_c214
+ din_214 dout_214 clk vdd gnd
+ dff
Xdff_r0_c215
+ din_215 dout_215 clk vdd gnd
+ dff
Xdff_r0_c216
+ din_216 dout_216 clk vdd gnd
+ dff
Xdff_r0_c217
+ din_217 dout_217 clk vdd gnd
+ dff
Xdff_r0_c218
+ din_218 dout_218 clk vdd gnd
+ dff
Xdff_r0_c219
+ din_219 dout_219 clk vdd gnd
+ dff
Xdff_r0_c220
+ din_220 dout_220 clk vdd gnd
+ dff
Xdff_r0_c221
+ din_221 dout_221 clk vdd gnd
+ dff
Xdff_r0_c222
+ din_222 dout_222 clk vdd gnd
+ dff
Xdff_r0_c223
+ din_223 dout_223 clk vdd gnd
+ dff
Xdff_r0_c224
+ din_224 dout_224 clk vdd gnd
+ dff
Xdff_r0_c225
+ din_225 dout_225 clk vdd gnd
+ dff
Xdff_r0_c226
+ din_226 dout_226 clk vdd gnd
+ dff
Xdff_r0_c227
+ din_227 dout_227 clk vdd gnd
+ dff
Xdff_r0_c228
+ din_228 dout_228 clk vdd gnd
+ dff
Xdff_r0_c229
+ din_229 dout_229 clk vdd gnd
+ dff
Xdff_r0_c230
+ din_230 dout_230 clk vdd gnd
+ dff
Xdff_r0_c231
+ din_231 dout_231 clk vdd gnd
+ dff
Xdff_r0_c232
+ din_232 dout_232 clk vdd gnd
+ dff
Xdff_r0_c233
+ din_233 dout_233 clk vdd gnd
+ dff
Xdff_r0_c234
+ din_234 dout_234 clk vdd gnd
+ dff
Xdff_r0_c235
+ din_235 dout_235 clk vdd gnd
+ dff
Xdff_r0_c236
+ din_236 dout_236 clk vdd gnd
+ dff
Xdff_r0_c237
+ din_237 dout_237 clk vdd gnd
+ dff
Xdff_r0_c238
+ din_238 dout_238 clk vdd gnd
+ dff
Xdff_r0_c239
+ din_239 dout_239 clk vdd gnd
+ dff
Xdff_r0_c240
+ din_240 dout_240 clk vdd gnd
+ dff
Xdff_r0_c241
+ din_241 dout_241 clk vdd gnd
+ dff
Xdff_r0_c242
+ din_242 dout_242 clk vdd gnd
+ dff
Xdff_r0_c243
+ din_243 dout_243 clk vdd gnd
+ dff
Xdff_r0_c244
+ din_244 dout_244 clk vdd gnd
+ dff
Xdff_r0_c245
+ din_245 dout_245 clk vdd gnd
+ dff
Xdff_r0_c246
+ din_246 dout_246 clk vdd gnd
+ dff
Xdff_r0_c247
+ din_247 dout_247 clk vdd gnd
+ dff
Xdff_r0_c248
+ din_248 dout_248 clk vdd gnd
+ dff
Xdff_r0_c249
+ din_249 dout_249 clk vdd gnd
+ dff
Xdff_r0_c250
+ din_250 dout_250 clk vdd gnd
+ dff
Xdff_r0_c251
+ din_251 dout_251 clk vdd gnd
+ dff
Xdff_r0_c252
+ din_252 dout_252 clk vdd gnd
+ dff
Xdff_r0_c253
+ din_253 dout_253 clk vdd gnd
+ dff
Xdff_r0_c254
+ din_254 dout_254 clk vdd gnd
+ dff
Xdff_r0_c255
+ din_255 dout_255 clk vdd gnd
+ dff
Xdff_r0_c256
+ din_256 dout_256 clk vdd gnd
+ dff
Xdff_r0_c257
+ din_257 dout_257 clk vdd gnd
+ dff
Xdff_r0_c258
+ din_258 dout_258 clk vdd gnd
+ dff
Xdff_r0_c259
+ din_259 dout_259 clk vdd gnd
+ dff
Xdff_r0_c260
+ din_260 dout_260 clk vdd gnd
+ dff
Xdff_r0_c261
+ din_261 dout_261 clk vdd gnd
+ dff
Xdff_r0_c262
+ din_262 dout_262 clk vdd gnd
+ dff
Xdff_r0_c263
+ din_263 dout_263 clk vdd gnd
+ dff
Xdff_r0_c264
+ din_264 dout_264 clk vdd gnd
+ dff
Xdff_r0_c265
+ din_265 dout_265 clk vdd gnd
+ dff
Xdff_r0_c266
+ din_266 dout_266 clk vdd gnd
+ dff
Xdff_r0_c267
+ din_267 dout_267 clk vdd gnd
+ dff
Xdff_r0_c268
+ din_268 dout_268 clk vdd gnd
+ dff
Xdff_r0_c269
+ din_269 dout_269 clk vdd gnd
+ dff
Xdff_r0_c270
+ din_270 dout_270 clk vdd gnd
+ dff
Xdff_r0_c271
+ din_271 dout_271 clk vdd gnd
+ dff
Xdff_r0_c272
+ din_272 dout_272 clk vdd gnd
+ dff
Xdff_r0_c273
+ din_273 dout_273 clk vdd gnd
+ dff
Xdff_r0_c274
+ din_274 dout_274 clk vdd gnd
+ dff
Xdff_r0_c275
+ din_275 dout_275 clk vdd gnd
+ dff
Xdff_r0_c276
+ din_276 dout_276 clk vdd gnd
+ dff
Xdff_r0_c277
+ din_277 dout_277 clk vdd gnd
+ dff
Xdff_r0_c278
+ din_278 dout_278 clk vdd gnd
+ dff
Xdff_r0_c279
+ din_279 dout_279 clk vdd gnd
+ dff
Xdff_r0_c280
+ din_280 dout_280 clk vdd gnd
+ dff
Xdff_r0_c281
+ din_281 dout_281 clk vdd gnd
+ dff
Xdff_r0_c282
+ din_282 dout_282 clk vdd gnd
+ dff
Xdff_r0_c283
+ din_283 dout_283 clk vdd gnd
+ dff
Xdff_r0_c284
+ din_284 dout_284 clk vdd gnd
+ dff
Xdff_r0_c285
+ din_285 dout_285 clk vdd gnd
+ dff
Xdff_r0_c286
+ din_286 dout_286 clk vdd gnd
+ dff
Xdff_r0_c287
+ din_287 dout_287 clk vdd gnd
+ dff
Xdff_r0_c288
+ din_288 dout_288 clk vdd gnd
+ dff
Xdff_r0_c289
+ din_289 dout_289 clk vdd gnd
+ dff
Xdff_r0_c290
+ din_290 dout_290 clk vdd gnd
+ dff
Xdff_r0_c291
+ din_291 dout_291 clk vdd gnd
+ dff
Xdff_r0_c292
+ din_292 dout_292 clk vdd gnd
+ dff
Xdff_r0_c293
+ din_293 dout_293 clk vdd gnd
+ dff
Xdff_r0_c294
+ din_294 dout_294 clk vdd gnd
+ dff
Xdff_r0_c295
+ din_295 dout_295 clk vdd gnd
+ dff
Xdff_r0_c296
+ din_296 dout_296 clk vdd gnd
+ dff
Xdff_r0_c297
+ din_297 dout_297 clk vdd gnd
+ dff
Xdff_r0_c298
+ din_298 dout_298 clk vdd gnd
+ dff
Xdff_r0_c299
+ din_299 dout_299 clk vdd gnd
+ dff
Xdff_r0_c300
+ din_300 dout_300 clk vdd gnd
+ dff
Xdff_r0_c301
+ din_301 dout_301 clk vdd gnd
+ dff
Xdff_r0_c302
+ din_302 dout_302 clk vdd gnd
+ dff
Xdff_r0_c303
+ din_303 dout_303 clk vdd gnd
+ dff
Xdff_r0_c304
+ din_304 dout_304 clk vdd gnd
+ dff
Xdff_r0_c305
+ din_305 dout_305 clk vdd gnd
+ dff
Xdff_r0_c306
+ din_306 dout_306 clk vdd gnd
+ dff
Xdff_r0_c307
+ din_307 dout_307 clk vdd gnd
+ dff
Xdff_r0_c308
+ din_308 dout_308 clk vdd gnd
+ dff
Xdff_r0_c309
+ din_309 dout_309 clk vdd gnd
+ dff
Xdff_r0_c310
+ din_310 dout_310 clk vdd gnd
+ dff
Xdff_r0_c311
+ din_311 dout_311 clk vdd gnd
+ dff
Xdff_r0_c312
+ din_312 dout_312 clk vdd gnd
+ dff
Xdff_r0_c313
+ din_313 dout_313 clk vdd gnd
+ dff
Xdff_r0_c314
+ din_314 dout_314 clk vdd gnd
+ dff
Xdff_r0_c315
+ din_315 dout_315 clk vdd gnd
+ dff
Xdff_r0_c316
+ din_316 dout_316 clk vdd gnd
+ dff
Xdff_r0_c317
+ din_317 dout_317 clk vdd gnd
+ dff
Xdff_r0_c318
+ din_318 dout_318 clk vdd gnd
+ dff
Xdff_r0_c319
+ din_319 dout_319 clk vdd gnd
+ dff
Xdff_r0_c320
+ din_320 dout_320 clk vdd gnd
+ dff
Xdff_r0_c321
+ din_321 dout_321 clk vdd gnd
+ dff
Xdff_r0_c322
+ din_322 dout_322 clk vdd gnd
+ dff
Xdff_r0_c323
+ din_323 dout_323 clk vdd gnd
+ dff
Xdff_r0_c324
+ din_324 dout_324 clk vdd gnd
+ dff
Xdff_r0_c325
+ din_325 dout_325 clk vdd gnd
+ dff
Xdff_r0_c326
+ din_326 dout_326 clk vdd gnd
+ dff
Xdff_r0_c327
+ din_327 dout_327 clk vdd gnd
+ dff
Xdff_r0_c328
+ din_328 dout_328 clk vdd gnd
+ dff
Xdff_r0_c329
+ din_329 dout_329 clk vdd gnd
+ dff
Xdff_r0_c330
+ din_330 dout_330 clk vdd gnd
+ dff
Xdff_r0_c331
+ din_331 dout_331 clk vdd gnd
+ dff
Xdff_r0_c332
+ din_332 dout_332 clk vdd gnd
+ dff
Xdff_r0_c333
+ din_333 dout_333 clk vdd gnd
+ dff
Xdff_r0_c334
+ din_334 dout_334 clk vdd gnd
+ dff
Xdff_r0_c335
+ din_335 dout_335 clk vdd gnd
+ dff
Xdff_r0_c336
+ din_336 dout_336 clk vdd gnd
+ dff
Xdff_r0_c337
+ din_337 dout_337 clk vdd gnd
+ dff
Xdff_r0_c338
+ din_338 dout_338 clk vdd gnd
+ dff
Xdff_r0_c339
+ din_339 dout_339 clk vdd gnd
+ dff
Xdff_r0_c340
+ din_340 dout_340 clk vdd gnd
+ dff
Xdff_r0_c341
+ din_341 dout_341 clk vdd gnd
+ dff
Xdff_r0_c342
+ din_342 dout_342 clk vdd gnd
+ dff
Xdff_r0_c343
+ din_343 dout_343 clk vdd gnd
+ dff
Xdff_r0_c344
+ din_344 dout_344 clk vdd gnd
+ dff
Xdff_r0_c345
+ din_345 dout_345 clk vdd gnd
+ dff
Xdff_r0_c346
+ din_346 dout_346 clk vdd gnd
+ dff
Xdff_r0_c347
+ din_347 dout_347 clk vdd gnd
+ dff
Xdff_r0_c348
+ din_348 dout_348 clk vdd gnd
+ dff
Xdff_r0_c349
+ din_349 dout_349 clk vdd gnd
+ dff
Xdff_r0_c350
+ din_350 dout_350 clk vdd gnd
+ dff
Xdff_r0_c351
+ din_351 dout_351 clk vdd gnd
+ dff
Xdff_r0_c352
+ din_352 dout_352 clk vdd gnd
+ dff
Xdff_r0_c353
+ din_353 dout_353 clk vdd gnd
+ dff
Xdff_r0_c354
+ din_354 dout_354 clk vdd gnd
+ dff
Xdff_r0_c355
+ din_355 dout_355 clk vdd gnd
+ dff
Xdff_r0_c356
+ din_356 dout_356 clk vdd gnd
+ dff
Xdff_r0_c357
+ din_357 dout_357 clk vdd gnd
+ dff
Xdff_r0_c358
+ din_358 dout_358 clk vdd gnd
+ dff
Xdff_r0_c359
+ din_359 dout_359 clk vdd gnd
+ dff
Xdff_r0_c360
+ din_360 dout_360 clk vdd gnd
+ dff
Xdff_r0_c361
+ din_361 dout_361 clk vdd gnd
+ dff
Xdff_r0_c362
+ din_362 dout_362 clk vdd gnd
+ dff
Xdff_r0_c363
+ din_363 dout_363 clk vdd gnd
+ dff
Xdff_r0_c364
+ din_364 dout_364 clk vdd gnd
+ dff
Xdff_r0_c365
+ din_365 dout_365 clk vdd gnd
+ dff
Xdff_r0_c366
+ din_366 dout_366 clk vdd gnd
+ dff
Xdff_r0_c367
+ din_367 dout_367 clk vdd gnd
+ dff
Xdff_r0_c368
+ din_368 dout_368 clk vdd gnd
+ dff
Xdff_r0_c369
+ din_369 dout_369 clk vdd gnd
+ dff
Xdff_r0_c370
+ din_370 dout_370 clk vdd gnd
+ dff
Xdff_r0_c371
+ din_371 dout_371 clk vdd gnd
+ dff
Xdff_r0_c372
+ din_372 dout_372 clk vdd gnd
+ dff
Xdff_r0_c373
+ din_373 dout_373 clk vdd gnd
+ dff
Xdff_r0_c374
+ din_374 dout_374 clk vdd gnd
+ dff
Xdff_r0_c375
+ din_375 dout_375 clk vdd gnd
+ dff
Xdff_r0_c376
+ din_376 dout_376 clk vdd gnd
+ dff
Xdff_r0_c377
+ din_377 dout_377 clk vdd gnd
+ dff
Xdff_r0_c378
+ din_378 dout_378 clk vdd gnd
+ dff
Xdff_r0_c379
+ din_379 dout_379 clk vdd gnd
+ dff
Xdff_r0_c380
+ din_380 dout_380 clk vdd gnd
+ dff
Xdff_r0_c381
+ din_381 dout_381 clk vdd gnd
+ dff
Xdff_r0_c382
+ din_382 dout_382 clk vdd gnd
+ dff
Xdff_r0_c383
+ din_383 dout_383 clk vdd gnd
+ dff
Xdff_r0_c384
+ din_384 dout_384 clk vdd gnd
+ dff
Xdff_r0_c385
+ din_385 dout_385 clk vdd gnd
+ dff
Xdff_r0_c386
+ din_386 dout_386 clk vdd gnd
+ dff
Xdff_r0_c387
+ din_387 dout_387 clk vdd gnd
+ dff
Xdff_r0_c388
+ din_388 dout_388 clk vdd gnd
+ dff
Xdff_r0_c389
+ din_389 dout_389 clk vdd gnd
+ dff
Xdff_r0_c390
+ din_390 dout_390 clk vdd gnd
+ dff
Xdff_r0_c391
+ din_391 dout_391 clk vdd gnd
+ dff
Xdff_r0_c392
+ din_392 dout_392 clk vdd gnd
+ dff
Xdff_r0_c393
+ din_393 dout_393 clk vdd gnd
+ dff
Xdff_r0_c394
+ din_394 dout_394 clk vdd gnd
+ dff
Xdff_r0_c395
+ din_395 dout_395 clk vdd gnd
+ dff
Xdff_r0_c396
+ din_396 dout_396 clk vdd gnd
+ dff
Xdff_r0_c397
+ din_397 dout_397 clk vdd gnd
+ dff
Xdff_r0_c398
+ din_398 dout_398 clk vdd gnd
+ dff
Xdff_r0_c399
+ din_399 dout_399 clk vdd gnd
+ dff
Xdff_r0_c400
+ din_400 dout_400 clk vdd gnd
+ dff
Xdff_r0_c401
+ din_401 dout_401 clk vdd gnd
+ dff
Xdff_r0_c402
+ din_402 dout_402 clk vdd gnd
+ dff
Xdff_r0_c403
+ din_403 dout_403 clk vdd gnd
+ dff
Xdff_r0_c404
+ din_404 dout_404 clk vdd gnd
+ dff
Xdff_r0_c405
+ din_405 dout_405 clk vdd gnd
+ dff
Xdff_r0_c406
+ din_406 dout_406 clk vdd gnd
+ dff
Xdff_r0_c407
+ din_407 dout_407 clk vdd gnd
+ dff
Xdff_r0_c408
+ din_408 dout_408 clk vdd gnd
+ dff
Xdff_r0_c409
+ din_409 dout_409 clk vdd gnd
+ dff
Xdff_r0_c410
+ din_410 dout_410 clk vdd gnd
+ dff
Xdff_r0_c411
+ din_411 dout_411 clk vdd gnd
+ dff
Xdff_r0_c412
+ din_412 dout_412 clk vdd gnd
+ dff
Xdff_r0_c413
+ din_413 dout_413 clk vdd gnd
+ dff
Xdff_r0_c414
+ din_414 dout_414 clk vdd gnd
+ dff
Xdff_r0_c415
+ din_415 dout_415 clk vdd gnd
+ dff
Xdff_r0_c416
+ din_416 dout_416 clk vdd gnd
+ dff
Xdff_r0_c417
+ din_417 dout_417 clk vdd gnd
+ dff
Xdff_r0_c418
+ din_418 dout_418 clk vdd gnd
+ dff
Xdff_r0_c419
+ din_419 dout_419 clk vdd gnd
+ dff
Xdff_r0_c420
+ din_420 dout_420 clk vdd gnd
+ dff
Xdff_r0_c421
+ din_421 dout_421 clk vdd gnd
+ dff
Xdff_r0_c422
+ din_422 dout_422 clk vdd gnd
+ dff
Xdff_r0_c423
+ din_423 dout_423 clk vdd gnd
+ dff
Xdff_r0_c424
+ din_424 dout_424 clk vdd gnd
+ dff
Xdff_r0_c425
+ din_425 dout_425 clk vdd gnd
+ dff
Xdff_r0_c426
+ din_426 dout_426 clk vdd gnd
+ dff
Xdff_r0_c427
+ din_427 dout_427 clk vdd gnd
+ dff
Xdff_r0_c428
+ din_428 dout_428 clk vdd gnd
+ dff
Xdff_r0_c429
+ din_429 dout_429 clk vdd gnd
+ dff
Xdff_r0_c430
+ din_430 dout_430 clk vdd gnd
+ dff
Xdff_r0_c431
+ din_431 dout_431 clk vdd gnd
+ dff
Xdff_r0_c432
+ din_432 dout_432 clk vdd gnd
+ dff
Xdff_r0_c433
+ din_433 dout_433 clk vdd gnd
+ dff
Xdff_r0_c434
+ din_434 dout_434 clk vdd gnd
+ dff
Xdff_r0_c435
+ din_435 dout_435 clk vdd gnd
+ dff
Xdff_r0_c436
+ din_436 dout_436 clk vdd gnd
+ dff
Xdff_r0_c437
+ din_437 dout_437 clk vdd gnd
+ dff
Xdff_r0_c438
+ din_438 dout_438 clk vdd gnd
+ dff
Xdff_r0_c439
+ din_439 dout_439 clk vdd gnd
+ dff
Xdff_r0_c440
+ din_440 dout_440 clk vdd gnd
+ dff
Xdff_r0_c441
+ din_441 dout_441 clk vdd gnd
+ dff
Xdff_r0_c442
+ din_442 dout_442 clk vdd gnd
+ dff
Xdff_r0_c443
+ din_443 dout_443 clk vdd gnd
+ dff
Xdff_r0_c444
+ din_444 dout_444 clk vdd gnd
+ dff
Xdff_r0_c445
+ din_445 dout_445 clk vdd gnd
+ dff
Xdff_r0_c446
+ din_446 dout_446 clk vdd gnd
+ dff
Xdff_r0_c447
+ din_447 dout_447 clk vdd gnd
+ dff
Xdff_r0_c448
+ din_448 dout_448 clk vdd gnd
+ dff
Xdff_r0_c449
+ din_449 dout_449 clk vdd gnd
+ dff
Xdff_r0_c450
+ din_450 dout_450 clk vdd gnd
+ dff
Xdff_r0_c451
+ din_451 dout_451 clk vdd gnd
+ dff
Xdff_r0_c452
+ din_452 dout_452 clk vdd gnd
+ dff
Xdff_r0_c453
+ din_453 dout_453 clk vdd gnd
+ dff
Xdff_r0_c454
+ din_454 dout_454 clk vdd gnd
+ dff
Xdff_r0_c455
+ din_455 dout_455 clk vdd gnd
+ dff
Xdff_r0_c456
+ din_456 dout_456 clk vdd gnd
+ dff
Xdff_r0_c457
+ din_457 dout_457 clk vdd gnd
+ dff
Xdff_r0_c458
+ din_458 dout_458 clk vdd gnd
+ dff
Xdff_r0_c459
+ din_459 dout_459 clk vdd gnd
+ dff
Xdff_r0_c460
+ din_460 dout_460 clk vdd gnd
+ dff
Xdff_r0_c461
+ din_461 dout_461 clk vdd gnd
+ dff
Xdff_r0_c462
+ din_462 dout_462 clk vdd gnd
+ dff
Xdff_r0_c463
+ din_463 dout_463 clk vdd gnd
+ dff
Xdff_r0_c464
+ din_464 dout_464 clk vdd gnd
+ dff
Xdff_r0_c465
+ din_465 dout_465 clk vdd gnd
+ dff
Xdff_r0_c466
+ din_466 dout_466 clk vdd gnd
+ dff
Xdff_r0_c467
+ din_467 dout_467 clk vdd gnd
+ dff
Xdff_r0_c468
+ din_468 dout_468 clk vdd gnd
+ dff
Xdff_r0_c469
+ din_469 dout_469 clk vdd gnd
+ dff
Xdff_r0_c470
+ din_470 dout_470 clk vdd gnd
+ dff
Xdff_r0_c471
+ din_471 dout_471 clk vdd gnd
+ dff
Xdff_r0_c472
+ din_472 dout_472 clk vdd gnd
+ dff
Xdff_r0_c473
+ din_473 dout_473 clk vdd gnd
+ dff
Xdff_r0_c474
+ din_474 dout_474 clk vdd gnd
+ dff
Xdff_r0_c475
+ din_475 dout_475 clk vdd gnd
+ dff
Xdff_r0_c476
+ din_476 dout_476 clk vdd gnd
+ dff
Xdff_r0_c477
+ din_477 dout_477 clk vdd gnd
+ dff
Xdff_r0_c478
+ din_478 dout_478 clk vdd gnd
+ dff
Xdff_r0_c479
+ din_479 dout_479 clk vdd gnd
+ dff
Xdff_r0_c480
+ din_480 dout_480 clk vdd gnd
+ dff
Xdff_r0_c481
+ din_481 dout_481 clk vdd gnd
+ dff
Xdff_r0_c482
+ din_482 dout_482 clk vdd gnd
+ dff
Xdff_r0_c483
+ din_483 dout_483 clk vdd gnd
+ dff
Xdff_r0_c484
+ din_484 dout_484 clk vdd gnd
+ dff
Xdff_r0_c485
+ din_485 dout_485 clk vdd gnd
+ dff
Xdff_r0_c486
+ din_486 dout_486 clk vdd gnd
+ dff
Xdff_r0_c487
+ din_487 dout_487 clk vdd gnd
+ dff
Xdff_r0_c488
+ din_488 dout_488 clk vdd gnd
+ dff
Xdff_r0_c489
+ din_489 dout_489 clk vdd gnd
+ dff
Xdff_r0_c490
+ din_490 dout_490 clk vdd gnd
+ dff
Xdff_r0_c491
+ din_491 dout_491 clk vdd gnd
+ dff
Xdff_r0_c492
+ din_492 dout_492 clk vdd gnd
+ dff
Xdff_r0_c493
+ din_493 dout_493 clk vdd gnd
+ dff
Xdff_r0_c494
+ din_494 dout_494 clk vdd gnd
+ dff
Xdff_r0_c495
+ din_495 dout_495 clk vdd gnd
+ dff
Xdff_r0_c496
+ din_496 dout_496 clk vdd gnd
+ dff
Xdff_r0_c497
+ din_497 dout_497 clk vdd gnd
+ dff
Xdff_r0_c498
+ din_498 dout_498 clk vdd gnd
+ dff
Xdff_r0_c499
+ din_499 dout_499 clk vdd gnd
+ dff
Xdff_r0_c500
+ din_500 dout_500 clk vdd gnd
+ dff
Xdff_r0_c501
+ din_501 dout_501 clk vdd gnd
+ dff
Xdff_r0_c502
+ din_502 dout_502 clk vdd gnd
+ dff
Xdff_r0_c503
+ din_503 dout_503 clk vdd gnd
+ dff
Xdff_r0_c504
+ din_504 dout_504 clk vdd gnd
+ dff
Xdff_r0_c505
+ din_505 dout_505 clk vdd gnd
+ dff
Xdff_r0_c506
+ din_506 dout_506 clk vdd gnd
+ dff
Xdff_r0_c507
+ din_507 dout_507 clk vdd gnd
+ dff
Xdff_r0_c508
+ din_508 dout_508 clk vdd gnd
+ dff
Xdff_r0_c509
+ din_509 dout_509 clk vdd gnd
+ dff
Xdff_r0_c510
+ din_510 dout_510 clk vdd gnd
+ dff
Xdff_r0_c511
+ din_511 dout_511 clk vdd gnd
+ dff
.ENDS freepdk45_sram_1rw0r_45x512_data_dff

* spice ptx M{0} {1} pmos_vtg m=153 w=0.9175u l=0.05u pd=1.94u ps=1.94u as=0.11p ad=0.11p

* spice ptx M{0} {1} nmos_vtg m=153 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_15
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=153 w=0.9175u l=0.05u pd=1.94u ps=1.94u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=153 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_15

.SUBCKT freepdk45_sram_1rw0r_45x512_pdriver_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [520]
Xbuf_inv1
+ A Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_15
.ENDS freepdk45_sram_1rw0r_45x512_pdriver_2

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* spice ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT freepdk45_sram_1rw0r_45x512_pnand3_0
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pnand3_0

.SUBCKT freepdk45_sram_1rw0r_45x512_pand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand
+ A B C zb_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pdriver_2
.ENDS freepdk45_sram_1rw0r_45x512_pand3

* spice ptx M{0} {1} nmos_vtg m=17 w=0.3025u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=17 w=0.905u l=0.05u pd=1.91u ps=1.91u as=0.11p ad=0.11p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_21
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=17 w=0.905u l=0.05u pd=1.91u ps=1.91u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=17 w=0.3025u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_21

* spice ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* spice ptx M{0} {1} nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_6
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_6

* spice ptx M{0} {1} nmos_vtg m=6 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=6 w=0.855u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_20
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=6 w=0.855u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=6 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_20

* spice ptx M{0} {1} pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_18
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_18

* spice ptx M{0} {1} pmos_vtg m=51 w=0.905u l=0.05u pd=1.91u ps=1.91u as=0.11p ad=0.11p

* spice ptx M{0} {1} nmos_vtg m=51 w=0.3025u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_22
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=51 w=0.905u l=0.05u pd=1.91u ps=1.91u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=51 w=0.3025u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_22

* spice ptx M{0} {1} nmos_vtg m=2 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* spice ptx M{0} {1} pmos_vtg m=2 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_19
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_19

.SUBCKT freepdk45_sram_1rw0r_45x512_pdriver_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 2, 6, 19, 57, 171]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_18
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_19
Xbuf_inv6
+ Zb5_int Zb6_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_20
Xbuf_inv7
+ Zb6_int Zb7_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_21
Xbuf_inv8
+ Zb7_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_22
.ENDS freepdk45_sram_1rw0r_45x512_pdriver_4

* spice ptx M{0} {1} nmos_vtg m=150 w=0.3075u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=150 w=0.9225u l=0.05u pd=1.95u ps=1.95u as=0.12p ad=0.12p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_16
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=150 w=0.9225u l=0.05u pd=1.95u ps=1.95u as=0.12p ad=0.12p
Mpinv_nmos Z A gnd gnd nmos_vtg m=150 w=0.3075u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_16

.SUBCKT freepdk45_sram_1rw0r_45x512_pdriver_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [512]
Xbuf_inv1
+ A Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_16
.ENDS freepdk45_sram_1rw0r_45x512_pdriver_3

.SUBCKT freepdk45_sram_1rw0r_45x512_pand3_0
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand
+ A B C zb_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pdriver_3
.ENDS freepdk45_sram_1rw0r_45x512_pand3_0

* spice ptx M{0} {1} pmos_vtg m=4 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

* spice ptx M{0} {1} nmos_vtg m=4 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=4 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=4 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_3

.SUBCKT freepdk45_sram_1rw0r_45x512_pdriver
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [12]
Xbuf_inv1
+ A Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_3
.ENDS freepdk45_sram_1rw0r_45x512_pdriver

.SUBCKT freepdk45_sram_1rw0r_45x512_pnand2_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pnand2_0

.SUBCKT freepdk45_sram_1rw0r_45x512_pand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand
+ A B zb_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand2_0
Xpand2_inv
+ zb_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pdriver
.ENDS freepdk45_sram_1rw0r_45x512_pand2

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_23
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_23

.SUBCKT freepdk45_sram_1rw0r_45x512_delay_chain
+ in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0
+ in dout_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_0_0
+ dout_1 n_0_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_0_1
+ dout_1 n_0_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_0_2
+ dout_1 n_0_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_0_3
+ dout_1 n_0_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv1
+ dout_1 dout_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_1_0
+ dout_2 n_1_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_1_1
+ dout_2 n_1_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_1_2
+ dout_2 n_1_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_1_3
+ dout_2 n_1_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv2
+ dout_2 dout_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_2_0
+ dout_3 n_2_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_2_1
+ dout_3 n_2_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_2_2
+ dout_3 n_2_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_2_3
+ dout_3 n_2_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv3
+ dout_3 dout_4 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_3_0
+ dout_4 n_3_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_3_1
+ dout_4 n_3_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_3_2
+ dout_4 n_3_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_3_3
+ dout_4 n_3_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv4
+ dout_4 dout_5 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_4_0
+ dout_5 n_4_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_4_1
+ dout_5 n_4_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_4_2
+ dout_5 n_4_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_4_3
+ dout_5 n_4_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv5
+ dout_5 dout_6 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_5_0
+ dout_6 n_5_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_5_1
+ dout_6 n_5_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_5_2
+ dout_6 n_5_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_5_3
+ dout_6 n_5_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv6
+ dout_6 dout_7 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_6_0
+ dout_7 n_6_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_6_1
+ dout_7 n_6_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_6_2
+ dout_7 n_6_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_6_3
+ dout_7 n_6_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv7
+ dout_7 dout_8 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_7_0
+ dout_8 n_7_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_7_1
+ dout_8 n_7_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_7_2
+ dout_8 n_7_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_7_3
+ dout_8 n_7_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdinv8
+ dout_8 out vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_8_0
+ out n_8_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_8_1
+ out n_8_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_8_2
+ out n_8_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
Xdload_8_3
+ out n_8_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_23
.ENDS freepdk45_sram_1rw0r_45x512_delay_chain

.SUBCKT freepdk45_sram_1rw0r_45x512_pnand2_1
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pnand2_1

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_1

* spice ptx M{0} {1} nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* spice ptx M{0} {1} pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_2

.SUBCKT freepdk45_sram_1rw0r_45x512_dff_buf_0
+ D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff
+ D qint clk vdd gnd
+ dff
Xdff_buf_inv1
+ qint Qb vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_1
Xdff_buf_inv2
+ Qb Q vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_2
.ENDS freepdk45_sram_1rw0r_45x512_dff_buf_0

.SUBCKT freepdk45_sram_1rw0r_45x512_dff_buf_array
+ din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_r0_c0
+ din_0 dout_0 dout_bar_0 clk vdd gnd
+ freepdk45_sram_1rw0r_45x512_dff_buf_0
Xdff_r1_c0
+ din_1 dout_1 dout_bar_1 clk vdd gnd
+ freepdk45_sram_1rw0r_45x512_dff_buf_0
.ENDS freepdk45_sram_1rw0r_45x512_dff_buf_array

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_17
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_17

* spice ptx M{0} {1} nmos_vtg m=5 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* spice ptx M{0} {1} pmos_vtg m=5 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_14
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=5 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=5 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_14

* spice ptx M{0} {1} pmos_vtg m=2 w=0.675u l=0.05u pd=1.45u ps=1.45u as=0.08p ad=0.08p

* spice ptx M{0} {1} nmos_vtg m=2 w=0.225u l=0.05u pd=0.55u ps=0.55u as=0.03p ad=0.03p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_13
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.675u l=0.05u pd=1.45u ps=1.45u as=0.08p ad=0.08p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.225u l=0.05u pd=0.55u ps=0.55u as=0.03p ad=0.03p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_13

.SUBCKT freepdk45_sram_1rw0r_45x512_pdriver_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [5, 15]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_13
Xbuf_inv2
+ Zb1_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_14
.ENDS freepdk45_sram_1rw0r_45x512_pdriver_1

* spice ptx M{0} {1} pmos_vtg m=254 w=0.9225u l=0.05u pd=1.95u ps=1.95u as=0.12p ad=0.12p

* spice ptx M{0} {1} nmos_vtg m=254 w=0.3075u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_12
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=254 w=0.9225u l=0.05u pd=1.95u ps=1.95u as=0.12p ad=0.12p
Mpinv_nmos Z A gnd gnd nmos_vtg m=254 w=0.3075u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_12

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_7
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_7

* spice ptx M{0} {1} nmos_vtg m=29 w=0.2975u l=0.05u pd=0.69u ps=0.69u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=29 w=0.895u l=0.05u pd=1.89u ps=1.89u as=0.11p ad=0.11p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_10
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=29 w=0.895u l=0.05u pd=1.89u ps=1.89u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=29 w=0.2975u l=0.05u pd=0.69u ps=0.69u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_10

* spice ptx M{0} {1} nmos_vtg m=10 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=10 w=0.865u l=0.05u pd=1.83u ps=1.83u as=0.11p ad=0.11p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_9
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=10 w=0.865u l=0.05u pd=1.83u ps=1.83u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=10 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_9

* spice ptx M{0} {1} nmos_vtg m=4 w=0.2475u l=0.05u pd=0.59u ps=0.59u as=0.03p ad=0.03p

* spice ptx M{0} {1} pmos_vtg m=4 w=0.7425u l=0.05u pd=1.59u ps=1.59u as=0.09p ad=0.09p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_8
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=4 w=0.7425u l=0.05u pd=1.59u ps=1.59u as=0.09p ad=0.09p
Mpinv_nmos Z A gnd gnd nmos_vtg m=4 w=0.2475u l=0.05u pd=0.59u ps=0.59u as=0.03p ad=0.03p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_8

* spice ptx M{0} {1} pmos_vtg m=85 w=0.9175u l=0.05u pd=1.94u ps=1.94u as=0.11p ad=0.11p

* spice ptx M{0} {1} nmos_vtg m=85 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_11
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=85 w=0.9175u l=0.05u pd=1.94u ps=1.94u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=85 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_11

.SUBCKT freepdk45_sram_1rw0r_45x512_pdriver_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 1, 1, 1, 1, 1, 4, 11, 32, 96, 289, 867]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv6
+ Zb5_int Zb6_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv7
+ Zb6_int Zb7_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv8
+ Zb7_int Zb8_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_6
Xbuf_inv9
+ Zb8_int Zb9_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_7
Xbuf_inv10
+ Zb9_int Zb10_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_8
Xbuf_inv11
+ Zb10_int Zb11_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_9
Xbuf_inv12
+ Zb11_int Zb12_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_10
Xbuf_inv13
+ Zb12_int Zb13_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_11
Xbuf_inv14
+ Zb13_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_12
.ENDS freepdk45_sram_1rw0r_45x512_pdriver_0

.SUBCKT freepdk45_sram_1rw0r_45x512_control_logic_rw
+ csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* word_size 512
Xctrl_dffs
+ csb web cs_bar cs we_bar we clk_buf vdd gnd
+ freepdk45_sram_1rw0r_45x512_dff_buf_array
Xclkbuf
+ clk clk_buf vdd gnd
+ freepdk45_sram_1rw0r_45x512_pdriver_0
Xinv_clk_bar
+ clk_buf clk_bar vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_17
Xand2_gated_clk_bar
+ clk_bar cs gated_clk_bar vdd gnd
+ freepdk45_sram_1rw0r_45x512_pand2
Xand2_gated_clk_buf
+ clk_buf cs gated_clk_buf vdd gnd
+ freepdk45_sram_1rw0r_45x512_pand2
Xbuf_wl_en
+ gated_clk_bar wl_en vdd gnd
+ freepdk45_sram_1rw0r_45x512_pdriver_1
Xrbl_bl_delay_inv
+ rbl_bl_delay rbl_bl_delay_bar vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_17
Xw_en_and
+ we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd
+ freepdk45_sram_1rw0r_45x512_pand3
Xbuf_s_en_and
+ rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd
+ freepdk45_sram_1rw0r_45x512_pand3_0
Xdelay_chain
+ rbl_bl rbl_bl_delay vdd gnd
+ freepdk45_sram_1rw0r_45x512_delay_chain
Xnand_p_en_bar
+ gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand2_1
Xbuf_p_en_bar
+ p_en_bar_unbuf p_en_bar vdd gnd
+ freepdk45_sram_1rw0r_45x512_pdriver_4
.ENDS freepdk45_sram_1rw0r_45x512_control_logic_rw

* spice ptx M{0} {1} nmos_vtg m=94 w=0.1225u l=0.05u pd=0.34u ps=0.34u as=0.02p ad=0.02p

* spice ptx M{0} {1} pmos_vtg m=94 w=0.3675u l=0.05u pd=0.83u ps=0.83u as=0.05p ad=0.05p

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=94 w=0.3675u l=0.05u pd=0.83u ps=0.83u as=0.05p ad=0.05p
Mpinv_nmos Z A gnd gnd nmos_vtg m=94 w=0.1225u l=0.05u pd=0.34u ps=0.34u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pinv_0

.SUBCKT freepdk45_sram_1rw0r_45x512_pnand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pnand2

.SUBCKT freepdk45_sram_1rw0r_45x512_and2_dec_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 128
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand2
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_0
.ENDS freepdk45_sram_1rw0r_45x512_and2_dec_0

.SUBCKT freepdk45_sram_1rw0r_45x512_wordline_driver
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xwld_nand
+ A B zb_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand2
Xwl_driver
+ zb_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv_0
.ENDS freepdk45_sram_1rw0r_45x512_wordline_driver

.SUBCKT freepdk45_sram_1rw0r_45x512_wordline_driver_array
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12
+ in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23
+ in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34
+ in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 wl_0 wl_1
+ wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14
+ wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25
+ wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36
+ wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 45 cols: 512
Xwl_driver_and0
+ in_0 en wl_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and1
+ in_1 en wl_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and2
+ in_2 en wl_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and3
+ in_3 en wl_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and4
+ in_4 en wl_4 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and5
+ in_5 en wl_5 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and6
+ in_6 en wl_6 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and7
+ in_7 en wl_7 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and8
+ in_8 en wl_8 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and9
+ in_9 en wl_9 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and10
+ in_10 en wl_10 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and11
+ in_11 en wl_11 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and12
+ in_12 en wl_12 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and13
+ in_13 en wl_13 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and14
+ in_14 en wl_14 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and15
+ in_15 en wl_15 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and16
+ in_16 en wl_16 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and17
+ in_17 en wl_17 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and18
+ in_18 en wl_18 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and19
+ in_19 en wl_19 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and20
+ in_20 en wl_20 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and21
+ in_21 en wl_21 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and22
+ in_22 en wl_22 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and23
+ in_23 en wl_23 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and24
+ in_24 en wl_24 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and25
+ in_25 en wl_25 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and26
+ in_26 en wl_26 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and27
+ in_27 en wl_27 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and28
+ in_28 en wl_28 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and29
+ in_29 en wl_29 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and30
+ in_30 en wl_30 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and31
+ in_31 en wl_31 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and32
+ in_32 en wl_32 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and33
+ in_33 en wl_33 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and34
+ in_34 en wl_34 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and35
+ in_35 en wl_35 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and36
+ in_36 en wl_36 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and37
+ in_37 en wl_37 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and38
+ in_38 en wl_38 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and39
+ in_39 en wl_39 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and40
+ in_40 en wl_40 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and41
+ in_41 en wl_41 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and42
+ in_42 en wl_42 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and43
+ in_43 en wl_43 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
Xwl_driver_and44
+ in_44 en wl_44 vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver
.ENDS freepdk45_sram_1rw0r_45x512_wordline_driver_array

.SUBCKT freepdk45_sram_1rw0r_45x512_pinv
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS freepdk45_sram_1rw0r_45x512_pinv

.SUBCKT freepdk45_sram_1rw0r_45x512_and2_dec
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand2
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv
.ENDS freepdk45_sram_1rw0r_45x512_and2_dec

.SUBCKT freepdk45_sram_1rw0r_45x512_hierarchical_predecode2x4
+ in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv
XXpre2x4_and_0
+ inbar_0 inbar_1 out_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and2_dec
XXpre2x4_and_1
+ in_0 inbar_1 out_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and2_dec
XXpre2x4_and_2
+ inbar_0 in_1 out_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and2_dec
XXpre2x4_and_3
+ in_0 in_1 out_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and2_dec
.ENDS freepdk45_sram_1rw0r_45x512_hierarchical_predecode2x4

.SUBCKT freepdk45_sram_1rw0r_45x512_pnand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS freepdk45_sram_1rw0r_45x512_pnand3

.SUBCKT freepdk45_sram_1rw0r_45x512_and3_dec
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_dec_nand
+ A B C zb_int vdd gnd
+ freepdk45_sram_1rw0r_45x512_pnand3
Xpand3_dec_inv
+ zb_int Z vdd gnd
+ freepdk45_sram_1rw0r_45x512_pinv
.ENDS freepdk45_sram_1rw0r_45x512_and3_dec

.SUBCKT freepdk45_sram_1rw0r_45x512_hierarchical_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 decode_0 decode_1 decode_2
+ decode_3 decode_4 decode_5 decode_6 decode_7 decode_8 decode_9
+ decode_10 decode_11 decode_12 decode_13 decode_14 decode_15 decode_16
+ decode_17 decode_18 decode_19 decode_20 decode_21 decode_22 decode_23
+ decode_24 decode_25 decode_26 decode_27 decode_28 decode_29 decode_30
+ decode_31 decode_32 decode_33 decode_34 decode_35 decode_36 decode_37
+ decode_38 decode_39 decode_40 decode_41 decode_42 decode_43 decode_44
+ vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* POWER : vdd 
* GROUND: gnd 
Xpre_0
+ addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_hierarchical_predecode2x4
Xpre_1
+ addr_2 addr_3 out_4 out_5 out_6 out_7 vdd gnd
+ freepdk45_sram_1rw0r_45x512_hierarchical_predecode2x4
Xpre_2
+ addr_4 addr_5 out_8 out_9 out_10 out_11 vdd gnd
+ freepdk45_sram_1rw0r_45x512_hierarchical_predecode2x4
XDEC_AND_0
+ out_0 out_4 out_8 decode_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_16
+ out_0 out_4 out_9 decode_16 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_32
+ out_0 out_4 out_10 decode_32 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_4
+ out_0 out_5 out_8 decode_4 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_20
+ out_0 out_5 out_9 decode_20 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_36
+ out_0 out_5 out_10 decode_36 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_8
+ out_0 out_6 out_8 decode_8 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_24
+ out_0 out_6 out_9 decode_24 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_40
+ out_0 out_6 out_10 decode_40 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_12
+ out_0 out_7 out_8 decode_12 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_28
+ out_0 out_7 out_9 decode_28 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_44
+ out_0 out_7 out_10 decode_44 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_1
+ out_1 out_4 out_8 decode_1 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_17
+ out_1 out_4 out_9 decode_17 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_33
+ out_1 out_4 out_10 decode_33 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_5
+ out_1 out_5 out_8 decode_5 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_21
+ out_1 out_5 out_9 decode_21 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_37
+ out_1 out_5 out_10 decode_37 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_9
+ out_1 out_6 out_8 decode_9 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_25
+ out_1 out_6 out_9 decode_25 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_41
+ out_1 out_6 out_10 decode_41 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_13
+ out_1 out_7 out_8 decode_13 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_29
+ out_1 out_7 out_9 decode_29 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_2
+ out_2 out_4 out_8 decode_2 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_18
+ out_2 out_4 out_9 decode_18 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_34
+ out_2 out_4 out_10 decode_34 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_6
+ out_2 out_5 out_8 decode_6 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_22
+ out_2 out_5 out_9 decode_22 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_38
+ out_2 out_5 out_10 decode_38 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_10
+ out_2 out_6 out_8 decode_10 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_26
+ out_2 out_6 out_9 decode_26 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_42
+ out_2 out_6 out_10 decode_42 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_14
+ out_2 out_7 out_8 decode_14 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_30
+ out_2 out_7 out_9 decode_30 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_3
+ out_3 out_4 out_8 decode_3 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_19
+ out_3 out_4 out_9 decode_19 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_35
+ out_3 out_4 out_10 decode_35 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_7
+ out_3 out_5 out_8 decode_7 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_23
+ out_3 out_5 out_9 decode_23 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_39
+ out_3 out_5 out_10 decode_39 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_11
+ out_3 out_6 out_8 decode_11 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_27
+ out_3 out_6 out_9 decode_27 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_43
+ out_3 out_6 out_10 decode_43 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_15
+ out_3 out_7 out_8 decode_15 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
XDEC_AND_31
+ out_3 out_7 out_9 decode_31 vdd gnd
+ freepdk45_sram_1rw0r_45x512_and3_dec
.ENDS freepdk45_sram_1rw0r_45x512_hierarchical_decoder

.SUBCKT freepdk45_sram_1rw0r_45x512_port_address
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 wl_en wl_0 wl_1 wl_2 wl_3
+ wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26
+ wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37
+ wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 rbl_wl vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: rbl_wl 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 dec_out_0 dec_out_1
+ dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8
+ dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14
+ dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20
+ dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26
+ dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32
+ dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38
+ dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 vdd
+ gnd
+ freepdk45_sram_1rw0r_45x512_hierarchical_decoder
Xwordline_driver
+ dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6
+ dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12
+ dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18
+ dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24
+ dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30
+ dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36
+ dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42
+ dec_out_43 dec_out_44 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8
+ wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20
+ wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31
+ wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42
+ wl_43 wl_44 wl_en vdd gnd
+ freepdk45_sram_1rw0r_45x512_wordline_driver_array
Xrbl_driver
+ wl_en vdd rbl_wl vdd gnd
+ freepdk45_sram_1rw0r_45x512_and2_dec_0
.ENDS freepdk45_sram_1rw0r_45x512_port_address

.SUBCKT freepdk45_sram_1rw0r_45x512_precharge_0
+ bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Mlower_pmos bl en_bar br vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos1 bl en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos2 br en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS freepdk45_sram_1rw0r_45x512_precharge_0

.SUBCKT freepdk45_sram_1rw0r_45x512_precharge_array
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67
+ bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73
+ br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78
+ bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84
+ br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89
+ bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95
+ br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100
+ bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105
+ bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110
+ bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115
+ bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120
+ bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125
+ bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130
+ bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135
+ bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140
+ bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145
+ bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150
+ bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155
+ bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160
+ bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165
+ bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170
+ bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175
+ bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180
+ bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185
+ bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190
+ bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195
+ bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200
+ bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205
+ bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210
+ bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215
+ bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220
+ bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225
+ bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230
+ bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235
+ bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240
+ bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245
+ bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250
+ bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255
+ bl_256 br_256 bl_257 br_257 bl_258 br_258 bl_259 br_259 bl_260 br_260
+ bl_261 br_261 bl_262 br_262 bl_263 br_263 bl_264 br_264 bl_265 br_265
+ bl_266 br_266 bl_267 br_267 bl_268 br_268 bl_269 br_269 bl_270 br_270
+ bl_271 br_271 bl_272 br_272 bl_273 br_273 bl_274 br_274 bl_275 br_275
+ bl_276 br_276 bl_277 br_277 bl_278 br_278 bl_279 br_279 bl_280 br_280
+ bl_281 br_281 bl_282 br_282 bl_283 br_283 bl_284 br_284 bl_285 br_285
+ bl_286 br_286 bl_287 br_287 bl_288 br_288 bl_289 br_289 bl_290 br_290
+ bl_291 br_291 bl_292 br_292 bl_293 br_293 bl_294 br_294 bl_295 br_295
+ bl_296 br_296 bl_297 br_297 bl_298 br_298 bl_299 br_299 bl_300 br_300
+ bl_301 br_301 bl_302 br_302 bl_303 br_303 bl_304 br_304 bl_305 br_305
+ bl_306 br_306 bl_307 br_307 bl_308 br_308 bl_309 br_309 bl_310 br_310
+ bl_311 br_311 bl_312 br_312 bl_313 br_313 bl_314 br_314 bl_315 br_315
+ bl_316 br_316 bl_317 br_317 bl_318 br_318 bl_319 br_319 bl_320 br_320
+ bl_321 br_321 bl_322 br_322 bl_323 br_323 bl_324 br_324 bl_325 br_325
+ bl_326 br_326 bl_327 br_327 bl_328 br_328 bl_329 br_329 bl_330 br_330
+ bl_331 br_331 bl_332 br_332 bl_333 br_333 bl_334 br_334 bl_335 br_335
+ bl_336 br_336 bl_337 br_337 bl_338 br_338 bl_339 br_339 bl_340 br_340
+ bl_341 br_341 bl_342 br_342 bl_343 br_343 bl_344 br_344 bl_345 br_345
+ bl_346 br_346 bl_347 br_347 bl_348 br_348 bl_349 br_349 bl_350 br_350
+ bl_351 br_351 bl_352 br_352 bl_353 br_353 bl_354 br_354 bl_355 br_355
+ bl_356 br_356 bl_357 br_357 bl_358 br_358 bl_359 br_359 bl_360 br_360
+ bl_361 br_361 bl_362 br_362 bl_363 br_363 bl_364 br_364 bl_365 br_365
+ bl_366 br_366 bl_367 br_367 bl_368 br_368 bl_369 br_369 bl_370 br_370
+ bl_371 br_371 bl_372 br_372 bl_373 br_373 bl_374 br_374 bl_375 br_375
+ bl_376 br_376 bl_377 br_377 bl_378 br_378 bl_379 br_379 bl_380 br_380
+ bl_381 br_381 bl_382 br_382 bl_383 br_383 bl_384 br_384 bl_385 br_385
+ bl_386 br_386 bl_387 br_387 bl_388 br_388 bl_389 br_389 bl_390 br_390
+ bl_391 br_391 bl_392 br_392 bl_393 br_393 bl_394 br_394 bl_395 br_395
+ bl_396 br_396 bl_397 br_397 bl_398 br_398 bl_399 br_399 bl_400 br_400
+ bl_401 br_401 bl_402 br_402 bl_403 br_403 bl_404 br_404 bl_405 br_405
+ bl_406 br_406 bl_407 br_407 bl_408 br_408 bl_409 br_409 bl_410 br_410
+ bl_411 br_411 bl_412 br_412 bl_413 br_413 bl_414 br_414 bl_415 br_415
+ bl_416 br_416 bl_417 br_417 bl_418 br_418 bl_419 br_419 bl_420 br_420
+ bl_421 br_421 bl_422 br_422 bl_423 br_423 bl_424 br_424 bl_425 br_425
+ bl_426 br_426 bl_427 br_427 bl_428 br_428 bl_429 br_429 bl_430 br_430
+ bl_431 br_431 bl_432 br_432 bl_433 br_433 bl_434 br_434 bl_435 br_435
+ bl_436 br_436 bl_437 br_437 bl_438 br_438 bl_439 br_439 bl_440 br_440
+ bl_441 br_441 bl_442 br_442 bl_443 br_443 bl_444 br_444 bl_445 br_445
+ bl_446 br_446 bl_447 br_447 bl_448 br_448 bl_449 br_449 bl_450 br_450
+ bl_451 br_451 bl_452 br_452 bl_453 br_453 bl_454 br_454 bl_455 br_455
+ bl_456 br_456 bl_457 br_457 bl_458 br_458 bl_459 br_459 bl_460 br_460
+ bl_461 br_461 bl_462 br_462 bl_463 br_463 bl_464 br_464 bl_465 br_465
+ bl_466 br_466 bl_467 br_467 bl_468 br_468 bl_469 br_469 bl_470 br_470
+ bl_471 br_471 bl_472 br_472 bl_473 br_473 bl_474 br_474 bl_475 br_475
+ bl_476 br_476 bl_477 br_477 bl_478 br_478 bl_479 br_479 bl_480 br_480
+ bl_481 br_481 bl_482 br_482 bl_483 br_483 bl_484 br_484 bl_485 br_485
+ bl_486 br_486 bl_487 br_487 bl_488 br_488 bl_489 br_489 bl_490 br_490
+ bl_491 br_491 bl_492 br_492 bl_493 br_493 bl_494 br_494 bl_495 br_495
+ bl_496 br_496 bl_497 br_497 bl_498 br_498 bl_499 br_499 bl_500 br_500
+ bl_501 br_501 bl_502 br_502 bl_503 br_503 bl_504 br_504 bl_505 br_505
+ bl_506 br_506 bl_507 br_507 bl_508 br_508 bl_509 br_509 bl_510 br_510
+ bl_511 br_511 bl_512 br_512 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* OUTPUT: bl_130 
* OUTPUT: br_130 
* OUTPUT: bl_131 
* OUTPUT: br_131 
* OUTPUT: bl_132 
* OUTPUT: br_132 
* OUTPUT: bl_133 
* OUTPUT: br_133 
* OUTPUT: bl_134 
* OUTPUT: br_134 
* OUTPUT: bl_135 
* OUTPUT: br_135 
* OUTPUT: bl_136 
* OUTPUT: br_136 
* OUTPUT: bl_137 
* OUTPUT: br_137 
* OUTPUT: bl_138 
* OUTPUT: br_138 
* OUTPUT: bl_139 
* OUTPUT: br_139 
* OUTPUT: bl_140 
* OUTPUT: br_140 
* OUTPUT: bl_141 
* OUTPUT: br_141 
* OUTPUT: bl_142 
* OUTPUT: br_142 
* OUTPUT: bl_143 
* OUTPUT: br_143 
* OUTPUT: bl_144 
* OUTPUT: br_144 
* OUTPUT: bl_145 
* OUTPUT: br_145 
* OUTPUT: bl_146 
* OUTPUT: br_146 
* OUTPUT: bl_147 
* OUTPUT: br_147 
* OUTPUT: bl_148 
* OUTPUT: br_148 
* OUTPUT: bl_149 
* OUTPUT: br_149 
* OUTPUT: bl_150 
* OUTPUT: br_150 
* OUTPUT: bl_151 
* OUTPUT: br_151 
* OUTPUT: bl_152 
* OUTPUT: br_152 
* OUTPUT: bl_153 
* OUTPUT: br_153 
* OUTPUT: bl_154 
* OUTPUT: br_154 
* OUTPUT: bl_155 
* OUTPUT: br_155 
* OUTPUT: bl_156 
* OUTPUT: br_156 
* OUTPUT: bl_157 
* OUTPUT: br_157 
* OUTPUT: bl_158 
* OUTPUT: br_158 
* OUTPUT: bl_159 
* OUTPUT: br_159 
* OUTPUT: bl_160 
* OUTPUT: br_160 
* OUTPUT: bl_161 
* OUTPUT: br_161 
* OUTPUT: bl_162 
* OUTPUT: br_162 
* OUTPUT: bl_163 
* OUTPUT: br_163 
* OUTPUT: bl_164 
* OUTPUT: br_164 
* OUTPUT: bl_165 
* OUTPUT: br_165 
* OUTPUT: bl_166 
* OUTPUT: br_166 
* OUTPUT: bl_167 
* OUTPUT: br_167 
* OUTPUT: bl_168 
* OUTPUT: br_168 
* OUTPUT: bl_169 
* OUTPUT: br_169 
* OUTPUT: bl_170 
* OUTPUT: br_170 
* OUTPUT: bl_171 
* OUTPUT: br_171 
* OUTPUT: bl_172 
* OUTPUT: br_172 
* OUTPUT: bl_173 
* OUTPUT: br_173 
* OUTPUT: bl_174 
* OUTPUT: br_174 
* OUTPUT: bl_175 
* OUTPUT: br_175 
* OUTPUT: bl_176 
* OUTPUT: br_176 
* OUTPUT: bl_177 
* OUTPUT: br_177 
* OUTPUT: bl_178 
* OUTPUT: br_178 
* OUTPUT: bl_179 
* OUTPUT: br_179 
* OUTPUT: bl_180 
* OUTPUT: br_180 
* OUTPUT: bl_181 
* OUTPUT: br_181 
* OUTPUT: bl_182 
* OUTPUT: br_182 
* OUTPUT: bl_183 
* OUTPUT: br_183 
* OUTPUT: bl_184 
* OUTPUT: br_184 
* OUTPUT: bl_185 
* OUTPUT: br_185 
* OUTPUT: bl_186 
* OUTPUT: br_186 
* OUTPUT: bl_187 
* OUTPUT: br_187 
* OUTPUT: bl_188 
* OUTPUT: br_188 
* OUTPUT: bl_189 
* OUTPUT: br_189 
* OUTPUT: bl_190 
* OUTPUT: br_190 
* OUTPUT: bl_191 
* OUTPUT: br_191 
* OUTPUT: bl_192 
* OUTPUT: br_192 
* OUTPUT: bl_193 
* OUTPUT: br_193 
* OUTPUT: bl_194 
* OUTPUT: br_194 
* OUTPUT: bl_195 
* OUTPUT: br_195 
* OUTPUT: bl_196 
* OUTPUT: br_196 
* OUTPUT: bl_197 
* OUTPUT: br_197 
* OUTPUT: bl_198 
* OUTPUT: br_198 
* OUTPUT: bl_199 
* OUTPUT: br_199 
* OUTPUT: bl_200 
* OUTPUT: br_200 
* OUTPUT: bl_201 
* OUTPUT: br_201 
* OUTPUT: bl_202 
* OUTPUT: br_202 
* OUTPUT: bl_203 
* OUTPUT: br_203 
* OUTPUT: bl_204 
* OUTPUT: br_204 
* OUTPUT: bl_205 
* OUTPUT: br_205 
* OUTPUT: bl_206 
* OUTPUT: br_206 
* OUTPUT: bl_207 
* OUTPUT: br_207 
* OUTPUT: bl_208 
* OUTPUT: br_208 
* OUTPUT: bl_209 
* OUTPUT: br_209 
* OUTPUT: bl_210 
* OUTPUT: br_210 
* OUTPUT: bl_211 
* OUTPUT: br_211 
* OUTPUT: bl_212 
* OUTPUT: br_212 
* OUTPUT: bl_213 
* OUTPUT: br_213 
* OUTPUT: bl_214 
* OUTPUT: br_214 
* OUTPUT: bl_215 
* OUTPUT: br_215 
* OUTPUT: bl_216 
* OUTPUT: br_216 
* OUTPUT: bl_217 
* OUTPUT: br_217 
* OUTPUT: bl_218 
* OUTPUT: br_218 
* OUTPUT: bl_219 
* OUTPUT: br_219 
* OUTPUT: bl_220 
* OUTPUT: br_220 
* OUTPUT: bl_221 
* OUTPUT: br_221 
* OUTPUT: bl_222 
* OUTPUT: br_222 
* OUTPUT: bl_223 
* OUTPUT: br_223 
* OUTPUT: bl_224 
* OUTPUT: br_224 
* OUTPUT: bl_225 
* OUTPUT: br_225 
* OUTPUT: bl_226 
* OUTPUT: br_226 
* OUTPUT: bl_227 
* OUTPUT: br_227 
* OUTPUT: bl_228 
* OUTPUT: br_228 
* OUTPUT: bl_229 
* OUTPUT: br_229 
* OUTPUT: bl_230 
* OUTPUT: br_230 
* OUTPUT: bl_231 
* OUTPUT: br_231 
* OUTPUT: bl_232 
* OUTPUT: br_232 
* OUTPUT: bl_233 
* OUTPUT: br_233 
* OUTPUT: bl_234 
* OUTPUT: br_234 
* OUTPUT: bl_235 
* OUTPUT: br_235 
* OUTPUT: bl_236 
* OUTPUT: br_236 
* OUTPUT: bl_237 
* OUTPUT: br_237 
* OUTPUT: bl_238 
* OUTPUT: br_238 
* OUTPUT: bl_239 
* OUTPUT: br_239 
* OUTPUT: bl_240 
* OUTPUT: br_240 
* OUTPUT: bl_241 
* OUTPUT: br_241 
* OUTPUT: bl_242 
* OUTPUT: br_242 
* OUTPUT: bl_243 
* OUTPUT: br_243 
* OUTPUT: bl_244 
* OUTPUT: br_244 
* OUTPUT: bl_245 
* OUTPUT: br_245 
* OUTPUT: bl_246 
* OUTPUT: br_246 
* OUTPUT: bl_247 
* OUTPUT: br_247 
* OUTPUT: bl_248 
* OUTPUT: br_248 
* OUTPUT: bl_249 
* OUTPUT: br_249 
* OUTPUT: bl_250 
* OUTPUT: br_250 
* OUTPUT: bl_251 
* OUTPUT: br_251 
* OUTPUT: bl_252 
* OUTPUT: br_252 
* OUTPUT: bl_253 
* OUTPUT: br_253 
* OUTPUT: bl_254 
* OUTPUT: br_254 
* OUTPUT: bl_255 
* OUTPUT: br_255 
* OUTPUT: bl_256 
* OUTPUT: br_256 
* OUTPUT: bl_257 
* OUTPUT: br_257 
* OUTPUT: bl_258 
* OUTPUT: br_258 
* OUTPUT: bl_259 
* OUTPUT: br_259 
* OUTPUT: bl_260 
* OUTPUT: br_260 
* OUTPUT: bl_261 
* OUTPUT: br_261 
* OUTPUT: bl_262 
* OUTPUT: br_262 
* OUTPUT: bl_263 
* OUTPUT: br_263 
* OUTPUT: bl_264 
* OUTPUT: br_264 
* OUTPUT: bl_265 
* OUTPUT: br_265 
* OUTPUT: bl_266 
* OUTPUT: br_266 
* OUTPUT: bl_267 
* OUTPUT: br_267 
* OUTPUT: bl_268 
* OUTPUT: br_268 
* OUTPUT: bl_269 
* OUTPUT: br_269 
* OUTPUT: bl_270 
* OUTPUT: br_270 
* OUTPUT: bl_271 
* OUTPUT: br_271 
* OUTPUT: bl_272 
* OUTPUT: br_272 
* OUTPUT: bl_273 
* OUTPUT: br_273 
* OUTPUT: bl_274 
* OUTPUT: br_274 
* OUTPUT: bl_275 
* OUTPUT: br_275 
* OUTPUT: bl_276 
* OUTPUT: br_276 
* OUTPUT: bl_277 
* OUTPUT: br_277 
* OUTPUT: bl_278 
* OUTPUT: br_278 
* OUTPUT: bl_279 
* OUTPUT: br_279 
* OUTPUT: bl_280 
* OUTPUT: br_280 
* OUTPUT: bl_281 
* OUTPUT: br_281 
* OUTPUT: bl_282 
* OUTPUT: br_282 
* OUTPUT: bl_283 
* OUTPUT: br_283 
* OUTPUT: bl_284 
* OUTPUT: br_284 
* OUTPUT: bl_285 
* OUTPUT: br_285 
* OUTPUT: bl_286 
* OUTPUT: br_286 
* OUTPUT: bl_287 
* OUTPUT: br_287 
* OUTPUT: bl_288 
* OUTPUT: br_288 
* OUTPUT: bl_289 
* OUTPUT: br_289 
* OUTPUT: bl_290 
* OUTPUT: br_290 
* OUTPUT: bl_291 
* OUTPUT: br_291 
* OUTPUT: bl_292 
* OUTPUT: br_292 
* OUTPUT: bl_293 
* OUTPUT: br_293 
* OUTPUT: bl_294 
* OUTPUT: br_294 
* OUTPUT: bl_295 
* OUTPUT: br_295 
* OUTPUT: bl_296 
* OUTPUT: br_296 
* OUTPUT: bl_297 
* OUTPUT: br_297 
* OUTPUT: bl_298 
* OUTPUT: br_298 
* OUTPUT: bl_299 
* OUTPUT: br_299 
* OUTPUT: bl_300 
* OUTPUT: br_300 
* OUTPUT: bl_301 
* OUTPUT: br_301 
* OUTPUT: bl_302 
* OUTPUT: br_302 
* OUTPUT: bl_303 
* OUTPUT: br_303 
* OUTPUT: bl_304 
* OUTPUT: br_304 
* OUTPUT: bl_305 
* OUTPUT: br_305 
* OUTPUT: bl_306 
* OUTPUT: br_306 
* OUTPUT: bl_307 
* OUTPUT: br_307 
* OUTPUT: bl_308 
* OUTPUT: br_308 
* OUTPUT: bl_309 
* OUTPUT: br_309 
* OUTPUT: bl_310 
* OUTPUT: br_310 
* OUTPUT: bl_311 
* OUTPUT: br_311 
* OUTPUT: bl_312 
* OUTPUT: br_312 
* OUTPUT: bl_313 
* OUTPUT: br_313 
* OUTPUT: bl_314 
* OUTPUT: br_314 
* OUTPUT: bl_315 
* OUTPUT: br_315 
* OUTPUT: bl_316 
* OUTPUT: br_316 
* OUTPUT: bl_317 
* OUTPUT: br_317 
* OUTPUT: bl_318 
* OUTPUT: br_318 
* OUTPUT: bl_319 
* OUTPUT: br_319 
* OUTPUT: bl_320 
* OUTPUT: br_320 
* OUTPUT: bl_321 
* OUTPUT: br_321 
* OUTPUT: bl_322 
* OUTPUT: br_322 
* OUTPUT: bl_323 
* OUTPUT: br_323 
* OUTPUT: bl_324 
* OUTPUT: br_324 
* OUTPUT: bl_325 
* OUTPUT: br_325 
* OUTPUT: bl_326 
* OUTPUT: br_326 
* OUTPUT: bl_327 
* OUTPUT: br_327 
* OUTPUT: bl_328 
* OUTPUT: br_328 
* OUTPUT: bl_329 
* OUTPUT: br_329 
* OUTPUT: bl_330 
* OUTPUT: br_330 
* OUTPUT: bl_331 
* OUTPUT: br_331 
* OUTPUT: bl_332 
* OUTPUT: br_332 
* OUTPUT: bl_333 
* OUTPUT: br_333 
* OUTPUT: bl_334 
* OUTPUT: br_334 
* OUTPUT: bl_335 
* OUTPUT: br_335 
* OUTPUT: bl_336 
* OUTPUT: br_336 
* OUTPUT: bl_337 
* OUTPUT: br_337 
* OUTPUT: bl_338 
* OUTPUT: br_338 
* OUTPUT: bl_339 
* OUTPUT: br_339 
* OUTPUT: bl_340 
* OUTPUT: br_340 
* OUTPUT: bl_341 
* OUTPUT: br_341 
* OUTPUT: bl_342 
* OUTPUT: br_342 
* OUTPUT: bl_343 
* OUTPUT: br_343 
* OUTPUT: bl_344 
* OUTPUT: br_344 
* OUTPUT: bl_345 
* OUTPUT: br_345 
* OUTPUT: bl_346 
* OUTPUT: br_346 
* OUTPUT: bl_347 
* OUTPUT: br_347 
* OUTPUT: bl_348 
* OUTPUT: br_348 
* OUTPUT: bl_349 
* OUTPUT: br_349 
* OUTPUT: bl_350 
* OUTPUT: br_350 
* OUTPUT: bl_351 
* OUTPUT: br_351 
* OUTPUT: bl_352 
* OUTPUT: br_352 
* OUTPUT: bl_353 
* OUTPUT: br_353 
* OUTPUT: bl_354 
* OUTPUT: br_354 
* OUTPUT: bl_355 
* OUTPUT: br_355 
* OUTPUT: bl_356 
* OUTPUT: br_356 
* OUTPUT: bl_357 
* OUTPUT: br_357 
* OUTPUT: bl_358 
* OUTPUT: br_358 
* OUTPUT: bl_359 
* OUTPUT: br_359 
* OUTPUT: bl_360 
* OUTPUT: br_360 
* OUTPUT: bl_361 
* OUTPUT: br_361 
* OUTPUT: bl_362 
* OUTPUT: br_362 
* OUTPUT: bl_363 
* OUTPUT: br_363 
* OUTPUT: bl_364 
* OUTPUT: br_364 
* OUTPUT: bl_365 
* OUTPUT: br_365 
* OUTPUT: bl_366 
* OUTPUT: br_366 
* OUTPUT: bl_367 
* OUTPUT: br_367 
* OUTPUT: bl_368 
* OUTPUT: br_368 
* OUTPUT: bl_369 
* OUTPUT: br_369 
* OUTPUT: bl_370 
* OUTPUT: br_370 
* OUTPUT: bl_371 
* OUTPUT: br_371 
* OUTPUT: bl_372 
* OUTPUT: br_372 
* OUTPUT: bl_373 
* OUTPUT: br_373 
* OUTPUT: bl_374 
* OUTPUT: br_374 
* OUTPUT: bl_375 
* OUTPUT: br_375 
* OUTPUT: bl_376 
* OUTPUT: br_376 
* OUTPUT: bl_377 
* OUTPUT: br_377 
* OUTPUT: bl_378 
* OUTPUT: br_378 
* OUTPUT: bl_379 
* OUTPUT: br_379 
* OUTPUT: bl_380 
* OUTPUT: br_380 
* OUTPUT: bl_381 
* OUTPUT: br_381 
* OUTPUT: bl_382 
* OUTPUT: br_382 
* OUTPUT: bl_383 
* OUTPUT: br_383 
* OUTPUT: bl_384 
* OUTPUT: br_384 
* OUTPUT: bl_385 
* OUTPUT: br_385 
* OUTPUT: bl_386 
* OUTPUT: br_386 
* OUTPUT: bl_387 
* OUTPUT: br_387 
* OUTPUT: bl_388 
* OUTPUT: br_388 
* OUTPUT: bl_389 
* OUTPUT: br_389 
* OUTPUT: bl_390 
* OUTPUT: br_390 
* OUTPUT: bl_391 
* OUTPUT: br_391 
* OUTPUT: bl_392 
* OUTPUT: br_392 
* OUTPUT: bl_393 
* OUTPUT: br_393 
* OUTPUT: bl_394 
* OUTPUT: br_394 
* OUTPUT: bl_395 
* OUTPUT: br_395 
* OUTPUT: bl_396 
* OUTPUT: br_396 
* OUTPUT: bl_397 
* OUTPUT: br_397 
* OUTPUT: bl_398 
* OUTPUT: br_398 
* OUTPUT: bl_399 
* OUTPUT: br_399 
* OUTPUT: bl_400 
* OUTPUT: br_400 
* OUTPUT: bl_401 
* OUTPUT: br_401 
* OUTPUT: bl_402 
* OUTPUT: br_402 
* OUTPUT: bl_403 
* OUTPUT: br_403 
* OUTPUT: bl_404 
* OUTPUT: br_404 
* OUTPUT: bl_405 
* OUTPUT: br_405 
* OUTPUT: bl_406 
* OUTPUT: br_406 
* OUTPUT: bl_407 
* OUTPUT: br_407 
* OUTPUT: bl_408 
* OUTPUT: br_408 
* OUTPUT: bl_409 
* OUTPUT: br_409 
* OUTPUT: bl_410 
* OUTPUT: br_410 
* OUTPUT: bl_411 
* OUTPUT: br_411 
* OUTPUT: bl_412 
* OUTPUT: br_412 
* OUTPUT: bl_413 
* OUTPUT: br_413 
* OUTPUT: bl_414 
* OUTPUT: br_414 
* OUTPUT: bl_415 
* OUTPUT: br_415 
* OUTPUT: bl_416 
* OUTPUT: br_416 
* OUTPUT: bl_417 
* OUTPUT: br_417 
* OUTPUT: bl_418 
* OUTPUT: br_418 
* OUTPUT: bl_419 
* OUTPUT: br_419 
* OUTPUT: bl_420 
* OUTPUT: br_420 
* OUTPUT: bl_421 
* OUTPUT: br_421 
* OUTPUT: bl_422 
* OUTPUT: br_422 
* OUTPUT: bl_423 
* OUTPUT: br_423 
* OUTPUT: bl_424 
* OUTPUT: br_424 
* OUTPUT: bl_425 
* OUTPUT: br_425 
* OUTPUT: bl_426 
* OUTPUT: br_426 
* OUTPUT: bl_427 
* OUTPUT: br_427 
* OUTPUT: bl_428 
* OUTPUT: br_428 
* OUTPUT: bl_429 
* OUTPUT: br_429 
* OUTPUT: bl_430 
* OUTPUT: br_430 
* OUTPUT: bl_431 
* OUTPUT: br_431 
* OUTPUT: bl_432 
* OUTPUT: br_432 
* OUTPUT: bl_433 
* OUTPUT: br_433 
* OUTPUT: bl_434 
* OUTPUT: br_434 
* OUTPUT: bl_435 
* OUTPUT: br_435 
* OUTPUT: bl_436 
* OUTPUT: br_436 
* OUTPUT: bl_437 
* OUTPUT: br_437 
* OUTPUT: bl_438 
* OUTPUT: br_438 
* OUTPUT: bl_439 
* OUTPUT: br_439 
* OUTPUT: bl_440 
* OUTPUT: br_440 
* OUTPUT: bl_441 
* OUTPUT: br_441 
* OUTPUT: bl_442 
* OUTPUT: br_442 
* OUTPUT: bl_443 
* OUTPUT: br_443 
* OUTPUT: bl_444 
* OUTPUT: br_444 
* OUTPUT: bl_445 
* OUTPUT: br_445 
* OUTPUT: bl_446 
* OUTPUT: br_446 
* OUTPUT: bl_447 
* OUTPUT: br_447 
* OUTPUT: bl_448 
* OUTPUT: br_448 
* OUTPUT: bl_449 
* OUTPUT: br_449 
* OUTPUT: bl_450 
* OUTPUT: br_450 
* OUTPUT: bl_451 
* OUTPUT: br_451 
* OUTPUT: bl_452 
* OUTPUT: br_452 
* OUTPUT: bl_453 
* OUTPUT: br_453 
* OUTPUT: bl_454 
* OUTPUT: br_454 
* OUTPUT: bl_455 
* OUTPUT: br_455 
* OUTPUT: bl_456 
* OUTPUT: br_456 
* OUTPUT: bl_457 
* OUTPUT: br_457 
* OUTPUT: bl_458 
* OUTPUT: br_458 
* OUTPUT: bl_459 
* OUTPUT: br_459 
* OUTPUT: bl_460 
* OUTPUT: br_460 
* OUTPUT: bl_461 
* OUTPUT: br_461 
* OUTPUT: bl_462 
* OUTPUT: br_462 
* OUTPUT: bl_463 
* OUTPUT: br_463 
* OUTPUT: bl_464 
* OUTPUT: br_464 
* OUTPUT: bl_465 
* OUTPUT: br_465 
* OUTPUT: bl_466 
* OUTPUT: br_466 
* OUTPUT: bl_467 
* OUTPUT: br_467 
* OUTPUT: bl_468 
* OUTPUT: br_468 
* OUTPUT: bl_469 
* OUTPUT: br_469 
* OUTPUT: bl_470 
* OUTPUT: br_470 
* OUTPUT: bl_471 
* OUTPUT: br_471 
* OUTPUT: bl_472 
* OUTPUT: br_472 
* OUTPUT: bl_473 
* OUTPUT: br_473 
* OUTPUT: bl_474 
* OUTPUT: br_474 
* OUTPUT: bl_475 
* OUTPUT: br_475 
* OUTPUT: bl_476 
* OUTPUT: br_476 
* OUTPUT: bl_477 
* OUTPUT: br_477 
* OUTPUT: bl_478 
* OUTPUT: br_478 
* OUTPUT: bl_479 
* OUTPUT: br_479 
* OUTPUT: bl_480 
* OUTPUT: br_480 
* OUTPUT: bl_481 
* OUTPUT: br_481 
* OUTPUT: bl_482 
* OUTPUT: br_482 
* OUTPUT: bl_483 
* OUTPUT: br_483 
* OUTPUT: bl_484 
* OUTPUT: br_484 
* OUTPUT: bl_485 
* OUTPUT: br_485 
* OUTPUT: bl_486 
* OUTPUT: br_486 
* OUTPUT: bl_487 
* OUTPUT: br_487 
* OUTPUT: bl_488 
* OUTPUT: br_488 
* OUTPUT: bl_489 
* OUTPUT: br_489 
* OUTPUT: bl_490 
* OUTPUT: br_490 
* OUTPUT: bl_491 
* OUTPUT: br_491 
* OUTPUT: bl_492 
* OUTPUT: br_492 
* OUTPUT: bl_493 
* OUTPUT: br_493 
* OUTPUT: bl_494 
* OUTPUT: br_494 
* OUTPUT: bl_495 
* OUTPUT: br_495 
* OUTPUT: bl_496 
* OUTPUT: br_496 
* OUTPUT: bl_497 
* OUTPUT: br_497 
* OUTPUT: bl_498 
* OUTPUT: br_498 
* OUTPUT: bl_499 
* OUTPUT: br_499 
* OUTPUT: bl_500 
* OUTPUT: br_500 
* OUTPUT: bl_501 
* OUTPUT: br_501 
* OUTPUT: bl_502 
* OUTPUT: br_502 
* OUTPUT: bl_503 
* OUTPUT: br_503 
* OUTPUT: bl_504 
* OUTPUT: br_504 
* OUTPUT: bl_505 
* OUTPUT: br_505 
* OUTPUT: bl_506 
* OUTPUT: br_506 
* OUTPUT: bl_507 
* OUTPUT: br_507 
* OUTPUT: bl_508 
* OUTPUT: br_508 
* OUTPUT: bl_509 
* OUTPUT: br_509 
* OUTPUT: bl_510 
* OUTPUT: br_510 
* OUTPUT: bl_511 
* OUTPUT: br_511 
* OUTPUT: bl_512 
* OUTPUT: br_512 
* INPUT : en_bar 
* POWER : vdd 
* cols: 513 size: 1 bl: bl br: br
Xpre_column_0
+ bl_0 br_0 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_1
+ bl_1 br_1 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_2
+ bl_2 br_2 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_3
+ bl_3 br_3 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_4
+ bl_4 br_4 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_5
+ bl_5 br_5 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_6
+ bl_6 br_6 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_7
+ bl_7 br_7 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_8
+ bl_8 br_8 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_9
+ bl_9 br_9 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_10
+ bl_10 br_10 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_11
+ bl_11 br_11 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_12
+ bl_12 br_12 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_13
+ bl_13 br_13 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_14
+ bl_14 br_14 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_15
+ bl_15 br_15 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_16
+ bl_16 br_16 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_17
+ bl_17 br_17 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_18
+ bl_18 br_18 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_19
+ bl_19 br_19 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_20
+ bl_20 br_20 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_21
+ bl_21 br_21 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_22
+ bl_22 br_22 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_23
+ bl_23 br_23 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_24
+ bl_24 br_24 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_25
+ bl_25 br_25 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_26
+ bl_26 br_26 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_27
+ bl_27 br_27 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_28
+ bl_28 br_28 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_29
+ bl_29 br_29 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_30
+ bl_30 br_30 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_31
+ bl_31 br_31 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_32
+ bl_32 br_32 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_33
+ bl_33 br_33 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_34
+ bl_34 br_34 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_35
+ bl_35 br_35 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_36
+ bl_36 br_36 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_37
+ bl_37 br_37 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_38
+ bl_38 br_38 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_39
+ bl_39 br_39 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_40
+ bl_40 br_40 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_41
+ bl_41 br_41 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_42
+ bl_42 br_42 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_43
+ bl_43 br_43 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_44
+ bl_44 br_44 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_45
+ bl_45 br_45 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_46
+ bl_46 br_46 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_47
+ bl_47 br_47 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_48
+ bl_48 br_48 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_49
+ bl_49 br_49 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_50
+ bl_50 br_50 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_51
+ bl_51 br_51 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_52
+ bl_52 br_52 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_53
+ bl_53 br_53 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_54
+ bl_54 br_54 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_55
+ bl_55 br_55 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_56
+ bl_56 br_56 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_57
+ bl_57 br_57 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_58
+ bl_58 br_58 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_59
+ bl_59 br_59 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_60
+ bl_60 br_60 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_61
+ bl_61 br_61 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_62
+ bl_62 br_62 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_63
+ bl_63 br_63 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_64
+ bl_64 br_64 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_65
+ bl_65 br_65 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_66
+ bl_66 br_66 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_67
+ bl_67 br_67 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_68
+ bl_68 br_68 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_69
+ bl_69 br_69 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_70
+ bl_70 br_70 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_71
+ bl_71 br_71 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_72
+ bl_72 br_72 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_73
+ bl_73 br_73 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_74
+ bl_74 br_74 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_75
+ bl_75 br_75 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_76
+ bl_76 br_76 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_77
+ bl_77 br_77 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_78
+ bl_78 br_78 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_79
+ bl_79 br_79 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_80
+ bl_80 br_80 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_81
+ bl_81 br_81 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_82
+ bl_82 br_82 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_83
+ bl_83 br_83 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_84
+ bl_84 br_84 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_85
+ bl_85 br_85 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_86
+ bl_86 br_86 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_87
+ bl_87 br_87 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_88
+ bl_88 br_88 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_89
+ bl_89 br_89 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_90
+ bl_90 br_90 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_91
+ bl_91 br_91 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_92
+ bl_92 br_92 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_93
+ bl_93 br_93 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_94
+ bl_94 br_94 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_95
+ bl_95 br_95 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_96
+ bl_96 br_96 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_97
+ bl_97 br_97 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_98
+ bl_98 br_98 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_99
+ bl_99 br_99 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_100
+ bl_100 br_100 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_101
+ bl_101 br_101 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_102
+ bl_102 br_102 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_103
+ bl_103 br_103 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_104
+ bl_104 br_104 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_105
+ bl_105 br_105 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_106
+ bl_106 br_106 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_107
+ bl_107 br_107 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_108
+ bl_108 br_108 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_109
+ bl_109 br_109 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_110
+ bl_110 br_110 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_111
+ bl_111 br_111 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_112
+ bl_112 br_112 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_113
+ bl_113 br_113 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_114
+ bl_114 br_114 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_115
+ bl_115 br_115 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_116
+ bl_116 br_116 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_117
+ bl_117 br_117 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_118
+ bl_118 br_118 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_119
+ bl_119 br_119 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_120
+ bl_120 br_120 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_121
+ bl_121 br_121 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_122
+ bl_122 br_122 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_123
+ bl_123 br_123 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_124
+ bl_124 br_124 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_125
+ bl_125 br_125 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_126
+ bl_126 br_126 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_127
+ bl_127 br_127 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_128
+ bl_128 br_128 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_129
+ bl_129 br_129 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_130
+ bl_130 br_130 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_131
+ bl_131 br_131 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_132
+ bl_132 br_132 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_133
+ bl_133 br_133 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_134
+ bl_134 br_134 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_135
+ bl_135 br_135 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_136
+ bl_136 br_136 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_137
+ bl_137 br_137 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_138
+ bl_138 br_138 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_139
+ bl_139 br_139 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_140
+ bl_140 br_140 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_141
+ bl_141 br_141 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_142
+ bl_142 br_142 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_143
+ bl_143 br_143 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_144
+ bl_144 br_144 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_145
+ bl_145 br_145 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_146
+ bl_146 br_146 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_147
+ bl_147 br_147 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_148
+ bl_148 br_148 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_149
+ bl_149 br_149 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_150
+ bl_150 br_150 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_151
+ bl_151 br_151 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_152
+ bl_152 br_152 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_153
+ bl_153 br_153 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_154
+ bl_154 br_154 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_155
+ bl_155 br_155 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_156
+ bl_156 br_156 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_157
+ bl_157 br_157 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_158
+ bl_158 br_158 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_159
+ bl_159 br_159 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_160
+ bl_160 br_160 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_161
+ bl_161 br_161 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_162
+ bl_162 br_162 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_163
+ bl_163 br_163 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_164
+ bl_164 br_164 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_165
+ bl_165 br_165 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_166
+ bl_166 br_166 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_167
+ bl_167 br_167 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_168
+ bl_168 br_168 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_169
+ bl_169 br_169 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_170
+ bl_170 br_170 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_171
+ bl_171 br_171 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_172
+ bl_172 br_172 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_173
+ bl_173 br_173 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_174
+ bl_174 br_174 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_175
+ bl_175 br_175 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_176
+ bl_176 br_176 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_177
+ bl_177 br_177 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_178
+ bl_178 br_178 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_179
+ bl_179 br_179 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_180
+ bl_180 br_180 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_181
+ bl_181 br_181 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_182
+ bl_182 br_182 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_183
+ bl_183 br_183 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_184
+ bl_184 br_184 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_185
+ bl_185 br_185 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_186
+ bl_186 br_186 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_187
+ bl_187 br_187 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_188
+ bl_188 br_188 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_189
+ bl_189 br_189 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_190
+ bl_190 br_190 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_191
+ bl_191 br_191 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_192
+ bl_192 br_192 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_193
+ bl_193 br_193 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_194
+ bl_194 br_194 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_195
+ bl_195 br_195 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_196
+ bl_196 br_196 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_197
+ bl_197 br_197 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_198
+ bl_198 br_198 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_199
+ bl_199 br_199 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_200
+ bl_200 br_200 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_201
+ bl_201 br_201 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_202
+ bl_202 br_202 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_203
+ bl_203 br_203 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_204
+ bl_204 br_204 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_205
+ bl_205 br_205 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_206
+ bl_206 br_206 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_207
+ bl_207 br_207 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_208
+ bl_208 br_208 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_209
+ bl_209 br_209 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_210
+ bl_210 br_210 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_211
+ bl_211 br_211 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_212
+ bl_212 br_212 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_213
+ bl_213 br_213 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_214
+ bl_214 br_214 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_215
+ bl_215 br_215 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_216
+ bl_216 br_216 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_217
+ bl_217 br_217 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_218
+ bl_218 br_218 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_219
+ bl_219 br_219 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_220
+ bl_220 br_220 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_221
+ bl_221 br_221 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_222
+ bl_222 br_222 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_223
+ bl_223 br_223 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_224
+ bl_224 br_224 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_225
+ bl_225 br_225 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_226
+ bl_226 br_226 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_227
+ bl_227 br_227 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_228
+ bl_228 br_228 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_229
+ bl_229 br_229 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_230
+ bl_230 br_230 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_231
+ bl_231 br_231 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_232
+ bl_232 br_232 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_233
+ bl_233 br_233 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_234
+ bl_234 br_234 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_235
+ bl_235 br_235 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_236
+ bl_236 br_236 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_237
+ bl_237 br_237 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_238
+ bl_238 br_238 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_239
+ bl_239 br_239 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_240
+ bl_240 br_240 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_241
+ bl_241 br_241 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_242
+ bl_242 br_242 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_243
+ bl_243 br_243 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_244
+ bl_244 br_244 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_245
+ bl_245 br_245 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_246
+ bl_246 br_246 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_247
+ bl_247 br_247 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_248
+ bl_248 br_248 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_249
+ bl_249 br_249 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_250
+ bl_250 br_250 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_251
+ bl_251 br_251 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_252
+ bl_252 br_252 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_253
+ bl_253 br_253 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_254
+ bl_254 br_254 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_255
+ bl_255 br_255 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_256
+ bl_256 br_256 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_257
+ bl_257 br_257 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_258
+ bl_258 br_258 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_259
+ bl_259 br_259 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_260
+ bl_260 br_260 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_261
+ bl_261 br_261 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_262
+ bl_262 br_262 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_263
+ bl_263 br_263 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_264
+ bl_264 br_264 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_265
+ bl_265 br_265 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_266
+ bl_266 br_266 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_267
+ bl_267 br_267 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_268
+ bl_268 br_268 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_269
+ bl_269 br_269 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_270
+ bl_270 br_270 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_271
+ bl_271 br_271 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_272
+ bl_272 br_272 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_273
+ bl_273 br_273 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_274
+ bl_274 br_274 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_275
+ bl_275 br_275 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_276
+ bl_276 br_276 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_277
+ bl_277 br_277 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_278
+ bl_278 br_278 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_279
+ bl_279 br_279 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_280
+ bl_280 br_280 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_281
+ bl_281 br_281 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_282
+ bl_282 br_282 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_283
+ bl_283 br_283 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_284
+ bl_284 br_284 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_285
+ bl_285 br_285 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_286
+ bl_286 br_286 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_287
+ bl_287 br_287 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_288
+ bl_288 br_288 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_289
+ bl_289 br_289 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_290
+ bl_290 br_290 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_291
+ bl_291 br_291 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_292
+ bl_292 br_292 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_293
+ bl_293 br_293 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_294
+ bl_294 br_294 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_295
+ bl_295 br_295 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_296
+ bl_296 br_296 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_297
+ bl_297 br_297 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_298
+ bl_298 br_298 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_299
+ bl_299 br_299 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_300
+ bl_300 br_300 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_301
+ bl_301 br_301 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_302
+ bl_302 br_302 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_303
+ bl_303 br_303 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_304
+ bl_304 br_304 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_305
+ bl_305 br_305 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_306
+ bl_306 br_306 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_307
+ bl_307 br_307 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_308
+ bl_308 br_308 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_309
+ bl_309 br_309 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_310
+ bl_310 br_310 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_311
+ bl_311 br_311 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_312
+ bl_312 br_312 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_313
+ bl_313 br_313 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_314
+ bl_314 br_314 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_315
+ bl_315 br_315 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_316
+ bl_316 br_316 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_317
+ bl_317 br_317 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_318
+ bl_318 br_318 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_319
+ bl_319 br_319 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_320
+ bl_320 br_320 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_321
+ bl_321 br_321 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_322
+ bl_322 br_322 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_323
+ bl_323 br_323 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_324
+ bl_324 br_324 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_325
+ bl_325 br_325 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_326
+ bl_326 br_326 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_327
+ bl_327 br_327 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_328
+ bl_328 br_328 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_329
+ bl_329 br_329 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_330
+ bl_330 br_330 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_331
+ bl_331 br_331 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_332
+ bl_332 br_332 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_333
+ bl_333 br_333 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_334
+ bl_334 br_334 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_335
+ bl_335 br_335 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_336
+ bl_336 br_336 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_337
+ bl_337 br_337 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_338
+ bl_338 br_338 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_339
+ bl_339 br_339 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_340
+ bl_340 br_340 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_341
+ bl_341 br_341 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_342
+ bl_342 br_342 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_343
+ bl_343 br_343 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_344
+ bl_344 br_344 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_345
+ bl_345 br_345 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_346
+ bl_346 br_346 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_347
+ bl_347 br_347 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_348
+ bl_348 br_348 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_349
+ bl_349 br_349 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_350
+ bl_350 br_350 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_351
+ bl_351 br_351 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_352
+ bl_352 br_352 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_353
+ bl_353 br_353 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_354
+ bl_354 br_354 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_355
+ bl_355 br_355 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_356
+ bl_356 br_356 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_357
+ bl_357 br_357 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_358
+ bl_358 br_358 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_359
+ bl_359 br_359 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_360
+ bl_360 br_360 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_361
+ bl_361 br_361 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_362
+ bl_362 br_362 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_363
+ bl_363 br_363 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_364
+ bl_364 br_364 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_365
+ bl_365 br_365 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_366
+ bl_366 br_366 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_367
+ bl_367 br_367 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_368
+ bl_368 br_368 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_369
+ bl_369 br_369 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_370
+ bl_370 br_370 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_371
+ bl_371 br_371 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_372
+ bl_372 br_372 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_373
+ bl_373 br_373 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_374
+ bl_374 br_374 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_375
+ bl_375 br_375 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_376
+ bl_376 br_376 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_377
+ bl_377 br_377 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_378
+ bl_378 br_378 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_379
+ bl_379 br_379 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_380
+ bl_380 br_380 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_381
+ bl_381 br_381 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_382
+ bl_382 br_382 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_383
+ bl_383 br_383 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_384
+ bl_384 br_384 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_385
+ bl_385 br_385 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_386
+ bl_386 br_386 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_387
+ bl_387 br_387 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_388
+ bl_388 br_388 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_389
+ bl_389 br_389 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_390
+ bl_390 br_390 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_391
+ bl_391 br_391 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_392
+ bl_392 br_392 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_393
+ bl_393 br_393 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_394
+ bl_394 br_394 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_395
+ bl_395 br_395 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_396
+ bl_396 br_396 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_397
+ bl_397 br_397 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_398
+ bl_398 br_398 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_399
+ bl_399 br_399 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_400
+ bl_400 br_400 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_401
+ bl_401 br_401 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_402
+ bl_402 br_402 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_403
+ bl_403 br_403 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_404
+ bl_404 br_404 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_405
+ bl_405 br_405 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_406
+ bl_406 br_406 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_407
+ bl_407 br_407 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_408
+ bl_408 br_408 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_409
+ bl_409 br_409 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_410
+ bl_410 br_410 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_411
+ bl_411 br_411 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_412
+ bl_412 br_412 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_413
+ bl_413 br_413 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_414
+ bl_414 br_414 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_415
+ bl_415 br_415 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_416
+ bl_416 br_416 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_417
+ bl_417 br_417 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_418
+ bl_418 br_418 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_419
+ bl_419 br_419 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_420
+ bl_420 br_420 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_421
+ bl_421 br_421 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_422
+ bl_422 br_422 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_423
+ bl_423 br_423 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_424
+ bl_424 br_424 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_425
+ bl_425 br_425 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_426
+ bl_426 br_426 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_427
+ bl_427 br_427 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_428
+ bl_428 br_428 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_429
+ bl_429 br_429 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_430
+ bl_430 br_430 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_431
+ bl_431 br_431 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_432
+ bl_432 br_432 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_433
+ bl_433 br_433 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_434
+ bl_434 br_434 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_435
+ bl_435 br_435 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_436
+ bl_436 br_436 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_437
+ bl_437 br_437 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_438
+ bl_438 br_438 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_439
+ bl_439 br_439 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_440
+ bl_440 br_440 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_441
+ bl_441 br_441 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_442
+ bl_442 br_442 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_443
+ bl_443 br_443 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_444
+ bl_444 br_444 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_445
+ bl_445 br_445 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_446
+ bl_446 br_446 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_447
+ bl_447 br_447 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_448
+ bl_448 br_448 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_449
+ bl_449 br_449 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_450
+ bl_450 br_450 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_451
+ bl_451 br_451 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_452
+ bl_452 br_452 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_453
+ bl_453 br_453 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_454
+ bl_454 br_454 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_455
+ bl_455 br_455 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_456
+ bl_456 br_456 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_457
+ bl_457 br_457 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_458
+ bl_458 br_458 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_459
+ bl_459 br_459 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_460
+ bl_460 br_460 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_461
+ bl_461 br_461 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_462
+ bl_462 br_462 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_463
+ bl_463 br_463 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_464
+ bl_464 br_464 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_465
+ bl_465 br_465 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_466
+ bl_466 br_466 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_467
+ bl_467 br_467 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_468
+ bl_468 br_468 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_469
+ bl_469 br_469 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_470
+ bl_470 br_470 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_471
+ bl_471 br_471 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_472
+ bl_472 br_472 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_473
+ bl_473 br_473 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_474
+ bl_474 br_474 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_475
+ bl_475 br_475 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_476
+ bl_476 br_476 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_477
+ bl_477 br_477 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_478
+ bl_478 br_478 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_479
+ bl_479 br_479 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_480
+ bl_480 br_480 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_481
+ bl_481 br_481 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_482
+ bl_482 br_482 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_483
+ bl_483 br_483 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_484
+ bl_484 br_484 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_485
+ bl_485 br_485 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_486
+ bl_486 br_486 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_487
+ bl_487 br_487 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_488
+ bl_488 br_488 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_489
+ bl_489 br_489 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_490
+ bl_490 br_490 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_491
+ bl_491 br_491 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_492
+ bl_492 br_492 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_493
+ bl_493 br_493 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_494
+ bl_494 br_494 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_495
+ bl_495 br_495 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_496
+ bl_496 br_496 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_497
+ bl_497 br_497 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_498
+ bl_498 br_498 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_499
+ bl_499 br_499 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_500
+ bl_500 br_500 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_501
+ bl_501 br_501 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_502
+ bl_502 br_502 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_503
+ bl_503 br_503 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_504
+ bl_504 br_504 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_505
+ bl_505 br_505 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_506
+ bl_506 br_506 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_507
+ bl_507 br_507 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_508
+ bl_508 br_508 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_509
+ bl_509 br_509 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_510
+ bl_510 br_510 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_511
+ bl_511 br_511 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
Xpre_column_512
+ bl_512 br_512 en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_0
.ENDS freepdk45_sram_1rw0r_45x512_precharge_array

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dout vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dout net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dout net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dout vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp


.SUBCKT freepdk45_sram_1rw0r_45x512_sense_amp_array
+ data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3
+ data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7
+ data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11
+ br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14
+ data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18
+ bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21
+ br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24
+ data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28
+ bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31
+ br_31 data_32 bl_32 br_32 data_33 bl_33 br_33 data_34 bl_34 br_34
+ data_35 bl_35 br_35 data_36 bl_36 br_36 data_37 bl_37 br_37 data_38
+ bl_38 br_38 data_39 bl_39 br_39 data_40 bl_40 br_40 data_41 bl_41
+ br_41 data_42 bl_42 br_42 data_43 bl_43 br_43 data_44 bl_44 br_44
+ data_45 bl_45 br_45 data_46 bl_46 br_46 data_47 bl_47 br_47 data_48
+ bl_48 br_48 data_49 bl_49 br_49 data_50 bl_50 br_50 data_51 bl_51
+ br_51 data_52 bl_52 br_52 data_53 bl_53 br_53 data_54 bl_54 br_54
+ data_55 bl_55 br_55 data_56 bl_56 br_56 data_57 bl_57 br_57 data_58
+ bl_58 br_58 data_59 bl_59 br_59 data_60 bl_60 br_60 data_61 bl_61
+ br_61 data_62 bl_62 br_62 data_63 bl_63 br_63 data_64 bl_64 br_64
+ data_65 bl_65 br_65 data_66 bl_66 br_66 data_67 bl_67 br_67 data_68
+ bl_68 br_68 data_69 bl_69 br_69 data_70 bl_70 br_70 data_71 bl_71
+ br_71 data_72 bl_72 br_72 data_73 bl_73 br_73 data_74 bl_74 br_74
+ data_75 bl_75 br_75 data_76 bl_76 br_76 data_77 bl_77 br_77 data_78
+ bl_78 br_78 data_79 bl_79 br_79 data_80 bl_80 br_80 data_81 bl_81
+ br_81 data_82 bl_82 br_82 data_83 bl_83 br_83 data_84 bl_84 br_84
+ data_85 bl_85 br_85 data_86 bl_86 br_86 data_87 bl_87 br_87 data_88
+ bl_88 br_88 data_89 bl_89 br_89 data_90 bl_90 br_90 data_91 bl_91
+ br_91 data_92 bl_92 br_92 data_93 bl_93 br_93 data_94 bl_94 br_94
+ data_95 bl_95 br_95 data_96 bl_96 br_96 data_97 bl_97 br_97 data_98
+ bl_98 br_98 data_99 bl_99 br_99 data_100 bl_100 br_100 data_101 bl_101
+ br_101 data_102 bl_102 br_102 data_103 bl_103 br_103 data_104 bl_104
+ br_104 data_105 bl_105 br_105 data_106 bl_106 br_106 data_107 bl_107
+ br_107 data_108 bl_108 br_108 data_109 bl_109 br_109 data_110 bl_110
+ br_110 data_111 bl_111 br_111 data_112 bl_112 br_112 data_113 bl_113
+ br_113 data_114 bl_114 br_114 data_115 bl_115 br_115 data_116 bl_116
+ br_116 data_117 bl_117 br_117 data_118 bl_118 br_118 data_119 bl_119
+ br_119 data_120 bl_120 br_120 data_121 bl_121 br_121 data_122 bl_122
+ br_122 data_123 bl_123 br_123 data_124 bl_124 br_124 data_125 bl_125
+ br_125 data_126 bl_126 br_126 data_127 bl_127 br_127 data_128 bl_128
+ br_128 data_129 bl_129 br_129 data_130 bl_130 br_130 data_131 bl_131
+ br_131 data_132 bl_132 br_132 data_133 bl_133 br_133 data_134 bl_134
+ br_134 data_135 bl_135 br_135 data_136 bl_136 br_136 data_137 bl_137
+ br_137 data_138 bl_138 br_138 data_139 bl_139 br_139 data_140 bl_140
+ br_140 data_141 bl_141 br_141 data_142 bl_142 br_142 data_143 bl_143
+ br_143 data_144 bl_144 br_144 data_145 bl_145 br_145 data_146 bl_146
+ br_146 data_147 bl_147 br_147 data_148 bl_148 br_148 data_149 bl_149
+ br_149 data_150 bl_150 br_150 data_151 bl_151 br_151 data_152 bl_152
+ br_152 data_153 bl_153 br_153 data_154 bl_154 br_154 data_155 bl_155
+ br_155 data_156 bl_156 br_156 data_157 bl_157 br_157 data_158 bl_158
+ br_158 data_159 bl_159 br_159 data_160 bl_160 br_160 data_161 bl_161
+ br_161 data_162 bl_162 br_162 data_163 bl_163 br_163 data_164 bl_164
+ br_164 data_165 bl_165 br_165 data_166 bl_166 br_166 data_167 bl_167
+ br_167 data_168 bl_168 br_168 data_169 bl_169 br_169 data_170 bl_170
+ br_170 data_171 bl_171 br_171 data_172 bl_172 br_172 data_173 bl_173
+ br_173 data_174 bl_174 br_174 data_175 bl_175 br_175 data_176 bl_176
+ br_176 data_177 bl_177 br_177 data_178 bl_178 br_178 data_179 bl_179
+ br_179 data_180 bl_180 br_180 data_181 bl_181 br_181 data_182 bl_182
+ br_182 data_183 bl_183 br_183 data_184 bl_184 br_184 data_185 bl_185
+ br_185 data_186 bl_186 br_186 data_187 bl_187 br_187 data_188 bl_188
+ br_188 data_189 bl_189 br_189 data_190 bl_190 br_190 data_191 bl_191
+ br_191 data_192 bl_192 br_192 data_193 bl_193 br_193 data_194 bl_194
+ br_194 data_195 bl_195 br_195 data_196 bl_196 br_196 data_197 bl_197
+ br_197 data_198 bl_198 br_198 data_199 bl_199 br_199 data_200 bl_200
+ br_200 data_201 bl_201 br_201 data_202 bl_202 br_202 data_203 bl_203
+ br_203 data_204 bl_204 br_204 data_205 bl_205 br_205 data_206 bl_206
+ br_206 data_207 bl_207 br_207 data_208 bl_208 br_208 data_209 bl_209
+ br_209 data_210 bl_210 br_210 data_211 bl_211 br_211 data_212 bl_212
+ br_212 data_213 bl_213 br_213 data_214 bl_214 br_214 data_215 bl_215
+ br_215 data_216 bl_216 br_216 data_217 bl_217 br_217 data_218 bl_218
+ br_218 data_219 bl_219 br_219 data_220 bl_220 br_220 data_221 bl_221
+ br_221 data_222 bl_222 br_222 data_223 bl_223 br_223 data_224 bl_224
+ br_224 data_225 bl_225 br_225 data_226 bl_226 br_226 data_227 bl_227
+ br_227 data_228 bl_228 br_228 data_229 bl_229 br_229 data_230 bl_230
+ br_230 data_231 bl_231 br_231 data_232 bl_232 br_232 data_233 bl_233
+ br_233 data_234 bl_234 br_234 data_235 bl_235 br_235 data_236 bl_236
+ br_236 data_237 bl_237 br_237 data_238 bl_238 br_238 data_239 bl_239
+ br_239 data_240 bl_240 br_240 data_241 bl_241 br_241 data_242 bl_242
+ br_242 data_243 bl_243 br_243 data_244 bl_244 br_244 data_245 bl_245
+ br_245 data_246 bl_246 br_246 data_247 bl_247 br_247 data_248 bl_248
+ br_248 data_249 bl_249 br_249 data_250 bl_250 br_250 data_251 bl_251
+ br_251 data_252 bl_252 br_252 data_253 bl_253 br_253 data_254 bl_254
+ br_254 data_255 bl_255 br_255 data_256 bl_256 br_256 data_257 bl_257
+ br_257 data_258 bl_258 br_258 data_259 bl_259 br_259 data_260 bl_260
+ br_260 data_261 bl_261 br_261 data_262 bl_262 br_262 data_263 bl_263
+ br_263 data_264 bl_264 br_264 data_265 bl_265 br_265 data_266 bl_266
+ br_266 data_267 bl_267 br_267 data_268 bl_268 br_268 data_269 bl_269
+ br_269 data_270 bl_270 br_270 data_271 bl_271 br_271 data_272 bl_272
+ br_272 data_273 bl_273 br_273 data_274 bl_274 br_274 data_275 bl_275
+ br_275 data_276 bl_276 br_276 data_277 bl_277 br_277 data_278 bl_278
+ br_278 data_279 bl_279 br_279 data_280 bl_280 br_280 data_281 bl_281
+ br_281 data_282 bl_282 br_282 data_283 bl_283 br_283 data_284 bl_284
+ br_284 data_285 bl_285 br_285 data_286 bl_286 br_286 data_287 bl_287
+ br_287 data_288 bl_288 br_288 data_289 bl_289 br_289 data_290 bl_290
+ br_290 data_291 bl_291 br_291 data_292 bl_292 br_292 data_293 bl_293
+ br_293 data_294 bl_294 br_294 data_295 bl_295 br_295 data_296 bl_296
+ br_296 data_297 bl_297 br_297 data_298 bl_298 br_298 data_299 bl_299
+ br_299 data_300 bl_300 br_300 data_301 bl_301 br_301 data_302 bl_302
+ br_302 data_303 bl_303 br_303 data_304 bl_304 br_304 data_305 bl_305
+ br_305 data_306 bl_306 br_306 data_307 bl_307 br_307 data_308 bl_308
+ br_308 data_309 bl_309 br_309 data_310 bl_310 br_310 data_311 bl_311
+ br_311 data_312 bl_312 br_312 data_313 bl_313 br_313 data_314 bl_314
+ br_314 data_315 bl_315 br_315 data_316 bl_316 br_316 data_317 bl_317
+ br_317 data_318 bl_318 br_318 data_319 bl_319 br_319 data_320 bl_320
+ br_320 data_321 bl_321 br_321 data_322 bl_322 br_322 data_323 bl_323
+ br_323 data_324 bl_324 br_324 data_325 bl_325 br_325 data_326 bl_326
+ br_326 data_327 bl_327 br_327 data_328 bl_328 br_328 data_329 bl_329
+ br_329 data_330 bl_330 br_330 data_331 bl_331 br_331 data_332 bl_332
+ br_332 data_333 bl_333 br_333 data_334 bl_334 br_334 data_335 bl_335
+ br_335 data_336 bl_336 br_336 data_337 bl_337 br_337 data_338 bl_338
+ br_338 data_339 bl_339 br_339 data_340 bl_340 br_340 data_341 bl_341
+ br_341 data_342 bl_342 br_342 data_343 bl_343 br_343 data_344 bl_344
+ br_344 data_345 bl_345 br_345 data_346 bl_346 br_346 data_347 bl_347
+ br_347 data_348 bl_348 br_348 data_349 bl_349 br_349 data_350 bl_350
+ br_350 data_351 bl_351 br_351 data_352 bl_352 br_352 data_353 bl_353
+ br_353 data_354 bl_354 br_354 data_355 bl_355 br_355 data_356 bl_356
+ br_356 data_357 bl_357 br_357 data_358 bl_358 br_358 data_359 bl_359
+ br_359 data_360 bl_360 br_360 data_361 bl_361 br_361 data_362 bl_362
+ br_362 data_363 bl_363 br_363 data_364 bl_364 br_364 data_365 bl_365
+ br_365 data_366 bl_366 br_366 data_367 bl_367 br_367 data_368 bl_368
+ br_368 data_369 bl_369 br_369 data_370 bl_370 br_370 data_371 bl_371
+ br_371 data_372 bl_372 br_372 data_373 bl_373 br_373 data_374 bl_374
+ br_374 data_375 bl_375 br_375 data_376 bl_376 br_376 data_377 bl_377
+ br_377 data_378 bl_378 br_378 data_379 bl_379 br_379 data_380 bl_380
+ br_380 data_381 bl_381 br_381 data_382 bl_382 br_382 data_383 bl_383
+ br_383 data_384 bl_384 br_384 data_385 bl_385 br_385 data_386 bl_386
+ br_386 data_387 bl_387 br_387 data_388 bl_388 br_388 data_389 bl_389
+ br_389 data_390 bl_390 br_390 data_391 bl_391 br_391 data_392 bl_392
+ br_392 data_393 bl_393 br_393 data_394 bl_394 br_394 data_395 bl_395
+ br_395 data_396 bl_396 br_396 data_397 bl_397 br_397 data_398 bl_398
+ br_398 data_399 bl_399 br_399 data_400 bl_400 br_400 data_401 bl_401
+ br_401 data_402 bl_402 br_402 data_403 bl_403 br_403 data_404 bl_404
+ br_404 data_405 bl_405 br_405 data_406 bl_406 br_406 data_407 bl_407
+ br_407 data_408 bl_408 br_408 data_409 bl_409 br_409 data_410 bl_410
+ br_410 data_411 bl_411 br_411 data_412 bl_412 br_412 data_413 bl_413
+ br_413 data_414 bl_414 br_414 data_415 bl_415 br_415 data_416 bl_416
+ br_416 data_417 bl_417 br_417 data_418 bl_418 br_418 data_419 bl_419
+ br_419 data_420 bl_420 br_420 data_421 bl_421 br_421 data_422 bl_422
+ br_422 data_423 bl_423 br_423 data_424 bl_424 br_424 data_425 bl_425
+ br_425 data_426 bl_426 br_426 data_427 bl_427 br_427 data_428 bl_428
+ br_428 data_429 bl_429 br_429 data_430 bl_430 br_430 data_431 bl_431
+ br_431 data_432 bl_432 br_432 data_433 bl_433 br_433 data_434 bl_434
+ br_434 data_435 bl_435 br_435 data_436 bl_436 br_436 data_437 bl_437
+ br_437 data_438 bl_438 br_438 data_439 bl_439 br_439 data_440 bl_440
+ br_440 data_441 bl_441 br_441 data_442 bl_442 br_442 data_443 bl_443
+ br_443 data_444 bl_444 br_444 data_445 bl_445 br_445 data_446 bl_446
+ br_446 data_447 bl_447 br_447 data_448 bl_448 br_448 data_449 bl_449
+ br_449 data_450 bl_450 br_450 data_451 bl_451 br_451 data_452 bl_452
+ br_452 data_453 bl_453 br_453 data_454 bl_454 br_454 data_455 bl_455
+ br_455 data_456 bl_456 br_456 data_457 bl_457 br_457 data_458 bl_458
+ br_458 data_459 bl_459 br_459 data_460 bl_460 br_460 data_461 bl_461
+ br_461 data_462 bl_462 br_462 data_463 bl_463 br_463 data_464 bl_464
+ br_464 data_465 bl_465 br_465 data_466 bl_466 br_466 data_467 bl_467
+ br_467 data_468 bl_468 br_468 data_469 bl_469 br_469 data_470 bl_470
+ br_470 data_471 bl_471 br_471 data_472 bl_472 br_472 data_473 bl_473
+ br_473 data_474 bl_474 br_474 data_475 bl_475 br_475 data_476 bl_476
+ br_476 data_477 bl_477 br_477 data_478 bl_478 br_478 data_479 bl_479
+ br_479 data_480 bl_480 br_480 data_481 bl_481 br_481 data_482 bl_482
+ br_482 data_483 bl_483 br_483 data_484 bl_484 br_484 data_485 bl_485
+ br_485 data_486 bl_486 br_486 data_487 bl_487 br_487 data_488 bl_488
+ br_488 data_489 bl_489 br_489 data_490 bl_490 br_490 data_491 bl_491
+ br_491 data_492 bl_492 br_492 data_493 bl_493 br_493 data_494 bl_494
+ br_494 data_495 bl_495 br_495 data_496 bl_496 br_496 data_497 bl_497
+ br_497 data_498 bl_498 br_498 data_499 bl_499 br_499 data_500 bl_500
+ br_500 data_501 bl_501 br_501 data_502 bl_502 br_502 data_503 bl_503
+ br_503 data_504 bl_504 br_504 data_505 bl_505 br_505 data_506 bl_506
+ br_506 data_507 bl_507 br_507 data_508 bl_508 br_508 data_509 bl_509
+ br_509 data_510 bl_510 br_510 data_511 bl_511 br_511 en vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* OUTPUT: data_32 
* INPUT : bl_32 
* INPUT : br_32 
* OUTPUT: data_33 
* INPUT : bl_33 
* INPUT : br_33 
* OUTPUT: data_34 
* INPUT : bl_34 
* INPUT : br_34 
* OUTPUT: data_35 
* INPUT : bl_35 
* INPUT : br_35 
* OUTPUT: data_36 
* INPUT : bl_36 
* INPUT : br_36 
* OUTPUT: data_37 
* INPUT : bl_37 
* INPUT : br_37 
* OUTPUT: data_38 
* INPUT : bl_38 
* INPUT : br_38 
* OUTPUT: data_39 
* INPUT : bl_39 
* INPUT : br_39 
* OUTPUT: data_40 
* INPUT : bl_40 
* INPUT : br_40 
* OUTPUT: data_41 
* INPUT : bl_41 
* INPUT : br_41 
* OUTPUT: data_42 
* INPUT : bl_42 
* INPUT : br_42 
* OUTPUT: data_43 
* INPUT : bl_43 
* INPUT : br_43 
* OUTPUT: data_44 
* INPUT : bl_44 
* INPUT : br_44 
* OUTPUT: data_45 
* INPUT : bl_45 
* INPUT : br_45 
* OUTPUT: data_46 
* INPUT : bl_46 
* INPUT : br_46 
* OUTPUT: data_47 
* INPUT : bl_47 
* INPUT : br_47 
* OUTPUT: data_48 
* INPUT : bl_48 
* INPUT : br_48 
* OUTPUT: data_49 
* INPUT : bl_49 
* INPUT : br_49 
* OUTPUT: data_50 
* INPUT : bl_50 
* INPUT : br_50 
* OUTPUT: data_51 
* INPUT : bl_51 
* INPUT : br_51 
* OUTPUT: data_52 
* INPUT : bl_52 
* INPUT : br_52 
* OUTPUT: data_53 
* INPUT : bl_53 
* INPUT : br_53 
* OUTPUT: data_54 
* INPUT : bl_54 
* INPUT : br_54 
* OUTPUT: data_55 
* INPUT : bl_55 
* INPUT : br_55 
* OUTPUT: data_56 
* INPUT : bl_56 
* INPUT : br_56 
* OUTPUT: data_57 
* INPUT : bl_57 
* INPUT : br_57 
* OUTPUT: data_58 
* INPUT : bl_58 
* INPUT : br_58 
* OUTPUT: data_59 
* INPUT : bl_59 
* INPUT : br_59 
* OUTPUT: data_60 
* INPUT : bl_60 
* INPUT : br_60 
* OUTPUT: data_61 
* INPUT : bl_61 
* INPUT : br_61 
* OUTPUT: data_62 
* INPUT : bl_62 
* INPUT : br_62 
* OUTPUT: data_63 
* INPUT : bl_63 
* INPUT : br_63 
* OUTPUT: data_64 
* INPUT : bl_64 
* INPUT : br_64 
* OUTPUT: data_65 
* INPUT : bl_65 
* INPUT : br_65 
* OUTPUT: data_66 
* INPUT : bl_66 
* INPUT : br_66 
* OUTPUT: data_67 
* INPUT : bl_67 
* INPUT : br_67 
* OUTPUT: data_68 
* INPUT : bl_68 
* INPUT : br_68 
* OUTPUT: data_69 
* INPUT : bl_69 
* INPUT : br_69 
* OUTPUT: data_70 
* INPUT : bl_70 
* INPUT : br_70 
* OUTPUT: data_71 
* INPUT : bl_71 
* INPUT : br_71 
* OUTPUT: data_72 
* INPUT : bl_72 
* INPUT : br_72 
* OUTPUT: data_73 
* INPUT : bl_73 
* INPUT : br_73 
* OUTPUT: data_74 
* INPUT : bl_74 
* INPUT : br_74 
* OUTPUT: data_75 
* INPUT : bl_75 
* INPUT : br_75 
* OUTPUT: data_76 
* INPUT : bl_76 
* INPUT : br_76 
* OUTPUT: data_77 
* INPUT : bl_77 
* INPUT : br_77 
* OUTPUT: data_78 
* INPUT : bl_78 
* INPUT : br_78 
* OUTPUT: data_79 
* INPUT : bl_79 
* INPUT : br_79 
* OUTPUT: data_80 
* INPUT : bl_80 
* INPUT : br_80 
* OUTPUT: data_81 
* INPUT : bl_81 
* INPUT : br_81 
* OUTPUT: data_82 
* INPUT : bl_82 
* INPUT : br_82 
* OUTPUT: data_83 
* INPUT : bl_83 
* INPUT : br_83 
* OUTPUT: data_84 
* INPUT : bl_84 
* INPUT : br_84 
* OUTPUT: data_85 
* INPUT : bl_85 
* INPUT : br_85 
* OUTPUT: data_86 
* INPUT : bl_86 
* INPUT : br_86 
* OUTPUT: data_87 
* INPUT : bl_87 
* INPUT : br_87 
* OUTPUT: data_88 
* INPUT : bl_88 
* INPUT : br_88 
* OUTPUT: data_89 
* INPUT : bl_89 
* INPUT : br_89 
* OUTPUT: data_90 
* INPUT : bl_90 
* INPUT : br_90 
* OUTPUT: data_91 
* INPUT : bl_91 
* INPUT : br_91 
* OUTPUT: data_92 
* INPUT : bl_92 
* INPUT : br_92 
* OUTPUT: data_93 
* INPUT : bl_93 
* INPUT : br_93 
* OUTPUT: data_94 
* INPUT : bl_94 
* INPUT : br_94 
* OUTPUT: data_95 
* INPUT : bl_95 
* INPUT : br_95 
* OUTPUT: data_96 
* INPUT : bl_96 
* INPUT : br_96 
* OUTPUT: data_97 
* INPUT : bl_97 
* INPUT : br_97 
* OUTPUT: data_98 
* INPUT : bl_98 
* INPUT : br_98 
* OUTPUT: data_99 
* INPUT : bl_99 
* INPUT : br_99 
* OUTPUT: data_100 
* INPUT : bl_100 
* INPUT : br_100 
* OUTPUT: data_101 
* INPUT : bl_101 
* INPUT : br_101 
* OUTPUT: data_102 
* INPUT : bl_102 
* INPUT : br_102 
* OUTPUT: data_103 
* INPUT : bl_103 
* INPUT : br_103 
* OUTPUT: data_104 
* INPUT : bl_104 
* INPUT : br_104 
* OUTPUT: data_105 
* INPUT : bl_105 
* INPUT : br_105 
* OUTPUT: data_106 
* INPUT : bl_106 
* INPUT : br_106 
* OUTPUT: data_107 
* INPUT : bl_107 
* INPUT : br_107 
* OUTPUT: data_108 
* INPUT : bl_108 
* INPUT : br_108 
* OUTPUT: data_109 
* INPUT : bl_109 
* INPUT : br_109 
* OUTPUT: data_110 
* INPUT : bl_110 
* INPUT : br_110 
* OUTPUT: data_111 
* INPUT : bl_111 
* INPUT : br_111 
* OUTPUT: data_112 
* INPUT : bl_112 
* INPUT : br_112 
* OUTPUT: data_113 
* INPUT : bl_113 
* INPUT : br_113 
* OUTPUT: data_114 
* INPUT : bl_114 
* INPUT : br_114 
* OUTPUT: data_115 
* INPUT : bl_115 
* INPUT : br_115 
* OUTPUT: data_116 
* INPUT : bl_116 
* INPUT : br_116 
* OUTPUT: data_117 
* INPUT : bl_117 
* INPUT : br_117 
* OUTPUT: data_118 
* INPUT : bl_118 
* INPUT : br_118 
* OUTPUT: data_119 
* INPUT : bl_119 
* INPUT : br_119 
* OUTPUT: data_120 
* INPUT : bl_120 
* INPUT : br_120 
* OUTPUT: data_121 
* INPUT : bl_121 
* INPUT : br_121 
* OUTPUT: data_122 
* INPUT : bl_122 
* INPUT : br_122 
* OUTPUT: data_123 
* INPUT : bl_123 
* INPUT : br_123 
* OUTPUT: data_124 
* INPUT : bl_124 
* INPUT : br_124 
* OUTPUT: data_125 
* INPUT : bl_125 
* INPUT : br_125 
* OUTPUT: data_126 
* INPUT : bl_126 
* INPUT : br_126 
* OUTPUT: data_127 
* INPUT : bl_127 
* INPUT : br_127 
* OUTPUT: data_128 
* INPUT : bl_128 
* INPUT : br_128 
* OUTPUT: data_129 
* INPUT : bl_129 
* INPUT : br_129 
* OUTPUT: data_130 
* INPUT : bl_130 
* INPUT : br_130 
* OUTPUT: data_131 
* INPUT : bl_131 
* INPUT : br_131 
* OUTPUT: data_132 
* INPUT : bl_132 
* INPUT : br_132 
* OUTPUT: data_133 
* INPUT : bl_133 
* INPUT : br_133 
* OUTPUT: data_134 
* INPUT : bl_134 
* INPUT : br_134 
* OUTPUT: data_135 
* INPUT : bl_135 
* INPUT : br_135 
* OUTPUT: data_136 
* INPUT : bl_136 
* INPUT : br_136 
* OUTPUT: data_137 
* INPUT : bl_137 
* INPUT : br_137 
* OUTPUT: data_138 
* INPUT : bl_138 
* INPUT : br_138 
* OUTPUT: data_139 
* INPUT : bl_139 
* INPUT : br_139 
* OUTPUT: data_140 
* INPUT : bl_140 
* INPUT : br_140 
* OUTPUT: data_141 
* INPUT : bl_141 
* INPUT : br_141 
* OUTPUT: data_142 
* INPUT : bl_142 
* INPUT : br_142 
* OUTPUT: data_143 
* INPUT : bl_143 
* INPUT : br_143 
* OUTPUT: data_144 
* INPUT : bl_144 
* INPUT : br_144 
* OUTPUT: data_145 
* INPUT : bl_145 
* INPUT : br_145 
* OUTPUT: data_146 
* INPUT : bl_146 
* INPUT : br_146 
* OUTPUT: data_147 
* INPUT : bl_147 
* INPUT : br_147 
* OUTPUT: data_148 
* INPUT : bl_148 
* INPUT : br_148 
* OUTPUT: data_149 
* INPUT : bl_149 
* INPUT : br_149 
* OUTPUT: data_150 
* INPUT : bl_150 
* INPUT : br_150 
* OUTPUT: data_151 
* INPUT : bl_151 
* INPUT : br_151 
* OUTPUT: data_152 
* INPUT : bl_152 
* INPUT : br_152 
* OUTPUT: data_153 
* INPUT : bl_153 
* INPUT : br_153 
* OUTPUT: data_154 
* INPUT : bl_154 
* INPUT : br_154 
* OUTPUT: data_155 
* INPUT : bl_155 
* INPUT : br_155 
* OUTPUT: data_156 
* INPUT : bl_156 
* INPUT : br_156 
* OUTPUT: data_157 
* INPUT : bl_157 
* INPUT : br_157 
* OUTPUT: data_158 
* INPUT : bl_158 
* INPUT : br_158 
* OUTPUT: data_159 
* INPUT : bl_159 
* INPUT : br_159 
* OUTPUT: data_160 
* INPUT : bl_160 
* INPUT : br_160 
* OUTPUT: data_161 
* INPUT : bl_161 
* INPUT : br_161 
* OUTPUT: data_162 
* INPUT : bl_162 
* INPUT : br_162 
* OUTPUT: data_163 
* INPUT : bl_163 
* INPUT : br_163 
* OUTPUT: data_164 
* INPUT : bl_164 
* INPUT : br_164 
* OUTPUT: data_165 
* INPUT : bl_165 
* INPUT : br_165 
* OUTPUT: data_166 
* INPUT : bl_166 
* INPUT : br_166 
* OUTPUT: data_167 
* INPUT : bl_167 
* INPUT : br_167 
* OUTPUT: data_168 
* INPUT : bl_168 
* INPUT : br_168 
* OUTPUT: data_169 
* INPUT : bl_169 
* INPUT : br_169 
* OUTPUT: data_170 
* INPUT : bl_170 
* INPUT : br_170 
* OUTPUT: data_171 
* INPUT : bl_171 
* INPUT : br_171 
* OUTPUT: data_172 
* INPUT : bl_172 
* INPUT : br_172 
* OUTPUT: data_173 
* INPUT : bl_173 
* INPUT : br_173 
* OUTPUT: data_174 
* INPUT : bl_174 
* INPUT : br_174 
* OUTPUT: data_175 
* INPUT : bl_175 
* INPUT : br_175 
* OUTPUT: data_176 
* INPUT : bl_176 
* INPUT : br_176 
* OUTPUT: data_177 
* INPUT : bl_177 
* INPUT : br_177 
* OUTPUT: data_178 
* INPUT : bl_178 
* INPUT : br_178 
* OUTPUT: data_179 
* INPUT : bl_179 
* INPUT : br_179 
* OUTPUT: data_180 
* INPUT : bl_180 
* INPUT : br_180 
* OUTPUT: data_181 
* INPUT : bl_181 
* INPUT : br_181 
* OUTPUT: data_182 
* INPUT : bl_182 
* INPUT : br_182 
* OUTPUT: data_183 
* INPUT : bl_183 
* INPUT : br_183 
* OUTPUT: data_184 
* INPUT : bl_184 
* INPUT : br_184 
* OUTPUT: data_185 
* INPUT : bl_185 
* INPUT : br_185 
* OUTPUT: data_186 
* INPUT : bl_186 
* INPUT : br_186 
* OUTPUT: data_187 
* INPUT : bl_187 
* INPUT : br_187 
* OUTPUT: data_188 
* INPUT : bl_188 
* INPUT : br_188 
* OUTPUT: data_189 
* INPUT : bl_189 
* INPUT : br_189 
* OUTPUT: data_190 
* INPUT : bl_190 
* INPUT : br_190 
* OUTPUT: data_191 
* INPUT : bl_191 
* INPUT : br_191 
* OUTPUT: data_192 
* INPUT : bl_192 
* INPUT : br_192 
* OUTPUT: data_193 
* INPUT : bl_193 
* INPUT : br_193 
* OUTPUT: data_194 
* INPUT : bl_194 
* INPUT : br_194 
* OUTPUT: data_195 
* INPUT : bl_195 
* INPUT : br_195 
* OUTPUT: data_196 
* INPUT : bl_196 
* INPUT : br_196 
* OUTPUT: data_197 
* INPUT : bl_197 
* INPUT : br_197 
* OUTPUT: data_198 
* INPUT : bl_198 
* INPUT : br_198 
* OUTPUT: data_199 
* INPUT : bl_199 
* INPUT : br_199 
* OUTPUT: data_200 
* INPUT : bl_200 
* INPUT : br_200 
* OUTPUT: data_201 
* INPUT : bl_201 
* INPUT : br_201 
* OUTPUT: data_202 
* INPUT : bl_202 
* INPUT : br_202 
* OUTPUT: data_203 
* INPUT : bl_203 
* INPUT : br_203 
* OUTPUT: data_204 
* INPUT : bl_204 
* INPUT : br_204 
* OUTPUT: data_205 
* INPUT : bl_205 
* INPUT : br_205 
* OUTPUT: data_206 
* INPUT : bl_206 
* INPUT : br_206 
* OUTPUT: data_207 
* INPUT : bl_207 
* INPUT : br_207 
* OUTPUT: data_208 
* INPUT : bl_208 
* INPUT : br_208 
* OUTPUT: data_209 
* INPUT : bl_209 
* INPUT : br_209 
* OUTPUT: data_210 
* INPUT : bl_210 
* INPUT : br_210 
* OUTPUT: data_211 
* INPUT : bl_211 
* INPUT : br_211 
* OUTPUT: data_212 
* INPUT : bl_212 
* INPUT : br_212 
* OUTPUT: data_213 
* INPUT : bl_213 
* INPUT : br_213 
* OUTPUT: data_214 
* INPUT : bl_214 
* INPUT : br_214 
* OUTPUT: data_215 
* INPUT : bl_215 
* INPUT : br_215 
* OUTPUT: data_216 
* INPUT : bl_216 
* INPUT : br_216 
* OUTPUT: data_217 
* INPUT : bl_217 
* INPUT : br_217 
* OUTPUT: data_218 
* INPUT : bl_218 
* INPUT : br_218 
* OUTPUT: data_219 
* INPUT : bl_219 
* INPUT : br_219 
* OUTPUT: data_220 
* INPUT : bl_220 
* INPUT : br_220 
* OUTPUT: data_221 
* INPUT : bl_221 
* INPUT : br_221 
* OUTPUT: data_222 
* INPUT : bl_222 
* INPUT : br_222 
* OUTPUT: data_223 
* INPUT : bl_223 
* INPUT : br_223 
* OUTPUT: data_224 
* INPUT : bl_224 
* INPUT : br_224 
* OUTPUT: data_225 
* INPUT : bl_225 
* INPUT : br_225 
* OUTPUT: data_226 
* INPUT : bl_226 
* INPUT : br_226 
* OUTPUT: data_227 
* INPUT : bl_227 
* INPUT : br_227 
* OUTPUT: data_228 
* INPUT : bl_228 
* INPUT : br_228 
* OUTPUT: data_229 
* INPUT : bl_229 
* INPUT : br_229 
* OUTPUT: data_230 
* INPUT : bl_230 
* INPUT : br_230 
* OUTPUT: data_231 
* INPUT : bl_231 
* INPUT : br_231 
* OUTPUT: data_232 
* INPUT : bl_232 
* INPUT : br_232 
* OUTPUT: data_233 
* INPUT : bl_233 
* INPUT : br_233 
* OUTPUT: data_234 
* INPUT : bl_234 
* INPUT : br_234 
* OUTPUT: data_235 
* INPUT : bl_235 
* INPUT : br_235 
* OUTPUT: data_236 
* INPUT : bl_236 
* INPUT : br_236 
* OUTPUT: data_237 
* INPUT : bl_237 
* INPUT : br_237 
* OUTPUT: data_238 
* INPUT : bl_238 
* INPUT : br_238 
* OUTPUT: data_239 
* INPUT : bl_239 
* INPUT : br_239 
* OUTPUT: data_240 
* INPUT : bl_240 
* INPUT : br_240 
* OUTPUT: data_241 
* INPUT : bl_241 
* INPUT : br_241 
* OUTPUT: data_242 
* INPUT : bl_242 
* INPUT : br_242 
* OUTPUT: data_243 
* INPUT : bl_243 
* INPUT : br_243 
* OUTPUT: data_244 
* INPUT : bl_244 
* INPUT : br_244 
* OUTPUT: data_245 
* INPUT : bl_245 
* INPUT : br_245 
* OUTPUT: data_246 
* INPUT : bl_246 
* INPUT : br_246 
* OUTPUT: data_247 
* INPUT : bl_247 
* INPUT : br_247 
* OUTPUT: data_248 
* INPUT : bl_248 
* INPUT : br_248 
* OUTPUT: data_249 
* INPUT : bl_249 
* INPUT : br_249 
* OUTPUT: data_250 
* INPUT : bl_250 
* INPUT : br_250 
* OUTPUT: data_251 
* INPUT : bl_251 
* INPUT : br_251 
* OUTPUT: data_252 
* INPUT : bl_252 
* INPUT : br_252 
* OUTPUT: data_253 
* INPUT : bl_253 
* INPUT : br_253 
* OUTPUT: data_254 
* INPUT : bl_254 
* INPUT : br_254 
* OUTPUT: data_255 
* INPUT : bl_255 
* INPUT : br_255 
* OUTPUT: data_256 
* INPUT : bl_256 
* INPUT : br_256 
* OUTPUT: data_257 
* INPUT : bl_257 
* INPUT : br_257 
* OUTPUT: data_258 
* INPUT : bl_258 
* INPUT : br_258 
* OUTPUT: data_259 
* INPUT : bl_259 
* INPUT : br_259 
* OUTPUT: data_260 
* INPUT : bl_260 
* INPUT : br_260 
* OUTPUT: data_261 
* INPUT : bl_261 
* INPUT : br_261 
* OUTPUT: data_262 
* INPUT : bl_262 
* INPUT : br_262 
* OUTPUT: data_263 
* INPUT : bl_263 
* INPUT : br_263 
* OUTPUT: data_264 
* INPUT : bl_264 
* INPUT : br_264 
* OUTPUT: data_265 
* INPUT : bl_265 
* INPUT : br_265 
* OUTPUT: data_266 
* INPUT : bl_266 
* INPUT : br_266 
* OUTPUT: data_267 
* INPUT : bl_267 
* INPUT : br_267 
* OUTPUT: data_268 
* INPUT : bl_268 
* INPUT : br_268 
* OUTPUT: data_269 
* INPUT : bl_269 
* INPUT : br_269 
* OUTPUT: data_270 
* INPUT : bl_270 
* INPUT : br_270 
* OUTPUT: data_271 
* INPUT : bl_271 
* INPUT : br_271 
* OUTPUT: data_272 
* INPUT : bl_272 
* INPUT : br_272 
* OUTPUT: data_273 
* INPUT : bl_273 
* INPUT : br_273 
* OUTPUT: data_274 
* INPUT : bl_274 
* INPUT : br_274 
* OUTPUT: data_275 
* INPUT : bl_275 
* INPUT : br_275 
* OUTPUT: data_276 
* INPUT : bl_276 
* INPUT : br_276 
* OUTPUT: data_277 
* INPUT : bl_277 
* INPUT : br_277 
* OUTPUT: data_278 
* INPUT : bl_278 
* INPUT : br_278 
* OUTPUT: data_279 
* INPUT : bl_279 
* INPUT : br_279 
* OUTPUT: data_280 
* INPUT : bl_280 
* INPUT : br_280 
* OUTPUT: data_281 
* INPUT : bl_281 
* INPUT : br_281 
* OUTPUT: data_282 
* INPUT : bl_282 
* INPUT : br_282 
* OUTPUT: data_283 
* INPUT : bl_283 
* INPUT : br_283 
* OUTPUT: data_284 
* INPUT : bl_284 
* INPUT : br_284 
* OUTPUT: data_285 
* INPUT : bl_285 
* INPUT : br_285 
* OUTPUT: data_286 
* INPUT : bl_286 
* INPUT : br_286 
* OUTPUT: data_287 
* INPUT : bl_287 
* INPUT : br_287 
* OUTPUT: data_288 
* INPUT : bl_288 
* INPUT : br_288 
* OUTPUT: data_289 
* INPUT : bl_289 
* INPUT : br_289 
* OUTPUT: data_290 
* INPUT : bl_290 
* INPUT : br_290 
* OUTPUT: data_291 
* INPUT : bl_291 
* INPUT : br_291 
* OUTPUT: data_292 
* INPUT : bl_292 
* INPUT : br_292 
* OUTPUT: data_293 
* INPUT : bl_293 
* INPUT : br_293 
* OUTPUT: data_294 
* INPUT : bl_294 
* INPUT : br_294 
* OUTPUT: data_295 
* INPUT : bl_295 
* INPUT : br_295 
* OUTPUT: data_296 
* INPUT : bl_296 
* INPUT : br_296 
* OUTPUT: data_297 
* INPUT : bl_297 
* INPUT : br_297 
* OUTPUT: data_298 
* INPUT : bl_298 
* INPUT : br_298 
* OUTPUT: data_299 
* INPUT : bl_299 
* INPUT : br_299 
* OUTPUT: data_300 
* INPUT : bl_300 
* INPUT : br_300 
* OUTPUT: data_301 
* INPUT : bl_301 
* INPUT : br_301 
* OUTPUT: data_302 
* INPUT : bl_302 
* INPUT : br_302 
* OUTPUT: data_303 
* INPUT : bl_303 
* INPUT : br_303 
* OUTPUT: data_304 
* INPUT : bl_304 
* INPUT : br_304 
* OUTPUT: data_305 
* INPUT : bl_305 
* INPUT : br_305 
* OUTPUT: data_306 
* INPUT : bl_306 
* INPUT : br_306 
* OUTPUT: data_307 
* INPUT : bl_307 
* INPUT : br_307 
* OUTPUT: data_308 
* INPUT : bl_308 
* INPUT : br_308 
* OUTPUT: data_309 
* INPUT : bl_309 
* INPUT : br_309 
* OUTPUT: data_310 
* INPUT : bl_310 
* INPUT : br_310 
* OUTPUT: data_311 
* INPUT : bl_311 
* INPUT : br_311 
* OUTPUT: data_312 
* INPUT : bl_312 
* INPUT : br_312 
* OUTPUT: data_313 
* INPUT : bl_313 
* INPUT : br_313 
* OUTPUT: data_314 
* INPUT : bl_314 
* INPUT : br_314 
* OUTPUT: data_315 
* INPUT : bl_315 
* INPUT : br_315 
* OUTPUT: data_316 
* INPUT : bl_316 
* INPUT : br_316 
* OUTPUT: data_317 
* INPUT : bl_317 
* INPUT : br_317 
* OUTPUT: data_318 
* INPUT : bl_318 
* INPUT : br_318 
* OUTPUT: data_319 
* INPUT : bl_319 
* INPUT : br_319 
* OUTPUT: data_320 
* INPUT : bl_320 
* INPUT : br_320 
* OUTPUT: data_321 
* INPUT : bl_321 
* INPUT : br_321 
* OUTPUT: data_322 
* INPUT : bl_322 
* INPUT : br_322 
* OUTPUT: data_323 
* INPUT : bl_323 
* INPUT : br_323 
* OUTPUT: data_324 
* INPUT : bl_324 
* INPUT : br_324 
* OUTPUT: data_325 
* INPUT : bl_325 
* INPUT : br_325 
* OUTPUT: data_326 
* INPUT : bl_326 
* INPUT : br_326 
* OUTPUT: data_327 
* INPUT : bl_327 
* INPUT : br_327 
* OUTPUT: data_328 
* INPUT : bl_328 
* INPUT : br_328 
* OUTPUT: data_329 
* INPUT : bl_329 
* INPUT : br_329 
* OUTPUT: data_330 
* INPUT : bl_330 
* INPUT : br_330 
* OUTPUT: data_331 
* INPUT : bl_331 
* INPUT : br_331 
* OUTPUT: data_332 
* INPUT : bl_332 
* INPUT : br_332 
* OUTPUT: data_333 
* INPUT : bl_333 
* INPUT : br_333 
* OUTPUT: data_334 
* INPUT : bl_334 
* INPUT : br_334 
* OUTPUT: data_335 
* INPUT : bl_335 
* INPUT : br_335 
* OUTPUT: data_336 
* INPUT : bl_336 
* INPUT : br_336 
* OUTPUT: data_337 
* INPUT : bl_337 
* INPUT : br_337 
* OUTPUT: data_338 
* INPUT : bl_338 
* INPUT : br_338 
* OUTPUT: data_339 
* INPUT : bl_339 
* INPUT : br_339 
* OUTPUT: data_340 
* INPUT : bl_340 
* INPUT : br_340 
* OUTPUT: data_341 
* INPUT : bl_341 
* INPUT : br_341 
* OUTPUT: data_342 
* INPUT : bl_342 
* INPUT : br_342 
* OUTPUT: data_343 
* INPUT : bl_343 
* INPUT : br_343 
* OUTPUT: data_344 
* INPUT : bl_344 
* INPUT : br_344 
* OUTPUT: data_345 
* INPUT : bl_345 
* INPUT : br_345 
* OUTPUT: data_346 
* INPUT : bl_346 
* INPUT : br_346 
* OUTPUT: data_347 
* INPUT : bl_347 
* INPUT : br_347 
* OUTPUT: data_348 
* INPUT : bl_348 
* INPUT : br_348 
* OUTPUT: data_349 
* INPUT : bl_349 
* INPUT : br_349 
* OUTPUT: data_350 
* INPUT : bl_350 
* INPUT : br_350 
* OUTPUT: data_351 
* INPUT : bl_351 
* INPUT : br_351 
* OUTPUT: data_352 
* INPUT : bl_352 
* INPUT : br_352 
* OUTPUT: data_353 
* INPUT : bl_353 
* INPUT : br_353 
* OUTPUT: data_354 
* INPUT : bl_354 
* INPUT : br_354 
* OUTPUT: data_355 
* INPUT : bl_355 
* INPUT : br_355 
* OUTPUT: data_356 
* INPUT : bl_356 
* INPUT : br_356 
* OUTPUT: data_357 
* INPUT : bl_357 
* INPUT : br_357 
* OUTPUT: data_358 
* INPUT : bl_358 
* INPUT : br_358 
* OUTPUT: data_359 
* INPUT : bl_359 
* INPUT : br_359 
* OUTPUT: data_360 
* INPUT : bl_360 
* INPUT : br_360 
* OUTPUT: data_361 
* INPUT : bl_361 
* INPUT : br_361 
* OUTPUT: data_362 
* INPUT : bl_362 
* INPUT : br_362 
* OUTPUT: data_363 
* INPUT : bl_363 
* INPUT : br_363 
* OUTPUT: data_364 
* INPUT : bl_364 
* INPUT : br_364 
* OUTPUT: data_365 
* INPUT : bl_365 
* INPUT : br_365 
* OUTPUT: data_366 
* INPUT : bl_366 
* INPUT : br_366 
* OUTPUT: data_367 
* INPUT : bl_367 
* INPUT : br_367 
* OUTPUT: data_368 
* INPUT : bl_368 
* INPUT : br_368 
* OUTPUT: data_369 
* INPUT : bl_369 
* INPUT : br_369 
* OUTPUT: data_370 
* INPUT : bl_370 
* INPUT : br_370 
* OUTPUT: data_371 
* INPUT : bl_371 
* INPUT : br_371 
* OUTPUT: data_372 
* INPUT : bl_372 
* INPUT : br_372 
* OUTPUT: data_373 
* INPUT : bl_373 
* INPUT : br_373 
* OUTPUT: data_374 
* INPUT : bl_374 
* INPUT : br_374 
* OUTPUT: data_375 
* INPUT : bl_375 
* INPUT : br_375 
* OUTPUT: data_376 
* INPUT : bl_376 
* INPUT : br_376 
* OUTPUT: data_377 
* INPUT : bl_377 
* INPUT : br_377 
* OUTPUT: data_378 
* INPUT : bl_378 
* INPUT : br_378 
* OUTPUT: data_379 
* INPUT : bl_379 
* INPUT : br_379 
* OUTPUT: data_380 
* INPUT : bl_380 
* INPUT : br_380 
* OUTPUT: data_381 
* INPUT : bl_381 
* INPUT : br_381 
* OUTPUT: data_382 
* INPUT : bl_382 
* INPUT : br_382 
* OUTPUT: data_383 
* INPUT : bl_383 
* INPUT : br_383 
* OUTPUT: data_384 
* INPUT : bl_384 
* INPUT : br_384 
* OUTPUT: data_385 
* INPUT : bl_385 
* INPUT : br_385 
* OUTPUT: data_386 
* INPUT : bl_386 
* INPUT : br_386 
* OUTPUT: data_387 
* INPUT : bl_387 
* INPUT : br_387 
* OUTPUT: data_388 
* INPUT : bl_388 
* INPUT : br_388 
* OUTPUT: data_389 
* INPUT : bl_389 
* INPUT : br_389 
* OUTPUT: data_390 
* INPUT : bl_390 
* INPUT : br_390 
* OUTPUT: data_391 
* INPUT : bl_391 
* INPUT : br_391 
* OUTPUT: data_392 
* INPUT : bl_392 
* INPUT : br_392 
* OUTPUT: data_393 
* INPUT : bl_393 
* INPUT : br_393 
* OUTPUT: data_394 
* INPUT : bl_394 
* INPUT : br_394 
* OUTPUT: data_395 
* INPUT : bl_395 
* INPUT : br_395 
* OUTPUT: data_396 
* INPUT : bl_396 
* INPUT : br_396 
* OUTPUT: data_397 
* INPUT : bl_397 
* INPUT : br_397 
* OUTPUT: data_398 
* INPUT : bl_398 
* INPUT : br_398 
* OUTPUT: data_399 
* INPUT : bl_399 
* INPUT : br_399 
* OUTPUT: data_400 
* INPUT : bl_400 
* INPUT : br_400 
* OUTPUT: data_401 
* INPUT : bl_401 
* INPUT : br_401 
* OUTPUT: data_402 
* INPUT : bl_402 
* INPUT : br_402 
* OUTPUT: data_403 
* INPUT : bl_403 
* INPUT : br_403 
* OUTPUT: data_404 
* INPUT : bl_404 
* INPUT : br_404 
* OUTPUT: data_405 
* INPUT : bl_405 
* INPUT : br_405 
* OUTPUT: data_406 
* INPUT : bl_406 
* INPUT : br_406 
* OUTPUT: data_407 
* INPUT : bl_407 
* INPUT : br_407 
* OUTPUT: data_408 
* INPUT : bl_408 
* INPUT : br_408 
* OUTPUT: data_409 
* INPUT : bl_409 
* INPUT : br_409 
* OUTPUT: data_410 
* INPUT : bl_410 
* INPUT : br_410 
* OUTPUT: data_411 
* INPUT : bl_411 
* INPUT : br_411 
* OUTPUT: data_412 
* INPUT : bl_412 
* INPUT : br_412 
* OUTPUT: data_413 
* INPUT : bl_413 
* INPUT : br_413 
* OUTPUT: data_414 
* INPUT : bl_414 
* INPUT : br_414 
* OUTPUT: data_415 
* INPUT : bl_415 
* INPUT : br_415 
* OUTPUT: data_416 
* INPUT : bl_416 
* INPUT : br_416 
* OUTPUT: data_417 
* INPUT : bl_417 
* INPUT : br_417 
* OUTPUT: data_418 
* INPUT : bl_418 
* INPUT : br_418 
* OUTPUT: data_419 
* INPUT : bl_419 
* INPUT : br_419 
* OUTPUT: data_420 
* INPUT : bl_420 
* INPUT : br_420 
* OUTPUT: data_421 
* INPUT : bl_421 
* INPUT : br_421 
* OUTPUT: data_422 
* INPUT : bl_422 
* INPUT : br_422 
* OUTPUT: data_423 
* INPUT : bl_423 
* INPUT : br_423 
* OUTPUT: data_424 
* INPUT : bl_424 
* INPUT : br_424 
* OUTPUT: data_425 
* INPUT : bl_425 
* INPUT : br_425 
* OUTPUT: data_426 
* INPUT : bl_426 
* INPUT : br_426 
* OUTPUT: data_427 
* INPUT : bl_427 
* INPUT : br_427 
* OUTPUT: data_428 
* INPUT : bl_428 
* INPUT : br_428 
* OUTPUT: data_429 
* INPUT : bl_429 
* INPUT : br_429 
* OUTPUT: data_430 
* INPUT : bl_430 
* INPUT : br_430 
* OUTPUT: data_431 
* INPUT : bl_431 
* INPUT : br_431 
* OUTPUT: data_432 
* INPUT : bl_432 
* INPUT : br_432 
* OUTPUT: data_433 
* INPUT : bl_433 
* INPUT : br_433 
* OUTPUT: data_434 
* INPUT : bl_434 
* INPUT : br_434 
* OUTPUT: data_435 
* INPUT : bl_435 
* INPUT : br_435 
* OUTPUT: data_436 
* INPUT : bl_436 
* INPUT : br_436 
* OUTPUT: data_437 
* INPUT : bl_437 
* INPUT : br_437 
* OUTPUT: data_438 
* INPUT : bl_438 
* INPUT : br_438 
* OUTPUT: data_439 
* INPUT : bl_439 
* INPUT : br_439 
* OUTPUT: data_440 
* INPUT : bl_440 
* INPUT : br_440 
* OUTPUT: data_441 
* INPUT : bl_441 
* INPUT : br_441 
* OUTPUT: data_442 
* INPUT : bl_442 
* INPUT : br_442 
* OUTPUT: data_443 
* INPUT : bl_443 
* INPUT : br_443 
* OUTPUT: data_444 
* INPUT : bl_444 
* INPUT : br_444 
* OUTPUT: data_445 
* INPUT : bl_445 
* INPUT : br_445 
* OUTPUT: data_446 
* INPUT : bl_446 
* INPUT : br_446 
* OUTPUT: data_447 
* INPUT : bl_447 
* INPUT : br_447 
* OUTPUT: data_448 
* INPUT : bl_448 
* INPUT : br_448 
* OUTPUT: data_449 
* INPUT : bl_449 
* INPUT : br_449 
* OUTPUT: data_450 
* INPUT : bl_450 
* INPUT : br_450 
* OUTPUT: data_451 
* INPUT : bl_451 
* INPUT : br_451 
* OUTPUT: data_452 
* INPUT : bl_452 
* INPUT : br_452 
* OUTPUT: data_453 
* INPUT : bl_453 
* INPUT : br_453 
* OUTPUT: data_454 
* INPUT : bl_454 
* INPUT : br_454 
* OUTPUT: data_455 
* INPUT : bl_455 
* INPUT : br_455 
* OUTPUT: data_456 
* INPUT : bl_456 
* INPUT : br_456 
* OUTPUT: data_457 
* INPUT : bl_457 
* INPUT : br_457 
* OUTPUT: data_458 
* INPUT : bl_458 
* INPUT : br_458 
* OUTPUT: data_459 
* INPUT : bl_459 
* INPUT : br_459 
* OUTPUT: data_460 
* INPUT : bl_460 
* INPUT : br_460 
* OUTPUT: data_461 
* INPUT : bl_461 
* INPUT : br_461 
* OUTPUT: data_462 
* INPUT : bl_462 
* INPUT : br_462 
* OUTPUT: data_463 
* INPUT : bl_463 
* INPUT : br_463 
* OUTPUT: data_464 
* INPUT : bl_464 
* INPUT : br_464 
* OUTPUT: data_465 
* INPUT : bl_465 
* INPUT : br_465 
* OUTPUT: data_466 
* INPUT : bl_466 
* INPUT : br_466 
* OUTPUT: data_467 
* INPUT : bl_467 
* INPUT : br_467 
* OUTPUT: data_468 
* INPUT : bl_468 
* INPUT : br_468 
* OUTPUT: data_469 
* INPUT : bl_469 
* INPUT : br_469 
* OUTPUT: data_470 
* INPUT : bl_470 
* INPUT : br_470 
* OUTPUT: data_471 
* INPUT : bl_471 
* INPUT : br_471 
* OUTPUT: data_472 
* INPUT : bl_472 
* INPUT : br_472 
* OUTPUT: data_473 
* INPUT : bl_473 
* INPUT : br_473 
* OUTPUT: data_474 
* INPUT : bl_474 
* INPUT : br_474 
* OUTPUT: data_475 
* INPUT : bl_475 
* INPUT : br_475 
* OUTPUT: data_476 
* INPUT : bl_476 
* INPUT : br_476 
* OUTPUT: data_477 
* INPUT : bl_477 
* INPUT : br_477 
* OUTPUT: data_478 
* INPUT : bl_478 
* INPUT : br_478 
* OUTPUT: data_479 
* INPUT : bl_479 
* INPUT : br_479 
* OUTPUT: data_480 
* INPUT : bl_480 
* INPUT : br_480 
* OUTPUT: data_481 
* INPUT : bl_481 
* INPUT : br_481 
* OUTPUT: data_482 
* INPUT : bl_482 
* INPUT : br_482 
* OUTPUT: data_483 
* INPUT : bl_483 
* INPUT : br_483 
* OUTPUT: data_484 
* INPUT : bl_484 
* INPUT : br_484 
* OUTPUT: data_485 
* INPUT : bl_485 
* INPUT : br_485 
* OUTPUT: data_486 
* INPUT : bl_486 
* INPUT : br_486 
* OUTPUT: data_487 
* INPUT : bl_487 
* INPUT : br_487 
* OUTPUT: data_488 
* INPUT : bl_488 
* INPUT : br_488 
* OUTPUT: data_489 
* INPUT : bl_489 
* INPUT : br_489 
* OUTPUT: data_490 
* INPUT : bl_490 
* INPUT : br_490 
* OUTPUT: data_491 
* INPUT : bl_491 
* INPUT : br_491 
* OUTPUT: data_492 
* INPUT : bl_492 
* INPUT : br_492 
* OUTPUT: data_493 
* INPUT : bl_493 
* INPUT : br_493 
* OUTPUT: data_494 
* INPUT : bl_494 
* INPUT : br_494 
* OUTPUT: data_495 
* INPUT : bl_495 
* INPUT : br_495 
* OUTPUT: data_496 
* INPUT : bl_496 
* INPUT : br_496 
* OUTPUT: data_497 
* INPUT : bl_497 
* INPUT : br_497 
* OUTPUT: data_498 
* INPUT : bl_498 
* INPUT : br_498 
* OUTPUT: data_499 
* INPUT : bl_499 
* INPUT : br_499 
* OUTPUT: data_500 
* INPUT : bl_500 
* INPUT : br_500 
* OUTPUT: data_501 
* INPUT : bl_501 
* INPUT : br_501 
* OUTPUT: data_502 
* INPUT : bl_502 
* INPUT : br_502 
* OUTPUT: data_503 
* INPUT : bl_503 
* INPUT : br_503 
* OUTPUT: data_504 
* INPUT : bl_504 
* INPUT : br_504 
* OUTPUT: data_505 
* INPUT : bl_505 
* INPUT : br_505 
* OUTPUT: data_506 
* INPUT : bl_506 
* INPUT : br_506 
* OUTPUT: data_507 
* INPUT : bl_507 
* INPUT : br_507 
* OUTPUT: data_508 
* INPUT : bl_508 
* INPUT : br_508 
* OUTPUT: data_509 
* INPUT : bl_509 
* INPUT : br_509 
* OUTPUT: data_510 
* INPUT : bl_510 
* INPUT : br_510 
* OUTPUT: data_511 
* INPUT : bl_511 
* INPUT : br_511 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* words_per_row: 1
Xsa_d0
+ bl_0 br_0 data_0 en vdd gnd
+ sense_amp
Xsa_d1
+ bl_1 br_1 data_1 en vdd gnd
+ sense_amp
Xsa_d2
+ bl_2 br_2 data_2 en vdd gnd
+ sense_amp
Xsa_d3
+ bl_3 br_3 data_3 en vdd gnd
+ sense_amp
Xsa_d4
+ bl_4 br_4 data_4 en vdd gnd
+ sense_amp
Xsa_d5
+ bl_5 br_5 data_5 en vdd gnd
+ sense_amp
Xsa_d6
+ bl_6 br_6 data_6 en vdd gnd
+ sense_amp
Xsa_d7
+ bl_7 br_7 data_7 en vdd gnd
+ sense_amp
Xsa_d8
+ bl_8 br_8 data_8 en vdd gnd
+ sense_amp
Xsa_d9
+ bl_9 br_9 data_9 en vdd gnd
+ sense_amp
Xsa_d10
+ bl_10 br_10 data_10 en vdd gnd
+ sense_amp
Xsa_d11
+ bl_11 br_11 data_11 en vdd gnd
+ sense_amp
Xsa_d12
+ bl_12 br_12 data_12 en vdd gnd
+ sense_amp
Xsa_d13
+ bl_13 br_13 data_13 en vdd gnd
+ sense_amp
Xsa_d14
+ bl_14 br_14 data_14 en vdd gnd
+ sense_amp
Xsa_d15
+ bl_15 br_15 data_15 en vdd gnd
+ sense_amp
Xsa_d16
+ bl_16 br_16 data_16 en vdd gnd
+ sense_amp
Xsa_d17
+ bl_17 br_17 data_17 en vdd gnd
+ sense_amp
Xsa_d18
+ bl_18 br_18 data_18 en vdd gnd
+ sense_amp
Xsa_d19
+ bl_19 br_19 data_19 en vdd gnd
+ sense_amp
Xsa_d20
+ bl_20 br_20 data_20 en vdd gnd
+ sense_amp
Xsa_d21
+ bl_21 br_21 data_21 en vdd gnd
+ sense_amp
Xsa_d22
+ bl_22 br_22 data_22 en vdd gnd
+ sense_amp
Xsa_d23
+ bl_23 br_23 data_23 en vdd gnd
+ sense_amp
Xsa_d24
+ bl_24 br_24 data_24 en vdd gnd
+ sense_amp
Xsa_d25
+ bl_25 br_25 data_25 en vdd gnd
+ sense_amp
Xsa_d26
+ bl_26 br_26 data_26 en vdd gnd
+ sense_amp
Xsa_d27
+ bl_27 br_27 data_27 en vdd gnd
+ sense_amp
Xsa_d28
+ bl_28 br_28 data_28 en vdd gnd
+ sense_amp
Xsa_d29
+ bl_29 br_29 data_29 en vdd gnd
+ sense_amp
Xsa_d30
+ bl_30 br_30 data_30 en vdd gnd
+ sense_amp
Xsa_d31
+ bl_31 br_31 data_31 en vdd gnd
+ sense_amp
Xsa_d32
+ bl_32 br_32 data_32 en vdd gnd
+ sense_amp
Xsa_d33
+ bl_33 br_33 data_33 en vdd gnd
+ sense_amp
Xsa_d34
+ bl_34 br_34 data_34 en vdd gnd
+ sense_amp
Xsa_d35
+ bl_35 br_35 data_35 en vdd gnd
+ sense_amp
Xsa_d36
+ bl_36 br_36 data_36 en vdd gnd
+ sense_amp
Xsa_d37
+ bl_37 br_37 data_37 en vdd gnd
+ sense_amp
Xsa_d38
+ bl_38 br_38 data_38 en vdd gnd
+ sense_amp
Xsa_d39
+ bl_39 br_39 data_39 en vdd gnd
+ sense_amp
Xsa_d40
+ bl_40 br_40 data_40 en vdd gnd
+ sense_amp
Xsa_d41
+ bl_41 br_41 data_41 en vdd gnd
+ sense_amp
Xsa_d42
+ bl_42 br_42 data_42 en vdd gnd
+ sense_amp
Xsa_d43
+ bl_43 br_43 data_43 en vdd gnd
+ sense_amp
Xsa_d44
+ bl_44 br_44 data_44 en vdd gnd
+ sense_amp
Xsa_d45
+ bl_45 br_45 data_45 en vdd gnd
+ sense_amp
Xsa_d46
+ bl_46 br_46 data_46 en vdd gnd
+ sense_amp
Xsa_d47
+ bl_47 br_47 data_47 en vdd gnd
+ sense_amp
Xsa_d48
+ bl_48 br_48 data_48 en vdd gnd
+ sense_amp
Xsa_d49
+ bl_49 br_49 data_49 en vdd gnd
+ sense_amp
Xsa_d50
+ bl_50 br_50 data_50 en vdd gnd
+ sense_amp
Xsa_d51
+ bl_51 br_51 data_51 en vdd gnd
+ sense_amp
Xsa_d52
+ bl_52 br_52 data_52 en vdd gnd
+ sense_amp
Xsa_d53
+ bl_53 br_53 data_53 en vdd gnd
+ sense_amp
Xsa_d54
+ bl_54 br_54 data_54 en vdd gnd
+ sense_amp
Xsa_d55
+ bl_55 br_55 data_55 en vdd gnd
+ sense_amp
Xsa_d56
+ bl_56 br_56 data_56 en vdd gnd
+ sense_amp
Xsa_d57
+ bl_57 br_57 data_57 en vdd gnd
+ sense_amp
Xsa_d58
+ bl_58 br_58 data_58 en vdd gnd
+ sense_amp
Xsa_d59
+ bl_59 br_59 data_59 en vdd gnd
+ sense_amp
Xsa_d60
+ bl_60 br_60 data_60 en vdd gnd
+ sense_amp
Xsa_d61
+ bl_61 br_61 data_61 en vdd gnd
+ sense_amp
Xsa_d62
+ bl_62 br_62 data_62 en vdd gnd
+ sense_amp
Xsa_d63
+ bl_63 br_63 data_63 en vdd gnd
+ sense_amp
Xsa_d64
+ bl_64 br_64 data_64 en vdd gnd
+ sense_amp
Xsa_d65
+ bl_65 br_65 data_65 en vdd gnd
+ sense_amp
Xsa_d66
+ bl_66 br_66 data_66 en vdd gnd
+ sense_amp
Xsa_d67
+ bl_67 br_67 data_67 en vdd gnd
+ sense_amp
Xsa_d68
+ bl_68 br_68 data_68 en vdd gnd
+ sense_amp
Xsa_d69
+ bl_69 br_69 data_69 en vdd gnd
+ sense_amp
Xsa_d70
+ bl_70 br_70 data_70 en vdd gnd
+ sense_amp
Xsa_d71
+ bl_71 br_71 data_71 en vdd gnd
+ sense_amp
Xsa_d72
+ bl_72 br_72 data_72 en vdd gnd
+ sense_amp
Xsa_d73
+ bl_73 br_73 data_73 en vdd gnd
+ sense_amp
Xsa_d74
+ bl_74 br_74 data_74 en vdd gnd
+ sense_amp
Xsa_d75
+ bl_75 br_75 data_75 en vdd gnd
+ sense_amp
Xsa_d76
+ bl_76 br_76 data_76 en vdd gnd
+ sense_amp
Xsa_d77
+ bl_77 br_77 data_77 en vdd gnd
+ sense_amp
Xsa_d78
+ bl_78 br_78 data_78 en vdd gnd
+ sense_amp
Xsa_d79
+ bl_79 br_79 data_79 en vdd gnd
+ sense_amp
Xsa_d80
+ bl_80 br_80 data_80 en vdd gnd
+ sense_amp
Xsa_d81
+ bl_81 br_81 data_81 en vdd gnd
+ sense_amp
Xsa_d82
+ bl_82 br_82 data_82 en vdd gnd
+ sense_amp
Xsa_d83
+ bl_83 br_83 data_83 en vdd gnd
+ sense_amp
Xsa_d84
+ bl_84 br_84 data_84 en vdd gnd
+ sense_amp
Xsa_d85
+ bl_85 br_85 data_85 en vdd gnd
+ sense_amp
Xsa_d86
+ bl_86 br_86 data_86 en vdd gnd
+ sense_amp
Xsa_d87
+ bl_87 br_87 data_87 en vdd gnd
+ sense_amp
Xsa_d88
+ bl_88 br_88 data_88 en vdd gnd
+ sense_amp
Xsa_d89
+ bl_89 br_89 data_89 en vdd gnd
+ sense_amp
Xsa_d90
+ bl_90 br_90 data_90 en vdd gnd
+ sense_amp
Xsa_d91
+ bl_91 br_91 data_91 en vdd gnd
+ sense_amp
Xsa_d92
+ bl_92 br_92 data_92 en vdd gnd
+ sense_amp
Xsa_d93
+ bl_93 br_93 data_93 en vdd gnd
+ sense_amp
Xsa_d94
+ bl_94 br_94 data_94 en vdd gnd
+ sense_amp
Xsa_d95
+ bl_95 br_95 data_95 en vdd gnd
+ sense_amp
Xsa_d96
+ bl_96 br_96 data_96 en vdd gnd
+ sense_amp
Xsa_d97
+ bl_97 br_97 data_97 en vdd gnd
+ sense_amp
Xsa_d98
+ bl_98 br_98 data_98 en vdd gnd
+ sense_amp
Xsa_d99
+ bl_99 br_99 data_99 en vdd gnd
+ sense_amp
Xsa_d100
+ bl_100 br_100 data_100 en vdd gnd
+ sense_amp
Xsa_d101
+ bl_101 br_101 data_101 en vdd gnd
+ sense_amp
Xsa_d102
+ bl_102 br_102 data_102 en vdd gnd
+ sense_amp
Xsa_d103
+ bl_103 br_103 data_103 en vdd gnd
+ sense_amp
Xsa_d104
+ bl_104 br_104 data_104 en vdd gnd
+ sense_amp
Xsa_d105
+ bl_105 br_105 data_105 en vdd gnd
+ sense_amp
Xsa_d106
+ bl_106 br_106 data_106 en vdd gnd
+ sense_amp
Xsa_d107
+ bl_107 br_107 data_107 en vdd gnd
+ sense_amp
Xsa_d108
+ bl_108 br_108 data_108 en vdd gnd
+ sense_amp
Xsa_d109
+ bl_109 br_109 data_109 en vdd gnd
+ sense_amp
Xsa_d110
+ bl_110 br_110 data_110 en vdd gnd
+ sense_amp
Xsa_d111
+ bl_111 br_111 data_111 en vdd gnd
+ sense_amp
Xsa_d112
+ bl_112 br_112 data_112 en vdd gnd
+ sense_amp
Xsa_d113
+ bl_113 br_113 data_113 en vdd gnd
+ sense_amp
Xsa_d114
+ bl_114 br_114 data_114 en vdd gnd
+ sense_amp
Xsa_d115
+ bl_115 br_115 data_115 en vdd gnd
+ sense_amp
Xsa_d116
+ bl_116 br_116 data_116 en vdd gnd
+ sense_amp
Xsa_d117
+ bl_117 br_117 data_117 en vdd gnd
+ sense_amp
Xsa_d118
+ bl_118 br_118 data_118 en vdd gnd
+ sense_amp
Xsa_d119
+ bl_119 br_119 data_119 en vdd gnd
+ sense_amp
Xsa_d120
+ bl_120 br_120 data_120 en vdd gnd
+ sense_amp
Xsa_d121
+ bl_121 br_121 data_121 en vdd gnd
+ sense_amp
Xsa_d122
+ bl_122 br_122 data_122 en vdd gnd
+ sense_amp
Xsa_d123
+ bl_123 br_123 data_123 en vdd gnd
+ sense_amp
Xsa_d124
+ bl_124 br_124 data_124 en vdd gnd
+ sense_amp
Xsa_d125
+ bl_125 br_125 data_125 en vdd gnd
+ sense_amp
Xsa_d126
+ bl_126 br_126 data_126 en vdd gnd
+ sense_amp
Xsa_d127
+ bl_127 br_127 data_127 en vdd gnd
+ sense_amp
Xsa_d128
+ bl_128 br_128 data_128 en vdd gnd
+ sense_amp
Xsa_d129
+ bl_129 br_129 data_129 en vdd gnd
+ sense_amp
Xsa_d130
+ bl_130 br_130 data_130 en vdd gnd
+ sense_amp
Xsa_d131
+ bl_131 br_131 data_131 en vdd gnd
+ sense_amp
Xsa_d132
+ bl_132 br_132 data_132 en vdd gnd
+ sense_amp
Xsa_d133
+ bl_133 br_133 data_133 en vdd gnd
+ sense_amp
Xsa_d134
+ bl_134 br_134 data_134 en vdd gnd
+ sense_amp
Xsa_d135
+ bl_135 br_135 data_135 en vdd gnd
+ sense_amp
Xsa_d136
+ bl_136 br_136 data_136 en vdd gnd
+ sense_amp
Xsa_d137
+ bl_137 br_137 data_137 en vdd gnd
+ sense_amp
Xsa_d138
+ bl_138 br_138 data_138 en vdd gnd
+ sense_amp
Xsa_d139
+ bl_139 br_139 data_139 en vdd gnd
+ sense_amp
Xsa_d140
+ bl_140 br_140 data_140 en vdd gnd
+ sense_amp
Xsa_d141
+ bl_141 br_141 data_141 en vdd gnd
+ sense_amp
Xsa_d142
+ bl_142 br_142 data_142 en vdd gnd
+ sense_amp
Xsa_d143
+ bl_143 br_143 data_143 en vdd gnd
+ sense_amp
Xsa_d144
+ bl_144 br_144 data_144 en vdd gnd
+ sense_amp
Xsa_d145
+ bl_145 br_145 data_145 en vdd gnd
+ sense_amp
Xsa_d146
+ bl_146 br_146 data_146 en vdd gnd
+ sense_amp
Xsa_d147
+ bl_147 br_147 data_147 en vdd gnd
+ sense_amp
Xsa_d148
+ bl_148 br_148 data_148 en vdd gnd
+ sense_amp
Xsa_d149
+ bl_149 br_149 data_149 en vdd gnd
+ sense_amp
Xsa_d150
+ bl_150 br_150 data_150 en vdd gnd
+ sense_amp
Xsa_d151
+ bl_151 br_151 data_151 en vdd gnd
+ sense_amp
Xsa_d152
+ bl_152 br_152 data_152 en vdd gnd
+ sense_amp
Xsa_d153
+ bl_153 br_153 data_153 en vdd gnd
+ sense_amp
Xsa_d154
+ bl_154 br_154 data_154 en vdd gnd
+ sense_amp
Xsa_d155
+ bl_155 br_155 data_155 en vdd gnd
+ sense_amp
Xsa_d156
+ bl_156 br_156 data_156 en vdd gnd
+ sense_amp
Xsa_d157
+ bl_157 br_157 data_157 en vdd gnd
+ sense_amp
Xsa_d158
+ bl_158 br_158 data_158 en vdd gnd
+ sense_amp
Xsa_d159
+ bl_159 br_159 data_159 en vdd gnd
+ sense_amp
Xsa_d160
+ bl_160 br_160 data_160 en vdd gnd
+ sense_amp
Xsa_d161
+ bl_161 br_161 data_161 en vdd gnd
+ sense_amp
Xsa_d162
+ bl_162 br_162 data_162 en vdd gnd
+ sense_amp
Xsa_d163
+ bl_163 br_163 data_163 en vdd gnd
+ sense_amp
Xsa_d164
+ bl_164 br_164 data_164 en vdd gnd
+ sense_amp
Xsa_d165
+ bl_165 br_165 data_165 en vdd gnd
+ sense_amp
Xsa_d166
+ bl_166 br_166 data_166 en vdd gnd
+ sense_amp
Xsa_d167
+ bl_167 br_167 data_167 en vdd gnd
+ sense_amp
Xsa_d168
+ bl_168 br_168 data_168 en vdd gnd
+ sense_amp
Xsa_d169
+ bl_169 br_169 data_169 en vdd gnd
+ sense_amp
Xsa_d170
+ bl_170 br_170 data_170 en vdd gnd
+ sense_amp
Xsa_d171
+ bl_171 br_171 data_171 en vdd gnd
+ sense_amp
Xsa_d172
+ bl_172 br_172 data_172 en vdd gnd
+ sense_amp
Xsa_d173
+ bl_173 br_173 data_173 en vdd gnd
+ sense_amp
Xsa_d174
+ bl_174 br_174 data_174 en vdd gnd
+ sense_amp
Xsa_d175
+ bl_175 br_175 data_175 en vdd gnd
+ sense_amp
Xsa_d176
+ bl_176 br_176 data_176 en vdd gnd
+ sense_amp
Xsa_d177
+ bl_177 br_177 data_177 en vdd gnd
+ sense_amp
Xsa_d178
+ bl_178 br_178 data_178 en vdd gnd
+ sense_amp
Xsa_d179
+ bl_179 br_179 data_179 en vdd gnd
+ sense_amp
Xsa_d180
+ bl_180 br_180 data_180 en vdd gnd
+ sense_amp
Xsa_d181
+ bl_181 br_181 data_181 en vdd gnd
+ sense_amp
Xsa_d182
+ bl_182 br_182 data_182 en vdd gnd
+ sense_amp
Xsa_d183
+ bl_183 br_183 data_183 en vdd gnd
+ sense_amp
Xsa_d184
+ bl_184 br_184 data_184 en vdd gnd
+ sense_amp
Xsa_d185
+ bl_185 br_185 data_185 en vdd gnd
+ sense_amp
Xsa_d186
+ bl_186 br_186 data_186 en vdd gnd
+ sense_amp
Xsa_d187
+ bl_187 br_187 data_187 en vdd gnd
+ sense_amp
Xsa_d188
+ bl_188 br_188 data_188 en vdd gnd
+ sense_amp
Xsa_d189
+ bl_189 br_189 data_189 en vdd gnd
+ sense_amp
Xsa_d190
+ bl_190 br_190 data_190 en vdd gnd
+ sense_amp
Xsa_d191
+ bl_191 br_191 data_191 en vdd gnd
+ sense_amp
Xsa_d192
+ bl_192 br_192 data_192 en vdd gnd
+ sense_amp
Xsa_d193
+ bl_193 br_193 data_193 en vdd gnd
+ sense_amp
Xsa_d194
+ bl_194 br_194 data_194 en vdd gnd
+ sense_amp
Xsa_d195
+ bl_195 br_195 data_195 en vdd gnd
+ sense_amp
Xsa_d196
+ bl_196 br_196 data_196 en vdd gnd
+ sense_amp
Xsa_d197
+ bl_197 br_197 data_197 en vdd gnd
+ sense_amp
Xsa_d198
+ bl_198 br_198 data_198 en vdd gnd
+ sense_amp
Xsa_d199
+ bl_199 br_199 data_199 en vdd gnd
+ sense_amp
Xsa_d200
+ bl_200 br_200 data_200 en vdd gnd
+ sense_amp
Xsa_d201
+ bl_201 br_201 data_201 en vdd gnd
+ sense_amp
Xsa_d202
+ bl_202 br_202 data_202 en vdd gnd
+ sense_amp
Xsa_d203
+ bl_203 br_203 data_203 en vdd gnd
+ sense_amp
Xsa_d204
+ bl_204 br_204 data_204 en vdd gnd
+ sense_amp
Xsa_d205
+ bl_205 br_205 data_205 en vdd gnd
+ sense_amp
Xsa_d206
+ bl_206 br_206 data_206 en vdd gnd
+ sense_amp
Xsa_d207
+ bl_207 br_207 data_207 en vdd gnd
+ sense_amp
Xsa_d208
+ bl_208 br_208 data_208 en vdd gnd
+ sense_amp
Xsa_d209
+ bl_209 br_209 data_209 en vdd gnd
+ sense_amp
Xsa_d210
+ bl_210 br_210 data_210 en vdd gnd
+ sense_amp
Xsa_d211
+ bl_211 br_211 data_211 en vdd gnd
+ sense_amp
Xsa_d212
+ bl_212 br_212 data_212 en vdd gnd
+ sense_amp
Xsa_d213
+ bl_213 br_213 data_213 en vdd gnd
+ sense_amp
Xsa_d214
+ bl_214 br_214 data_214 en vdd gnd
+ sense_amp
Xsa_d215
+ bl_215 br_215 data_215 en vdd gnd
+ sense_amp
Xsa_d216
+ bl_216 br_216 data_216 en vdd gnd
+ sense_amp
Xsa_d217
+ bl_217 br_217 data_217 en vdd gnd
+ sense_amp
Xsa_d218
+ bl_218 br_218 data_218 en vdd gnd
+ sense_amp
Xsa_d219
+ bl_219 br_219 data_219 en vdd gnd
+ sense_amp
Xsa_d220
+ bl_220 br_220 data_220 en vdd gnd
+ sense_amp
Xsa_d221
+ bl_221 br_221 data_221 en vdd gnd
+ sense_amp
Xsa_d222
+ bl_222 br_222 data_222 en vdd gnd
+ sense_amp
Xsa_d223
+ bl_223 br_223 data_223 en vdd gnd
+ sense_amp
Xsa_d224
+ bl_224 br_224 data_224 en vdd gnd
+ sense_amp
Xsa_d225
+ bl_225 br_225 data_225 en vdd gnd
+ sense_amp
Xsa_d226
+ bl_226 br_226 data_226 en vdd gnd
+ sense_amp
Xsa_d227
+ bl_227 br_227 data_227 en vdd gnd
+ sense_amp
Xsa_d228
+ bl_228 br_228 data_228 en vdd gnd
+ sense_amp
Xsa_d229
+ bl_229 br_229 data_229 en vdd gnd
+ sense_amp
Xsa_d230
+ bl_230 br_230 data_230 en vdd gnd
+ sense_amp
Xsa_d231
+ bl_231 br_231 data_231 en vdd gnd
+ sense_amp
Xsa_d232
+ bl_232 br_232 data_232 en vdd gnd
+ sense_amp
Xsa_d233
+ bl_233 br_233 data_233 en vdd gnd
+ sense_amp
Xsa_d234
+ bl_234 br_234 data_234 en vdd gnd
+ sense_amp
Xsa_d235
+ bl_235 br_235 data_235 en vdd gnd
+ sense_amp
Xsa_d236
+ bl_236 br_236 data_236 en vdd gnd
+ sense_amp
Xsa_d237
+ bl_237 br_237 data_237 en vdd gnd
+ sense_amp
Xsa_d238
+ bl_238 br_238 data_238 en vdd gnd
+ sense_amp
Xsa_d239
+ bl_239 br_239 data_239 en vdd gnd
+ sense_amp
Xsa_d240
+ bl_240 br_240 data_240 en vdd gnd
+ sense_amp
Xsa_d241
+ bl_241 br_241 data_241 en vdd gnd
+ sense_amp
Xsa_d242
+ bl_242 br_242 data_242 en vdd gnd
+ sense_amp
Xsa_d243
+ bl_243 br_243 data_243 en vdd gnd
+ sense_amp
Xsa_d244
+ bl_244 br_244 data_244 en vdd gnd
+ sense_amp
Xsa_d245
+ bl_245 br_245 data_245 en vdd gnd
+ sense_amp
Xsa_d246
+ bl_246 br_246 data_246 en vdd gnd
+ sense_amp
Xsa_d247
+ bl_247 br_247 data_247 en vdd gnd
+ sense_amp
Xsa_d248
+ bl_248 br_248 data_248 en vdd gnd
+ sense_amp
Xsa_d249
+ bl_249 br_249 data_249 en vdd gnd
+ sense_amp
Xsa_d250
+ bl_250 br_250 data_250 en vdd gnd
+ sense_amp
Xsa_d251
+ bl_251 br_251 data_251 en vdd gnd
+ sense_amp
Xsa_d252
+ bl_252 br_252 data_252 en vdd gnd
+ sense_amp
Xsa_d253
+ bl_253 br_253 data_253 en vdd gnd
+ sense_amp
Xsa_d254
+ bl_254 br_254 data_254 en vdd gnd
+ sense_amp
Xsa_d255
+ bl_255 br_255 data_255 en vdd gnd
+ sense_amp
Xsa_d256
+ bl_256 br_256 data_256 en vdd gnd
+ sense_amp
Xsa_d257
+ bl_257 br_257 data_257 en vdd gnd
+ sense_amp
Xsa_d258
+ bl_258 br_258 data_258 en vdd gnd
+ sense_amp
Xsa_d259
+ bl_259 br_259 data_259 en vdd gnd
+ sense_amp
Xsa_d260
+ bl_260 br_260 data_260 en vdd gnd
+ sense_amp
Xsa_d261
+ bl_261 br_261 data_261 en vdd gnd
+ sense_amp
Xsa_d262
+ bl_262 br_262 data_262 en vdd gnd
+ sense_amp
Xsa_d263
+ bl_263 br_263 data_263 en vdd gnd
+ sense_amp
Xsa_d264
+ bl_264 br_264 data_264 en vdd gnd
+ sense_amp
Xsa_d265
+ bl_265 br_265 data_265 en vdd gnd
+ sense_amp
Xsa_d266
+ bl_266 br_266 data_266 en vdd gnd
+ sense_amp
Xsa_d267
+ bl_267 br_267 data_267 en vdd gnd
+ sense_amp
Xsa_d268
+ bl_268 br_268 data_268 en vdd gnd
+ sense_amp
Xsa_d269
+ bl_269 br_269 data_269 en vdd gnd
+ sense_amp
Xsa_d270
+ bl_270 br_270 data_270 en vdd gnd
+ sense_amp
Xsa_d271
+ bl_271 br_271 data_271 en vdd gnd
+ sense_amp
Xsa_d272
+ bl_272 br_272 data_272 en vdd gnd
+ sense_amp
Xsa_d273
+ bl_273 br_273 data_273 en vdd gnd
+ sense_amp
Xsa_d274
+ bl_274 br_274 data_274 en vdd gnd
+ sense_amp
Xsa_d275
+ bl_275 br_275 data_275 en vdd gnd
+ sense_amp
Xsa_d276
+ bl_276 br_276 data_276 en vdd gnd
+ sense_amp
Xsa_d277
+ bl_277 br_277 data_277 en vdd gnd
+ sense_amp
Xsa_d278
+ bl_278 br_278 data_278 en vdd gnd
+ sense_amp
Xsa_d279
+ bl_279 br_279 data_279 en vdd gnd
+ sense_amp
Xsa_d280
+ bl_280 br_280 data_280 en vdd gnd
+ sense_amp
Xsa_d281
+ bl_281 br_281 data_281 en vdd gnd
+ sense_amp
Xsa_d282
+ bl_282 br_282 data_282 en vdd gnd
+ sense_amp
Xsa_d283
+ bl_283 br_283 data_283 en vdd gnd
+ sense_amp
Xsa_d284
+ bl_284 br_284 data_284 en vdd gnd
+ sense_amp
Xsa_d285
+ bl_285 br_285 data_285 en vdd gnd
+ sense_amp
Xsa_d286
+ bl_286 br_286 data_286 en vdd gnd
+ sense_amp
Xsa_d287
+ bl_287 br_287 data_287 en vdd gnd
+ sense_amp
Xsa_d288
+ bl_288 br_288 data_288 en vdd gnd
+ sense_amp
Xsa_d289
+ bl_289 br_289 data_289 en vdd gnd
+ sense_amp
Xsa_d290
+ bl_290 br_290 data_290 en vdd gnd
+ sense_amp
Xsa_d291
+ bl_291 br_291 data_291 en vdd gnd
+ sense_amp
Xsa_d292
+ bl_292 br_292 data_292 en vdd gnd
+ sense_amp
Xsa_d293
+ bl_293 br_293 data_293 en vdd gnd
+ sense_amp
Xsa_d294
+ bl_294 br_294 data_294 en vdd gnd
+ sense_amp
Xsa_d295
+ bl_295 br_295 data_295 en vdd gnd
+ sense_amp
Xsa_d296
+ bl_296 br_296 data_296 en vdd gnd
+ sense_amp
Xsa_d297
+ bl_297 br_297 data_297 en vdd gnd
+ sense_amp
Xsa_d298
+ bl_298 br_298 data_298 en vdd gnd
+ sense_amp
Xsa_d299
+ bl_299 br_299 data_299 en vdd gnd
+ sense_amp
Xsa_d300
+ bl_300 br_300 data_300 en vdd gnd
+ sense_amp
Xsa_d301
+ bl_301 br_301 data_301 en vdd gnd
+ sense_amp
Xsa_d302
+ bl_302 br_302 data_302 en vdd gnd
+ sense_amp
Xsa_d303
+ bl_303 br_303 data_303 en vdd gnd
+ sense_amp
Xsa_d304
+ bl_304 br_304 data_304 en vdd gnd
+ sense_amp
Xsa_d305
+ bl_305 br_305 data_305 en vdd gnd
+ sense_amp
Xsa_d306
+ bl_306 br_306 data_306 en vdd gnd
+ sense_amp
Xsa_d307
+ bl_307 br_307 data_307 en vdd gnd
+ sense_amp
Xsa_d308
+ bl_308 br_308 data_308 en vdd gnd
+ sense_amp
Xsa_d309
+ bl_309 br_309 data_309 en vdd gnd
+ sense_amp
Xsa_d310
+ bl_310 br_310 data_310 en vdd gnd
+ sense_amp
Xsa_d311
+ bl_311 br_311 data_311 en vdd gnd
+ sense_amp
Xsa_d312
+ bl_312 br_312 data_312 en vdd gnd
+ sense_amp
Xsa_d313
+ bl_313 br_313 data_313 en vdd gnd
+ sense_amp
Xsa_d314
+ bl_314 br_314 data_314 en vdd gnd
+ sense_amp
Xsa_d315
+ bl_315 br_315 data_315 en vdd gnd
+ sense_amp
Xsa_d316
+ bl_316 br_316 data_316 en vdd gnd
+ sense_amp
Xsa_d317
+ bl_317 br_317 data_317 en vdd gnd
+ sense_amp
Xsa_d318
+ bl_318 br_318 data_318 en vdd gnd
+ sense_amp
Xsa_d319
+ bl_319 br_319 data_319 en vdd gnd
+ sense_amp
Xsa_d320
+ bl_320 br_320 data_320 en vdd gnd
+ sense_amp
Xsa_d321
+ bl_321 br_321 data_321 en vdd gnd
+ sense_amp
Xsa_d322
+ bl_322 br_322 data_322 en vdd gnd
+ sense_amp
Xsa_d323
+ bl_323 br_323 data_323 en vdd gnd
+ sense_amp
Xsa_d324
+ bl_324 br_324 data_324 en vdd gnd
+ sense_amp
Xsa_d325
+ bl_325 br_325 data_325 en vdd gnd
+ sense_amp
Xsa_d326
+ bl_326 br_326 data_326 en vdd gnd
+ sense_amp
Xsa_d327
+ bl_327 br_327 data_327 en vdd gnd
+ sense_amp
Xsa_d328
+ bl_328 br_328 data_328 en vdd gnd
+ sense_amp
Xsa_d329
+ bl_329 br_329 data_329 en vdd gnd
+ sense_amp
Xsa_d330
+ bl_330 br_330 data_330 en vdd gnd
+ sense_amp
Xsa_d331
+ bl_331 br_331 data_331 en vdd gnd
+ sense_amp
Xsa_d332
+ bl_332 br_332 data_332 en vdd gnd
+ sense_amp
Xsa_d333
+ bl_333 br_333 data_333 en vdd gnd
+ sense_amp
Xsa_d334
+ bl_334 br_334 data_334 en vdd gnd
+ sense_amp
Xsa_d335
+ bl_335 br_335 data_335 en vdd gnd
+ sense_amp
Xsa_d336
+ bl_336 br_336 data_336 en vdd gnd
+ sense_amp
Xsa_d337
+ bl_337 br_337 data_337 en vdd gnd
+ sense_amp
Xsa_d338
+ bl_338 br_338 data_338 en vdd gnd
+ sense_amp
Xsa_d339
+ bl_339 br_339 data_339 en vdd gnd
+ sense_amp
Xsa_d340
+ bl_340 br_340 data_340 en vdd gnd
+ sense_amp
Xsa_d341
+ bl_341 br_341 data_341 en vdd gnd
+ sense_amp
Xsa_d342
+ bl_342 br_342 data_342 en vdd gnd
+ sense_amp
Xsa_d343
+ bl_343 br_343 data_343 en vdd gnd
+ sense_amp
Xsa_d344
+ bl_344 br_344 data_344 en vdd gnd
+ sense_amp
Xsa_d345
+ bl_345 br_345 data_345 en vdd gnd
+ sense_amp
Xsa_d346
+ bl_346 br_346 data_346 en vdd gnd
+ sense_amp
Xsa_d347
+ bl_347 br_347 data_347 en vdd gnd
+ sense_amp
Xsa_d348
+ bl_348 br_348 data_348 en vdd gnd
+ sense_amp
Xsa_d349
+ bl_349 br_349 data_349 en vdd gnd
+ sense_amp
Xsa_d350
+ bl_350 br_350 data_350 en vdd gnd
+ sense_amp
Xsa_d351
+ bl_351 br_351 data_351 en vdd gnd
+ sense_amp
Xsa_d352
+ bl_352 br_352 data_352 en vdd gnd
+ sense_amp
Xsa_d353
+ bl_353 br_353 data_353 en vdd gnd
+ sense_amp
Xsa_d354
+ bl_354 br_354 data_354 en vdd gnd
+ sense_amp
Xsa_d355
+ bl_355 br_355 data_355 en vdd gnd
+ sense_amp
Xsa_d356
+ bl_356 br_356 data_356 en vdd gnd
+ sense_amp
Xsa_d357
+ bl_357 br_357 data_357 en vdd gnd
+ sense_amp
Xsa_d358
+ bl_358 br_358 data_358 en vdd gnd
+ sense_amp
Xsa_d359
+ bl_359 br_359 data_359 en vdd gnd
+ sense_amp
Xsa_d360
+ bl_360 br_360 data_360 en vdd gnd
+ sense_amp
Xsa_d361
+ bl_361 br_361 data_361 en vdd gnd
+ sense_amp
Xsa_d362
+ bl_362 br_362 data_362 en vdd gnd
+ sense_amp
Xsa_d363
+ bl_363 br_363 data_363 en vdd gnd
+ sense_amp
Xsa_d364
+ bl_364 br_364 data_364 en vdd gnd
+ sense_amp
Xsa_d365
+ bl_365 br_365 data_365 en vdd gnd
+ sense_amp
Xsa_d366
+ bl_366 br_366 data_366 en vdd gnd
+ sense_amp
Xsa_d367
+ bl_367 br_367 data_367 en vdd gnd
+ sense_amp
Xsa_d368
+ bl_368 br_368 data_368 en vdd gnd
+ sense_amp
Xsa_d369
+ bl_369 br_369 data_369 en vdd gnd
+ sense_amp
Xsa_d370
+ bl_370 br_370 data_370 en vdd gnd
+ sense_amp
Xsa_d371
+ bl_371 br_371 data_371 en vdd gnd
+ sense_amp
Xsa_d372
+ bl_372 br_372 data_372 en vdd gnd
+ sense_amp
Xsa_d373
+ bl_373 br_373 data_373 en vdd gnd
+ sense_amp
Xsa_d374
+ bl_374 br_374 data_374 en vdd gnd
+ sense_amp
Xsa_d375
+ bl_375 br_375 data_375 en vdd gnd
+ sense_amp
Xsa_d376
+ bl_376 br_376 data_376 en vdd gnd
+ sense_amp
Xsa_d377
+ bl_377 br_377 data_377 en vdd gnd
+ sense_amp
Xsa_d378
+ bl_378 br_378 data_378 en vdd gnd
+ sense_amp
Xsa_d379
+ bl_379 br_379 data_379 en vdd gnd
+ sense_amp
Xsa_d380
+ bl_380 br_380 data_380 en vdd gnd
+ sense_amp
Xsa_d381
+ bl_381 br_381 data_381 en vdd gnd
+ sense_amp
Xsa_d382
+ bl_382 br_382 data_382 en vdd gnd
+ sense_amp
Xsa_d383
+ bl_383 br_383 data_383 en vdd gnd
+ sense_amp
Xsa_d384
+ bl_384 br_384 data_384 en vdd gnd
+ sense_amp
Xsa_d385
+ bl_385 br_385 data_385 en vdd gnd
+ sense_amp
Xsa_d386
+ bl_386 br_386 data_386 en vdd gnd
+ sense_amp
Xsa_d387
+ bl_387 br_387 data_387 en vdd gnd
+ sense_amp
Xsa_d388
+ bl_388 br_388 data_388 en vdd gnd
+ sense_amp
Xsa_d389
+ bl_389 br_389 data_389 en vdd gnd
+ sense_amp
Xsa_d390
+ bl_390 br_390 data_390 en vdd gnd
+ sense_amp
Xsa_d391
+ bl_391 br_391 data_391 en vdd gnd
+ sense_amp
Xsa_d392
+ bl_392 br_392 data_392 en vdd gnd
+ sense_amp
Xsa_d393
+ bl_393 br_393 data_393 en vdd gnd
+ sense_amp
Xsa_d394
+ bl_394 br_394 data_394 en vdd gnd
+ sense_amp
Xsa_d395
+ bl_395 br_395 data_395 en vdd gnd
+ sense_amp
Xsa_d396
+ bl_396 br_396 data_396 en vdd gnd
+ sense_amp
Xsa_d397
+ bl_397 br_397 data_397 en vdd gnd
+ sense_amp
Xsa_d398
+ bl_398 br_398 data_398 en vdd gnd
+ sense_amp
Xsa_d399
+ bl_399 br_399 data_399 en vdd gnd
+ sense_amp
Xsa_d400
+ bl_400 br_400 data_400 en vdd gnd
+ sense_amp
Xsa_d401
+ bl_401 br_401 data_401 en vdd gnd
+ sense_amp
Xsa_d402
+ bl_402 br_402 data_402 en vdd gnd
+ sense_amp
Xsa_d403
+ bl_403 br_403 data_403 en vdd gnd
+ sense_amp
Xsa_d404
+ bl_404 br_404 data_404 en vdd gnd
+ sense_amp
Xsa_d405
+ bl_405 br_405 data_405 en vdd gnd
+ sense_amp
Xsa_d406
+ bl_406 br_406 data_406 en vdd gnd
+ sense_amp
Xsa_d407
+ bl_407 br_407 data_407 en vdd gnd
+ sense_amp
Xsa_d408
+ bl_408 br_408 data_408 en vdd gnd
+ sense_amp
Xsa_d409
+ bl_409 br_409 data_409 en vdd gnd
+ sense_amp
Xsa_d410
+ bl_410 br_410 data_410 en vdd gnd
+ sense_amp
Xsa_d411
+ bl_411 br_411 data_411 en vdd gnd
+ sense_amp
Xsa_d412
+ bl_412 br_412 data_412 en vdd gnd
+ sense_amp
Xsa_d413
+ bl_413 br_413 data_413 en vdd gnd
+ sense_amp
Xsa_d414
+ bl_414 br_414 data_414 en vdd gnd
+ sense_amp
Xsa_d415
+ bl_415 br_415 data_415 en vdd gnd
+ sense_amp
Xsa_d416
+ bl_416 br_416 data_416 en vdd gnd
+ sense_amp
Xsa_d417
+ bl_417 br_417 data_417 en vdd gnd
+ sense_amp
Xsa_d418
+ bl_418 br_418 data_418 en vdd gnd
+ sense_amp
Xsa_d419
+ bl_419 br_419 data_419 en vdd gnd
+ sense_amp
Xsa_d420
+ bl_420 br_420 data_420 en vdd gnd
+ sense_amp
Xsa_d421
+ bl_421 br_421 data_421 en vdd gnd
+ sense_amp
Xsa_d422
+ bl_422 br_422 data_422 en vdd gnd
+ sense_amp
Xsa_d423
+ bl_423 br_423 data_423 en vdd gnd
+ sense_amp
Xsa_d424
+ bl_424 br_424 data_424 en vdd gnd
+ sense_amp
Xsa_d425
+ bl_425 br_425 data_425 en vdd gnd
+ sense_amp
Xsa_d426
+ bl_426 br_426 data_426 en vdd gnd
+ sense_amp
Xsa_d427
+ bl_427 br_427 data_427 en vdd gnd
+ sense_amp
Xsa_d428
+ bl_428 br_428 data_428 en vdd gnd
+ sense_amp
Xsa_d429
+ bl_429 br_429 data_429 en vdd gnd
+ sense_amp
Xsa_d430
+ bl_430 br_430 data_430 en vdd gnd
+ sense_amp
Xsa_d431
+ bl_431 br_431 data_431 en vdd gnd
+ sense_amp
Xsa_d432
+ bl_432 br_432 data_432 en vdd gnd
+ sense_amp
Xsa_d433
+ bl_433 br_433 data_433 en vdd gnd
+ sense_amp
Xsa_d434
+ bl_434 br_434 data_434 en vdd gnd
+ sense_amp
Xsa_d435
+ bl_435 br_435 data_435 en vdd gnd
+ sense_amp
Xsa_d436
+ bl_436 br_436 data_436 en vdd gnd
+ sense_amp
Xsa_d437
+ bl_437 br_437 data_437 en vdd gnd
+ sense_amp
Xsa_d438
+ bl_438 br_438 data_438 en vdd gnd
+ sense_amp
Xsa_d439
+ bl_439 br_439 data_439 en vdd gnd
+ sense_amp
Xsa_d440
+ bl_440 br_440 data_440 en vdd gnd
+ sense_amp
Xsa_d441
+ bl_441 br_441 data_441 en vdd gnd
+ sense_amp
Xsa_d442
+ bl_442 br_442 data_442 en vdd gnd
+ sense_amp
Xsa_d443
+ bl_443 br_443 data_443 en vdd gnd
+ sense_amp
Xsa_d444
+ bl_444 br_444 data_444 en vdd gnd
+ sense_amp
Xsa_d445
+ bl_445 br_445 data_445 en vdd gnd
+ sense_amp
Xsa_d446
+ bl_446 br_446 data_446 en vdd gnd
+ sense_amp
Xsa_d447
+ bl_447 br_447 data_447 en vdd gnd
+ sense_amp
Xsa_d448
+ bl_448 br_448 data_448 en vdd gnd
+ sense_amp
Xsa_d449
+ bl_449 br_449 data_449 en vdd gnd
+ sense_amp
Xsa_d450
+ bl_450 br_450 data_450 en vdd gnd
+ sense_amp
Xsa_d451
+ bl_451 br_451 data_451 en vdd gnd
+ sense_amp
Xsa_d452
+ bl_452 br_452 data_452 en vdd gnd
+ sense_amp
Xsa_d453
+ bl_453 br_453 data_453 en vdd gnd
+ sense_amp
Xsa_d454
+ bl_454 br_454 data_454 en vdd gnd
+ sense_amp
Xsa_d455
+ bl_455 br_455 data_455 en vdd gnd
+ sense_amp
Xsa_d456
+ bl_456 br_456 data_456 en vdd gnd
+ sense_amp
Xsa_d457
+ bl_457 br_457 data_457 en vdd gnd
+ sense_amp
Xsa_d458
+ bl_458 br_458 data_458 en vdd gnd
+ sense_amp
Xsa_d459
+ bl_459 br_459 data_459 en vdd gnd
+ sense_amp
Xsa_d460
+ bl_460 br_460 data_460 en vdd gnd
+ sense_amp
Xsa_d461
+ bl_461 br_461 data_461 en vdd gnd
+ sense_amp
Xsa_d462
+ bl_462 br_462 data_462 en vdd gnd
+ sense_amp
Xsa_d463
+ bl_463 br_463 data_463 en vdd gnd
+ sense_amp
Xsa_d464
+ bl_464 br_464 data_464 en vdd gnd
+ sense_amp
Xsa_d465
+ bl_465 br_465 data_465 en vdd gnd
+ sense_amp
Xsa_d466
+ bl_466 br_466 data_466 en vdd gnd
+ sense_amp
Xsa_d467
+ bl_467 br_467 data_467 en vdd gnd
+ sense_amp
Xsa_d468
+ bl_468 br_468 data_468 en vdd gnd
+ sense_amp
Xsa_d469
+ bl_469 br_469 data_469 en vdd gnd
+ sense_amp
Xsa_d470
+ bl_470 br_470 data_470 en vdd gnd
+ sense_amp
Xsa_d471
+ bl_471 br_471 data_471 en vdd gnd
+ sense_amp
Xsa_d472
+ bl_472 br_472 data_472 en vdd gnd
+ sense_amp
Xsa_d473
+ bl_473 br_473 data_473 en vdd gnd
+ sense_amp
Xsa_d474
+ bl_474 br_474 data_474 en vdd gnd
+ sense_amp
Xsa_d475
+ bl_475 br_475 data_475 en vdd gnd
+ sense_amp
Xsa_d476
+ bl_476 br_476 data_476 en vdd gnd
+ sense_amp
Xsa_d477
+ bl_477 br_477 data_477 en vdd gnd
+ sense_amp
Xsa_d478
+ bl_478 br_478 data_478 en vdd gnd
+ sense_amp
Xsa_d479
+ bl_479 br_479 data_479 en vdd gnd
+ sense_amp
Xsa_d480
+ bl_480 br_480 data_480 en vdd gnd
+ sense_amp
Xsa_d481
+ bl_481 br_481 data_481 en vdd gnd
+ sense_amp
Xsa_d482
+ bl_482 br_482 data_482 en vdd gnd
+ sense_amp
Xsa_d483
+ bl_483 br_483 data_483 en vdd gnd
+ sense_amp
Xsa_d484
+ bl_484 br_484 data_484 en vdd gnd
+ sense_amp
Xsa_d485
+ bl_485 br_485 data_485 en vdd gnd
+ sense_amp
Xsa_d486
+ bl_486 br_486 data_486 en vdd gnd
+ sense_amp
Xsa_d487
+ bl_487 br_487 data_487 en vdd gnd
+ sense_amp
Xsa_d488
+ bl_488 br_488 data_488 en vdd gnd
+ sense_amp
Xsa_d489
+ bl_489 br_489 data_489 en vdd gnd
+ sense_amp
Xsa_d490
+ bl_490 br_490 data_490 en vdd gnd
+ sense_amp
Xsa_d491
+ bl_491 br_491 data_491 en vdd gnd
+ sense_amp
Xsa_d492
+ bl_492 br_492 data_492 en vdd gnd
+ sense_amp
Xsa_d493
+ bl_493 br_493 data_493 en vdd gnd
+ sense_amp
Xsa_d494
+ bl_494 br_494 data_494 en vdd gnd
+ sense_amp
Xsa_d495
+ bl_495 br_495 data_495 en vdd gnd
+ sense_amp
Xsa_d496
+ bl_496 br_496 data_496 en vdd gnd
+ sense_amp
Xsa_d497
+ bl_497 br_497 data_497 en vdd gnd
+ sense_amp
Xsa_d498
+ bl_498 br_498 data_498 en vdd gnd
+ sense_amp
Xsa_d499
+ bl_499 br_499 data_499 en vdd gnd
+ sense_amp
Xsa_d500
+ bl_500 br_500 data_500 en vdd gnd
+ sense_amp
Xsa_d501
+ bl_501 br_501 data_501 en vdd gnd
+ sense_amp
Xsa_d502
+ bl_502 br_502 data_502 en vdd gnd
+ sense_amp
Xsa_d503
+ bl_503 br_503 data_503 en vdd gnd
+ sense_amp
Xsa_d504
+ bl_504 br_504 data_504 en vdd gnd
+ sense_amp
Xsa_d505
+ bl_505 br_505 data_505 en vdd gnd
+ sense_amp
Xsa_d506
+ bl_506 br_506 data_506 en vdd gnd
+ sense_amp
Xsa_d507
+ bl_507 br_507 data_507 en vdd gnd
+ sense_amp
Xsa_d508
+ bl_508 br_508 data_508 en vdd gnd
+ sense_amp
Xsa_d509
+ bl_509 br_509 data_509 en vdd gnd
+ sense_amp
Xsa_d510
+ bl_510 br_510 data_510 en vdd gnd
+ sense_amp
Xsa_d511
+ bl_511 br_511 data_511 en vdd gnd
+ sense_amp
.ENDS freepdk45_sram_1rw0r_45x512_sense_amp_array

.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pmos_vtg w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nmos_vtg w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pmos_vtg w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pmos_vtg w=360.000000n l=50.000000n
mout0N bl en int2 gnd nmos_vtg w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pmos_vtg w=360.000000n l=50.000000n
mout1N br en int4 gnd nmos_vtg w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nmos_vtg w=180.000000n l=50.000000n
.ENDS write_driver


.SUBCKT freepdk45_sram_1rw0r_45x512_write_driver_array
+ data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9
+ data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17
+ data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25
+ data_26 data_27 data_28 data_29 data_30 data_31 data_32 data_33
+ data_34 data_35 data_36 data_37 data_38 data_39 data_40 data_41
+ data_42 data_43 data_44 data_45 data_46 data_47 data_48 data_49
+ data_50 data_51 data_52 data_53 data_54 data_55 data_56 data_57
+ data_58 data_59 data_60 data_61 data_62 data_63 data_64 data_65
+ data_66 data_67 data_68 data_69 data_70 data_71 data_72 data_73
+ data_74 data_75 data_76 data_77 data_78 data_79 data_80 data_81
+ data_82 data_83 data_84 data_85 data_86 data_87 data_88 data_89
+ data_90 data_91 data_92 data_93 data_94 data_95 data_96 data_97
+ data_98 data_99 data_100 data_101 data_102 data_103 data_104 data_105
+ data_106 data_107 data_108 data_109 data_110 data_111 data_112
+ data_113 data_114 data_115 data_116 data_117 data_118 data_119
+ data_120 data_121 data_122 data_123 data_124 data_125 data_126
+ data_127 data_128 data_129 data_130 data_131 data_132 data_133
+ data_134 data_135 data_136 data_137 data_138 data_139 data_140
+ data_141 data_142 data_143 data_144 data_145 data_146 data_147
+ data_148 data_149 data_150 data_151 data_152 data_153 data_154
+ data_155 data_156 data_157 data_158 data_159 data_160 data_161
+ data_162 data_163 data_164 data_165 data_166 data_167 data_168
+ data_169 data_170 data_171 data_172 data_173 data_174 data_175
+ data_176 data_177 data_178 data_179 data_180 data_181 data_182
+ data_183 data_184 data_185 data_186 data_187 data_188 data_189
+ data_190 data_191 data_192 data_193 data_194 data_195 data_196
+ data_197 data_198 data_199 data_200 data_201 data_202 data_203
+ data_204 data_205 data_206 data_207 data_208 data_209 data_210
+ data_211 data_212 data_213 data_214 data_215 data_216 data_217
+ data_218 data_219 data_220 data_221 data_222 data_223 data_224
+ data_225 data_226 data_227 data_228 data_229 data_230 data_231
+ data_232 data_233 data_234 data_235 data_236 data_237 data_238
+ data_239 data_240 data_241 data_242 data_243 data_244 data_245
+ data_246 data_247 data_248 data_249 data_250 data_251 data_252
+ data_253 data_254 data_255 data_256 data_257 data_258 data_259
+ data_260 data_261 data_262 data_263 data_264 data_265 data_266
+ data_267 data_268 data_269 data_270 data_271 data_272 data_273
+ data_274 data_275 data_276 data_277 data_278 data_279 data_280
+ data_281 data_282 data_283 data_284 data_285 data_286 data_287
+ data_288 data_289 data_290 data_291 data_292 data_293 data_294
+ data_295 data_296 data_297 data_298 data_299 data_300 data_301
+ data_302 data_303 data_304 data_305 data_306 data_307 data_308
+ data_309 data_310 data_311 data_312 data_313 data_314 data_315
+ data_316 data_317 data_318 data_319 data_320 data_321 data_322
+ data_323 data_324 data_325 data_326 data_327 data_328 data_329
+ data_330 data_331 data_332 data_333 data_334 data_335 data_336
+ data_337 data_338 data_339 data_340 data_341 data_342 data_343
+ data_344 data_345 data_346 data_347 data_348 data_349 data_350
+ data_351 data_352 data_353 data_354 data_355 data_356 data_357
+ data_358 data_359 data_360 data_361 data_362 data_363 data_364
+ data_365 data_366 data_367 data_368 data_369 data_370 data_371
+ data_372 data_373 data_374 data_375 data_376 data_377 data_378
+ data_379 data_380 data_381 data_382 data_383 data_384 data_385
+ data_386 data_387 data_388 data_389 data_390 data_391 data_392
+ data_393 data_394 data_395 data_396 data_397 data_398 data_399
+ data_400 data_401 data_402 data_403 data_404 data_405 data_406
+ data_407 data_408 data_409 data_410 data_411 data_412 data_413
+ data_414 data_415 data_416 data_417 data_418 data_419 data_420
+ data_421 data_422 data_423 data_424 data_425 data_426 data_427
+ data_428 data_429 data_430 data_431 data_432 data_433 data_434
+ data_435 data_436 data_437 data_438 data_439 data_440 data_441
+ data_442 data_443 data_444 data_445 data_446 data_447 data_448
+ data_449 data_450 data_451 data_452 data_453 data_454 data_455
+ data_456 data_457 data_458 data_459 data_460 data_461 data_462
+ data_463 data_464 data_465 data_466 data_467 data_468 data_469
+ data_470 data_471 data_472 data_473 data_474 data_475 data_476
+ data_477 data_478 data_479 data_480 data_481 data_482 data_483
+ data_484 data_485 data_486 data_487 data_488 data_489 data_490
+ data_491 data_492 data_493 data_494 data_495 data_496 data_497
+ data_498 data_499 data_500 data_501 data_502 data_503 data_504
+ data_505 data_506 data_507 data_508 data_509 data_510 data_511 bl_0
+ br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7
+ br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13
+ br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18
+ bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24
+ br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29
+ bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35
+ br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40
+ bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46
+ br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51
+ bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57
+ br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62
+ bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68
+ br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73
+ bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79
+ br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84
+ bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90
+ br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95
+ bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101
+ br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106
+ br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111
+ br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116
+ br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121
+ br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126
+ br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131
+ br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136
+ br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141
+ br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146
+ br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151
+ br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156
+ br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161
+ br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166
+ br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171
+ br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176
+ br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181
+ br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186
+ br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191
+ br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196
+ br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201
+ br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206
+ br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211
+ br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216
+ br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221
+ br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226
+ br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231
+ br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236
+ br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241
+ br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246
+ br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251
+ br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 bl_256
+ br_256 bl_257 br_257 bl_258 br_258 bl_259 br_259 bl_260 br_260 bl_261
+ br_261 bl_262 br_262 bl_263 br_263 bl_264 br_264 bl_265 br_265 bl_266
+ br_266 bl_267 br_267 bl_268 br_268 bl_269 br_269 bl_270 br_270 bl_271
+ br_271 bl_272 br_272 bl_273 br_273 bl_274 br_274 bl_275 br_275 bl_276
+ br_276 bl_277 br_277 bl_278 br_278 bl_279 br_279 bl_280 br_280 bl_281
+ br_281 bl_282 br_282 bl_283 br_283 bl_284 br_284 bl_285 br_285 bl_286
+ br_286 bl_287 br_287 bl_288 br_288 bl_289 br_289 bl_290 br_290 bl_291
+ br_291 bl_292 br_292 bl_293 br_293 bl_294 br_294 bl_295 br_295 bl_296
+ br_296 bl_297 br_297 bl_298 br_298 bl_299 br_299 bl_300 br_300 bl_301
+ br_301 bl_302 br_302 bl_303 br_303 bl_304 br_304 bl_305 br_305 bl_306
+ br_306 bl_307 br_307 bl_308 br_308 bl_309 br_309 bl_310 br_310 bl_311
+ br_311 bl_312 br_312 bl_313 br_313 bl_314 br_314 bl_315 br_315 bl_316
+ br_316 bl_317 br_317 bl_318 br_318 bl_319 br_319 bl_320 br_320 bl_321
+ br_321 bl_322 br_322 bl_323 br_323 bl_324 br_324 bl_325 br_325 bl_326
+ br_326 bl_327 br_327 bl_328 br_328 bl_329 br_329 bl_330 br_330 bl_331
+ br_331 bl_332 br_332 bl_333 br_333 bl_334 br_334 bl_335 br_335 bl_336
+ br_336 bl_337 br_337 bl_338 br_338 bl_339 br_339 bl_340 br_340 bl_341
+ br_341 bl_342 br_342 bl_343 br_343 bl_344 br_344 bl_345 br_345 bl_346
+ br_346 bl_347 br_347 bl_348 br_348 bl_349 br_349 bl_350 br_350 bl_351
+ br_351 bl_352 br_352 bl_353 br_353 bl_354 br_354 bl_355 br_355 bl_356
+ br_356 bl_357 br_357 bl_358 br_358 bl_359 br_359 bl_360 br_360 bl_361
+ br_361 bl_362 br_362 bl_363 br_363 bl_364 br_364 bl_365 br_365 bl_366
+ br_366 bl_367 br_367 bl_368 br_368 bl_369 br_369 bl_370 br_370 bl_371
+ br_371 bl_372 br_372 bl_373 br_373 bl_374 br_374 bl_375 br_375 bl_376
+ br_376 bl_377 br_377 bl_378 br_378 bl_379 br_379 bl_380 br_380 bl_381
+ br_381 bl_382 br_382 bl_383 br_383 bl_384 br_384 bl_385 br_385 bl_386
+ br_386 bl_387 br_387 bl_388 br_388 bl_389 br_389 bl_390 br_390 bl_391
+ br_391 bl_392 br_392 bl_393 br_393 bl_394 br_394 bl_395 br_395 bl_396
+ br_396 bl_397 br_397 bl_398 br_398 bl_399 br_399 bl_400 br_400 bl_401
+ br_401 bl_402 br_402 bl_403 br_403 bl_404 br_404 bl_405 br_405 bl_406
+ br_406 bl_407 br_407 bl_408 br_408 bl_409 br_409 bl_410 br_410 bl_411
+ br_411 bl_412 br_412 bl_413 br_413 bl_414 br_414 bl_415 br_415 bl_416
+ br_416 bl_417 br_417 bl_418 br_418 bl_419 br_419 bl_420 br_420 bl_421
+ br_421 bl_422 br_422 bl_423 br_423 bl_424 br_424 bl_425 br_425 bl_426
+ br_426 bl_427 br_427 bl_428 br_428 bl_429 br_429 bl_430 br_430 bl_431
+ br_431 bl_432 br_432 bl_433 br_433 bl_434 br_434 bl_435 br_435 bl_436
+ br_436 bl_437 br_437 bl_438 br_438 bl_439 br_439 bl_440 br_440 bl_441
+ br_441 bl_442 br_442 bl_443 br_443 bl_444 br_444 bl_445 br_445 bl_446
+ br_446 bl_447 br_447 bl_448 br_448 bl_449 br_449 bl_450 br_450 bl_451
+ br_451 bl_452 br_452 bl_453 br_453 bl_454 br_454 bl_455 br_455 bl_456
+ br_456 bl_457 br_457 bl_458 br_458 bl_459 br_459 bl_460 br_460 bl_461
+ br_461 bl_462 br_462 bl_463 br_463 bl_464 br_464 bl_465 br_465 bl_466
+ br_466 bl_467 br_467 bl_468 br_468 bl_469 br_469 bl_470 br_470 bl_471
+ br_471 bl_472 br_472 bl_473 br_473 bl_474 br_474 bl_475 br_475 bl_476
+ br_476 bl_477 br_477 bl_478 br_478 bl_479 br_479 bl_480 br_480 bl_481
+ br_481 bl_482 br_482 bl_483 br_483 bl_484 br_484 bl_485 br_485 bl_486
+ br_486 bl_487 br_487 bl_488 br_488 bl_489 br_489 bl_490 br_490 bl_491
+ br_491 bl_492 br_492 bl_493 br_493 bl_494 br_494 bl_495 br_495 bl_496
+ br_496 bl_497 br_497 bl_498 br_498 bl_499 br_499 bl_500 br_500 bl_501
+ br_501 bl_502 br_502 bl_503 br_503 bl_504 br_504 bl_505 br_505 bl_506
+ br_506 bl_507 br_507 bl_508 br_508 bl_509 br_509 bl_510 br_510 bl_511
+ br_511 en vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* INPUT : data_32 
* INPUT : data_33 
* INPUT : data_34 
* INPUT : data_35 
* INPUT : data_36 
* INPUT : data_37 
* INPUT : data_38 
* INPUT : data_39 
* INPUT : data_40 
* INPUT : data_41 
* INPUT : data_42 
* INPUT : data_43 
* INPUT : data_44 
* INPUT : data_45 
* INPUT : data_46 
* INPUT : data_47 
* INPUT : data_48 
* INPUT : data_49 
* INPUT : data_50 
* INPUT : data_51 
* INPUT : data_52 
* INPUT : data_53 
* INPUT : data_54 
* INPUT : data_55 
* INPUT : data_56 
* INPUT : data_57 
* INPUT : data_58 
* INPUT : data_59 
* INPUT : data_60 
* INPUT : data_61 
* INPUT : data_62 
* INPUT : data_63 
* INPUT : data_64 
* INPUT : data_65 
* INPUT : data_66 
* INPUT : data_67 
* INPUT : data_68 
* INPUT : data_69 
* INPUT : data_70 
* INPUT : data_71 
* INPUT : data_72 
* INPUT : data_73 
* INPUT : data_74 
* INPUT : data_75 
* INPUT : data_76 
* INPUT : data_77 
* INPUT : data_78 
* INPUT : data_79 
* INPUT : data_80 
* INPUT : data_81 
* INPUT : data_82 
* INPUT : data_83 
* INPUT : data_84 
* INPUT : data_85 
* INPUT : data_86 
* INPUT : data_87 
* INPUT : data_88 
* INPUT : data_89 
* INPUT : data_90 
* INPUT : data_91 
* INPUT : data_92 
* INPUT : data_93 
* INPUT : data_94 
* INPUT : data_95 
* INPUT : data_96 
* INPUT : data_97 
* INPUT : data_98 
* INPUT : data_99 
* INPUT : data_100 
* INPUT : data_101 
* INPUT : data_102 
* INPUT : data_103 
* INPUT : data_104 
* INPUT : data_105 
* INPUT : data_106 
* INPUT : data_107 
* INPUT : data_108 
* INPUT : data_109 
* INPUT : data_110 
* INPUT : data_111 
* INPUT : data_112 
* INPUT : data_113 
* INPUT : data_114 
* INPUT : data_115 
* INPUT : data_116 
* INPUT : data_117 
* INPUT : data_118 
* INPUT : data_119 
* INPUT : data_120 
* INPUT : data_121 
* INPUT : data_122 
* INPUT : data_123 
* INPUT : data_124 
* INPUT : data_125 
* INPUT : data_126 
* INPUT : data_127 
* INPUT : data_128 
* INPUT : data_129 
* INPUT : data_130 
* INPUT : data_131 
* INPUT : data_132 
* INPUT : data_133 
* INPUT : data_134 
* INPUT : data_135 
* INPUT : data_136 
* INPUT : data_137 
* INPUT : data_138 
* INPUT : data_139 
* INPUT : data_140 
* INPUT : data_141 
* INPUT : data_142 
* INPUT : data_143 
* INPUT : data_144 
* INPUT : data_145 
* INPUT : data_146 
* INPUT : data_147 
* INPUT : data_148 
* INPUT : data_149 
* INPUT : data_150 
* INPUT : data_151 
* INPUT : data_152 
* INPUT : data_153 
* INPUT : data_154 
* INPUT : data_155 
* INPUT : data_156 
* INPUT : data_157 
* INPUT : data_158 
* INPUT : data_159 
* INPUT : data_160 
* INPUT : data_161 
* INPUT : data_162 
* INPUT : data_163 
* INPUT : data_164 
* INPUT : data_165 
* INPUT : data_166 
* INPUT : data_167 
* INPUT : data_168 
* INPUT : data_169 
* INPUT : data_170 
* INPUT : data_171 
* INPUT : data_172 
* INPUT : data_173 
* INPUT : data_174 
* INPUT : data_175 
* INPUT : data_176 
* INPUT : data_177 
* INPUT : data_178 
* INPUT : data_179 
* INPUT : data_180 
* INPUT : data_181 
* INPUT : data_182 
* INPUT : data_183 
* INPUT : data_184 
* INPUT : data_185 
* INPUT : data_186 
* INPUT : data_187 
* INPUT : data_188 
* INPUT : data_189 
* INPUT : data_190 
* INPUT : data_191 
* INPUT : data_192 
* INPUT : data_193 
* INPUT : data_194 
* INPUT : data_195 
* INPUT : data_196 
* INPUT : data_197 
* INPUT : data_198 
* INPUT : data_199 
* INPUT : data_200 
* INPUT : data_201 
* INPUT : data_202 
* INPUT : data_203 
* INPUT : data_204 
* INPUT : data_205 
* INPUT : data_206 
* INPUT : data_207 
* INPUT : data_208 
* INPUT : data_209 
* INPUT : data_210 
* INPUT : data_211 
* INPUT : data_212 
* INPUT : data_213 
* INPUT : data_214 
* INPUT : data_215 
* INPUT : data_216 
* INPUT : data_217 
* INPUT : data_218 
* INPUT : data_219 
* INPUT : data_220 
* INPUT : data_221 
* INPUT : data_222 
* INPUT : data_223 
* INPUT : data_224 
* INPUT : data_225 
* INPUT : data_226 
* INPUT : data_227 
* INPUT : data_228 
* INPUT : data_229 
* INPUT : data_230 
* INPUT : data_231 
* INPUT : data_232 
* INPUT : data_233 
* INPUT : data_234 
* INPUT : data_235 
* INPUT : data_236 
* INPUT : data_237 
* INPUT : data_238 
* INPUT : data_239 
* INPUT : data_240 
* INPUT : data_241 
* INPUT : data_242 
* INPUT : data_243 
* INPUT : data_244 
* INPUT : data_245 
* INPUT : data_246 
* INPUT : data_247 
* INPUT : data_248 
* INPUT : data_249 
* INPUT : data_250 
* INPUT : data_251 
* INPUT : data_252 
* INPUT : data_253 
* INPUT : data_254 
* INPUT : data_255 
* INPUT : data_256 
* INPUT : data_257 
* INPUT : data_258 
* INPUT : data_259 
* INPUT : data_260 
* INPUT : data_261 
* INPUT : data_262 
* INPUT : data_263 
* INPUT : data_264 
* INPUT : data_265 
* INPUT : data_266 
* INPUT : data_267 
* INPUT : data_268 
* INPUT : data_269 
* INPUT : data_270 
* INPUT : data_271 
* INPUT : data_272 
* INPUT : data_273 
* INPUT : data_274 
* INPUT : data_275 
* INPUT : data_276 
* INPUT : data_277 
* INPUT : data_278 
* INPUT : data_279 
* INPUT : data_280 
* INPUT : data_281 
* INPUT : data_282 
* INPUT : data_283 
* INPUT : data_284 
* INPUT : data_285 
* INPUT : data_286 
* INPUT : data_287 
* INPUT : data_288 
* INPUT : data_289 
* INPUT : data_290 
* INPUT : data_291 
* INPUT : data_292 
* INPUT : data_293 
* INPUT : data_294 
* INPUT : data_295 
* INPUT : data_296 
* INPUT : data_297 
* INPUT : data_298 
* INPUT : data_299 
* INPUT : data_300 
* INPUT : data_301 
* INPUT : data_302 
* INPUT : data_303 
* INPUT : data_304 
* INPUT : data_305 
* INPUT : data_306 
* INPUT : data_307 
* INPUT : data_308 
* INPUT : data_309 
* INPUT : data_310 
* INPUT : data_311 
* INPUT : data_312 
* INPUT : data_313 
* INPUT : data_314 
* INPUT : data_315 
* INPUT : data_316 
* INPUT : data_317 
* INPUT : data_318 
* INPUT : data_319 
* INPUT : data_320 
* INPUT : data_321 
* INPUT : data_322 
* INPUT : data_323 
* INPUT : data_324 
* INPUT : data_325 
* INPUT : data_326 
* INPUT : data_327 
* INPUT : data_328 
* INPUT : data_329 
* INPUT : data_330 
* INPUT : data_331 
* INPUT : data_332 
* INPUT : data_333 
* INPUT : data_334 
* INPUT : data_335 
* INPUT : data_336 
* INPUT : data_337 
* INPUT : data_338 
* INPUT : data_339 
* INPUT : data_340 
* INPUT : data_341 
* INPUT : data_342 
* INPUT : data_343 
* INPUT : data_344 
* INPUT : data_345 
* INPUT : data_346 
* INPUT : data_347 
* INPUT : data_348 
* INPUT : data_349 
* INPUT : data_350 
* INPUT : data_351 
* INPUT : data_352 
* INPUT : data_353 
* INPUT : data_354 
* INPUT : data_355 
* INPUT : data_356 
* INPUT : data_357 
* INPUT : data_358 
* INPUT : data_359 
* INPUT : data_360 
* INPUT : data_361 
* INPUT : data_362 
* INPUT : data_363 
* INPUT : data_364 
* INPUT : data_365 
* INPUT : data_366 
* INPUT : data_367 
* INPUT : data_368 
* INPUT : data_369 
* INPUT : data_370 
* INPUT : data_371 
* INPUT : data_372 
* INPUT : data_373 
* INPUT : data_374 
* INPUT : data_375 
* INPUT : data_376 
* INPUT : data_377 
* INPUT : data_378 
* INPUT : data_379 
* INPUT : data_380 
* INPUT : data_381 
* INPUT : data_382 
* INPUT : data_383 
* INPUT : data_384 
* INPUT : data_385 
* INPUT : data_386 
* INPUT : data_387 
* INPUT : data_388 
* INPUT : data_389 
* INPUT : data_390 
* INPUT : data_391 
* INPUT : data_392 
* INPUT : data_393 
* INPUT : data_394 
* INPUT : data_395 
* INPUT : data_396 
* INPUT : data_397 
* INPUT : data_398 
* INPUT : data_399 
* INPUT : data_400 
* INPUT : data_401 
* INPUT : data_402 
* INPUT : data_403 
* INPUT : data_404 
* INPUT : data_405 
* INPUT : data_406 
* INPUT : data_407 
* INPUT : data_408 
* INPUT : data_409 
* INPUT : data_410 
* INPUT : data_411 
* INPUT : data_412 
* INPUT : data_413 
* INPUT : data_414 
* INPUT : data_415 
* INPUT : data_416 
* INPUT : data_417 
* INPUT : data_418 
* INPUT : data_419 
* INPUT : data_420 
* INPUT : data_421 
* INPUT : data_422 
* INPUT : data_423 
* INPUT : data_424 
* INPUT : data_425 
* INPUT : data_426 
* INPUT : data_427 
* INPUT : data_428 
* INPUT : data_429 
* INPUT : data_430 
* INPUT : data_431 
* INPUT : data_432 
* INPUT : data_433 
* INPUT : data_434 
* INPUT : data_435 
* INPUT : data_436 
* INPUT : data_437 
* INPUT : data_438 
* INPUT : data_439 
* INPUT : data_440 
* INPUT : data_441 
* INPUT : data_442 
* INPUT : data_443 
* INPUT : data_444 
* INPUT : data_445 
* INPUT : data_446 
* INPUT : data_447 
* INPUT : data_448 
* INPUT : data_449 
* INPUT : data_450 
* INPUT : data_451 
* INPUT : data_452 
* INPUT : data_453 
* INPUT : data_454 
* INPUT : data_455 
* INPUT : data_456 
* INPUT : data_457 
* INPUT : data_458 
* INPUT : data_459 
* INPUT : data_460 
* INPUT : data_461 
* INPUT : data_462 
* INPUT : data_463 
* INPUT : data_464 
* INPUT : data_465 
* INPUT : data_466 
* INPUT : data_467 
* INPUT : data_468 
* INPUT : data_469 
* INPUT : data_470 
* INPUT : data_471 
* INPUT : data_472 
* INPUT : data_473 
* INPUT : data_474 
* INPUT : data_475 
* INPUT : data_476 
* INPUT : data_477 
* INPUT : data_478 
* INPUT : data_479 
* INPUT : data_480 
* INPUT : data_481 
* INPUT : data_482 
* INPUT : data_483 
* INPUT : data_484 
* INPUT : data_485 
* INPUT : data_486 
* INPUT : data_487 
* INPUT : data_488 
* INPUT : data_489 
* INPUT : data_490 
* INPUT : data_491 
* INPUT : data_492 
* INPUT : data_493 
* INPUT : data_494 
* INPUT : data_495 
* INPUT : data_496 
* INPUT : data_497 
* INPUT : data_498 
* INPUT : data_499 
* INPUT : data_500 
* INPUT : data_501 
* INPUT : data_502 
* INPUT : data_503 
* INPUT : data_504 
* INPUT : data_505 
* INPUT : data_506 
* INPUT : data_507 
* INPUT : data_508 
* INPUT : data_509 
* INPUT : data_510 
* INPUT : data_511 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* OUTPUT: bl_130 
* OUTPUT: br_130 
* OUTPUT: bl_131 
* OUTPUT: br_131 
* OUTPUT: bl_132 
* OUTPUT: br_132 
* OUTPUT: bl_133 
* OUTPUT: br_133 
* OUTPUT: bl_134 
* OUTPUT: br_134 
* OUTPUT: bl_135 
* OUTPUT: br_135 
* OUTPUT: bl_136 
* OUTPUT: br_136 
* OUTPUT: bl_137 
* OUTPUT: br_137 
* OUTPUT: bl_138 
* OUTPUT: br_138 
* OUTPUT: bl_139 
* OUTPUT: br_139 
* OUTPUT: bl_140 
* OUTPUT: br_140 
* OUTPUT: bl_141 
* OUTPUT: br_141 
* OUTPUT: bl_142 
* OUTPUT: br_142 
* OUTPUT: bl_143 
* OUTPUT: br_143 
* OUTPUT: bl_144 
* OUTPUT: br_144 
* OUTPUT: bl_145 
* OUTPUT: br_145 
* OUTPUT: bl_146 
* OUTPUT: br_146 
* OUTPUT: bl_147 
* OUTPUT: br_147 
* OUTPUT: bl_148 
* OUTPUT: br_148 
* OUTPUT: bl_149 
* OUTPUT: br_149 
* OUTPUT: bl_150 
* OUTPUT: br_150 
* OUTPUT: bl_151 
* OUTPUT: br_151 
* OUTPUT: bl_152 
* OUTPUT: br_152 
* OUTPUT: bl_153 
* OUTPUT: br_153 
* OUTPUT: bl_154 
* OUTPUT: br_154 
* OUTPUT: bl_155 
* OUTPUT: br_155 
* OUTPUT: bl_156 
* OUTPUT: br_156 
* OUTPUT: bl_157 
* OUTPUT: br_157 
* OUTPUT: bl_158 
* OUTPUT: br_158 
* OUTPUT: bl_159 
* OUTPUT: br_159 
* OUTPUT: bl_160 
* OUTPUT: br_160 
* OUTPUT: bl_161 
* OUTPUT: br_161 
* OUTPUT: bl_162 
* OUTPUT: br_162 
* OUTPUT: bl_163 
* OUTPUT: br_163 
* OUTPUT: bl_164 
* OUTPUT: br_164 
* OUTPUT: bl_165 
* OUTPUT: br_165 
* OUTPUT: bl_166 
* OUTPUT: br_166 
* OUTPUT: bl_167 
* OUTPUT: br_167 
* OUTPUT: bl_168 
* OUTPUT: br_168 
* OUTPUT: bl_169 
* OUTPUT: br_169 
* OUTPUT: bl_170 
* OUTPUT: br_170 
* OUTPUT: bl_171 
* OUTPUT: br_171 
* OUTPUT: bl_172 
* OUTPUT: br_172 
* OUTPUT: bl_173 
* OUTPUT: br_173 
* OUTPUT: bl_174 
* OUTPUT: br_174 
* OUTPUT: bl_175 
* OUTPUT: br_175 
* OUTPUT: bl_176 
* OUTPUT: br_176 
* OUTPUT: bl_177 
* OUTPUT: br_177 
* OUTPUT: bl_178 
* OUTPUT: br_178 
* OUTPUT: bl_179 
* OUTPUT: br_179 
* OUTPUT: bl_180 
* OUTPUT: br_180 
* OUTPUT: bl_181 
* OUTPUT: br_181 
* OUTPUT: bl_182 
* OUTPUT: br_182 
* OUTPUT: bl_183 
* OUTPUT: br_183 
* OUTPUT: bl_184 
* OUTPUT: br_184 
* OUTPUT: bl_185 
* OUTPUT: br_185 
* OUTPUT: bl_186 
* OUTPUT: br_186 
* OUTPUT: bl_187 
* OUTPUT: br_187 
* OUTPUT: bl_188 
* OUTPUT: br_188 
* OUTPUT: bl_189 
* OUTPUT: br_189 
* OUTPUT: bl_190 
* OUTPUT: br_190 
* OUTPUT: bl_191 
* OUTPUT: br_191 
* OUTPUT: bl_192 
* OUTPUT: br_192 
* OUTPUT: bl_193 
* OUTPUT: br_193 
* OUTPUT: bl_194 
* OUTPUT: br_194 
* OUTPUT: bl_195 
* OUTPUT: br_195 
* OUTPUT: bl_196 
* OUTPUT: br_196 
* OUTPUT: bl_197 
* OUTPUT: br_197 
* OUTPUT: bl_198 
* OUTPUT: br_198 
* OUTPUT: bl_199 
* OUTPUT: br_199 
* OUTPUT: bl_200 
* OUTPUT: br_200 
* OUTPUT: bl_201 
* OUTPUT: br_201 
* OUTPUT: bl_202 
* OUTPUT: br_202 
* OUTPUT: bl_203 
* OUTPUT: br_203 
* OUTPUT: bl_204 
* OUTPUT: br_204 
* OUTPUT: bl_205 
* OUTPUT: br_205 
* OUTPUT: bl_206 
* OUTPUT: br_206 
* OUTPUT: bl_207 
* OUTPUT: br_207 
* OUTPUT: bl_208 
* OUTPUT: br_208 
* OUTPUT: bl_209 
* OUTPUT: br_209 
* OUTPUT: bl_210 
* OUTPUT: br_210 
* OUTPUT: bl_211 
* OUTPUT: br_211 
* OUTPUT: bl_212 
* OUTPUT: br_212 
* OUTPUT: bl_213 
* OUTPUT: br_213 
* OUTPUT: bl_214 
* OUTPUT: br_214 
* OUTPUT: bl_215 
* OUTPUT: br_215 
* OUTPUT: bl_216 
* OUTPUT: br_216 
* OUTPUT: bl_217 
* OUTPUT: br_217 
* OUTPUT: bl_218 
* OUTPUT: br_218 
* OUTPUT: bl_219 
* OUTPUT: br_219 
* OUTPUT: bl_220 
* OUTPUT: br_220 
* OUTPUT: bl_221 
* OUTPUT: br_221 
* OUTPUT: bl_222 
* OUTPUT: br_222 
* OUTPUT: bl_223 
* OUTPUT: br_223 
* OUTPUT: bl_224 
* OUTPUT: br_224 
* OUTPUT: bl_225 
* OUTPUT: br_225 
* OUTPUT: bl_226 
* OUTPUT: br_226 
* OUTPUT: bl_227 
* OUTPUT: br_227 
* OUTPUT: bl_228 
* OUTPUT: br_228 
* OUTPUT: bl_229 
* OUTPUT: br_229 
* OUTPUT: bl_230 
* OUTPUT: br_230 
* OUTPUT: bl_231 
* OUTPUT: br_231 
* OUTPUT: bl_232 
* OUTPUT: br_232 
* OUTPUT: bl_233 
* OUTPUT: br_233 
* OUTPUT: bl_234 
* OUTPUT: br_234 
* OUTPUT: bl_235 
* OUTPUT: br_235 
* OUTPUT: bl_236 
* OUTPUT: br_236 
* OUTPUT: bl_237 
* OUTPUT: br_237 
* OUTPUT: bl_238 
* OUTPUT: br_238 
* OUTPUT: bl_239 
* OUTPUT: br_239 
* OUTPUT: bl_240 
* OUTPUT: br_240 
* OUTPUT: bl_241 
* OUTPUT: br_241 
* OUTPUT: bl_242 
* OUTPUT: br_242 
* OUTPUT: bl_243 
* OUTPUT: br_243 
* OUTPUT: bl_244 
* OUTPUT: br_244 
* OUTPUT: bl_245 
* OUTPUT: br_245 
* OUTPUT: bl_246 
* OUTPUT: br_246 
* OUTPUT: bl_247 
* OUTPUT: br_247 
* OUTPUT: bl_248 
* OUTPUT: br_248 
* OUTPUT: bl_249 
* OUTPUT: br_249 
* OUTPUT: bl_250 
* OUTPUT: br_250 
* OUTPUT: bl_251 
* OUTPUT: br_251 
* OUTPUT: bl_252 
* OUTPUT: br_252 
* OUTPUT: bl_253 
* OUTPUT: br_253 
* OUTPUT: bl_254 
* OUTPUT: br_254 
* OUTPUT: bl_255 
* OUTPUT: br_255 
* OUTPUT: bl_256 
* OUTPUT: br_256 
* OUTPUT: bl_257 
* OUTPUT: br_257 
* OUTPUT: bl_258 
* OUTPUT: br_258 
* OUTPUT: bl_259 
* OUTPUT: br_259 
* OUTPUT: bl_260 
* OUTPUT: br_260 
* OUTPUT: bl_261 
* OUTPUT: br_261 
* OUTPUT: bl_262 
* OUTPUT: br_262 
* OUTPUT: bl_263 
* OUTPUT: br_263 
* OUTPUT: bl_264 
* OUTPUT: br_264 
* OUTPUT: bl_265 
* OUTPUT: br_265 
* OUTPUT: bl_266 
* OUTPUT: br_266 
* OUTPUT: bl_267 
* OUTPUT: br_267 
* OUTPUT: bl_268 
* OUTPUT: br_268 
* OUTPUT: bl_269 
* OUTPUT: br_269 
* OUTPUT: bl_270 
* OUTPUT: br_270 
* OUTPUT: bl_271 
* OUTPUT: br_271 
* OUTPUT: bl_272 
* OUTPUT: br_272 
* OUTPUT: bl_273 
* OUTPUT: br_273 
* OUTPUT: bl_274 
* OUTPUT: br_274 
* OUTPUT: bl_275 
* OUTPUT: br_275 
* OUTPUT: bl_276 
* OUTPUT: br_276 
* OUTPUT: bl_277 
* OUTPUT: br_277 
* OUTPUT: bl_278 
* OUTPUT: br_278 
* OUTPUT: bl_279 
* OUTPUT: br_279 
* OUTPUT: bl_280 
* OUTPUT: br_280 
* OUTPUT: bl_281 
* OUTPUT: br_281 
* OUTPUT: bl_282 
* OUTPUT: br_282 
* OUTPUT: bl_283 
* OUTPUT: br_283 
* OUTPUT: bl_284 
* OUTPUT: br_284 
* OUTPUT: bl_285 
* OUTPUT: br_285 
* OUTPUT: bl_286 
* OUTPUT: br_286 
* OUTPUT: bl_287 
* OUTPUT: br_287 
* OUTPUT: bl_288 
* OUTPUT: br_288 
* OUTPUT: bl_289 
* OUTPUT: br_289 
* OUTPUT: bl_290 
* OUTPUT: br_290 
* OUTPUT: bl_291 
* OUTPUT: br_291 
* OUTPUT: bl_292 
* OUTPUT: br_292 
* OUTPUT: bl_293 
* OUTPUT: br_293 
* OUTPUT: bl_294 
* OUTPUT: br_294 
* OUTPUT: bl_295 
* OUTPUT: br_295 
* OUTPUT: bl_296 
* OUTPUT: br_296 
* OUTPUT: bl_297 
* OUTPUT: br_297 
* OUTPUT: bl_298 
* OUTPUT: br_298 
* OUTPUT: bl_299 
* OUTPUT: br_299 
* OUTPUT: bl_300 
* OUTPUT: br_300 
* OUTPUT: bl_301 
* OUTPUT: br_301 
* OUTPUT: bl_302 
* OUTPUT: br_302 
* OUTPUT: bl_303 
* OUTPUT: br_303 
* OUTPUT: bl_304 
* OUTPUT: br_304 
* OUTPUT: bl_305 
* OUTPUT: br_305 
* OUTPUT: bl_306 
* OUTPUT: br_306 
* OUTPUT: bl_307 
* OUTPUT: br_307 
* OUTPUT: bl_308 
* OUTPUT: br_308 
* OUTPUT: bl_309 
* OUTPUT: br_309 
* OUTPUT: bl_310 
* OUTPUT: br_310 
* OUTPUT: bl_311 
* OUTPUT: br_311 
* OUTPUT: bl_312 
* OUTPUT: br_312 
* OUTPUT: bl_313 
* OUTPUT: br_313 
* OUTPUT: bl_314 
* OUTPUT: br_314 
* OUTPUT: bl_315 
* OUTPUT: br_315 
* OUTPUT: bl_316 
* OUTPUT: br_316 
* OUTPUT: bl_317 
* OUTPUT: br_317 
* OUTPUT: bl_318 
* OUTPUT: br_318 
* OUTPUT: bl_319 
* OUTPUT: br_319 
* OUTPUT: bl_320 
* OUTPUT: br_320 
* OUTPUT: bl_321 
* OUTPUT: br_321 
* OUTPUT: bl_322 
* OUTPUT: br_322 
* OUTPUT: bl_323 
* OUTPUT: br_323 
* OUTPUT: bl_324 
* OUTPUT: br_324 
* OUTPUT: bl_325 
* OUTPUT: br_325 
* OUTPUT: bl_326 
* OUTPUT: br_326 
* OUTPUT: bl_327 
* OUTPUT: br_327 
* OUTPUT: bl_328 
* OUTPUT: br_328 
* OUTPUT: bl_329 
* OUTPUT: br_329 
* OUTPUT: bl_330 
* OUTPUT: br_330 
* OUTPUT: bl_331 
* OUTPUT: br_331 
* OUTPUT: bl_332 
* OUTPUT: br_332 
* OUTPUT: bl_333 
* OUTPUT: br_333 
* OUTPUT: bl_334 
* OUTPUT: br_334 
* OUTPUT: bl_335 
* OUTPUT: br_335 
* OUTPUT: bl_336 
* OUTPUT: br_336 
* OUTPUT: bl_337 
* OUTPUT: br_337 
* OUTPUT: bl_338 
* OUTPUT: br_338 
* OUTPUT: bl_339 
* OUTPUT: br_339 
* OUTPUT: bl_340 
* OUTPUT: br_340 
* OUTPUT: bl_341 
* OUTPUT: br_341 
* OUTPUT: bl_342 
* OUTPUT: br_342 
* OUTPUT: bl_343 
* OUTPUT: br_343 
* OUTPUT: bl_344 
* OUTPUT: br_344 
* OUTPUT: bl_345 
* OUTPUT: br_345 
* OUTPUT: bl_346 
* OUTPUT: br_346 
* OUTPUT: bl_347 
* OUTPUT: br_347 
* OUTPUT: bl_348 
* OUTPUT: br_348 
* OUTPUT: bl_349 
* OUTPUT: br_349 
* OUTPUT: bl_350 
* OUTPUT: br_350 
* OUTPUT: bl_351 
* OUTPUT: br_351 
* OUTPUT: bl_352 
* OUTPUT: br_352 
* OUTPUT: bl_353 
* OUTPUT: br_353 
* OUTPUT: bl_354 
* OUTPUT: br_354 
* OUTPUT: bl_355 
* OUTPUT: br_355 
* OUTPUT: bl_356 
* OUTPUT: br_356 
* OUTPUT: bl_357 
* OUTPUT: br_357 
* OUTPUT: bl_358 
* OUTPUT: br_358 
* OUTPUT: bl_359 
* OUTPUT: br_359 
* OUTPUT: bl_360 
* OUTPUT: br_360 
* OUTPUT: bl_361 
* OUTPUT: br_361 
* OUTPUT: bl_362 
* OUTPUT: br_362 
* OUTPUT: bl_363 
* OUTPUT: br_363 
* OUTPUT: bl_364 
* OUTPUT: br_364 
* OUTPUT: bl_365 
* OUTPUT: br_365 
* OUTPUT: bl_366 
* OUTPUT: br_366 
* OUTPUT: bl_367 
* OUTPUT: br_367 
* OUTPUT: bl_368 
* OUTPUT: br_368 
* OUTPUT: bl_369 
* OUTPUT: br_369 
* OUTPUT: bl_370 
* OUTPUT: br_370 
* OUTPUT: bl_371 
* OUTPUT: br_371 
* OUTPUT: bl_372 
* OUTPUT: br_372 
* OUTPUT: bl_373 
* OUTPUT: br_373 
* OUTPUT: bl_374 
* OUTPUT: br_374 
* OUTPUT: bl_375 
* OUTPUT: br_375 
* OUTPUT: bl_376 
* OUTPUT: br_376 
* OUTPUT: bl_377 
* OUTPUT: br_377 
* OUTPUT: bl_378 
* OUTPUT: br_378 
* OUTPUT: bl_379 
* OUTPUT: br_379 
* OUTPUT: bl_380 
* OUTPUT: br_380 
* OUTPUT: bl_381 
* OUTPUT: br_381 
* OUTPUT: bl_382 
* OUTPUT: br_382 
* OUTPUT: bl_383 
* OUTPUT: br_383 
* OUTPUT: bl_384 
* OUTPUT: br_384 
* OUTPUT: bl_385 
* OUTPUT: br_385 
* OUTPUT: bl_386 
* OUTPUT: br_386 
* OUTPUT: bl_387 
* OUTPUT: br_387 
* OUTPUT: bl_388 
* OUTPUT: br_388 
* OUTPUT: bl_389 
* OUTPUT: br_389 
* OUTPUT: bl_390 
* OUTPUT: br_390 
* OUTPUT: bl_391 
* OUTPUT: br_391 
* OUTPUT: bl_392 
* OUTPUT: br_392 
* OUTPUT: bl_393 
* OUTPUT: br_393 
* OUTPUT: bl_394 
* OUTPUT: br_394 
* OUTPUT: bl_395 
* OUTPUT: br_395 
* OUTPUT: bl_396 
* OUTPUT: br_396 
* OUTPUT: bl_397 
* OUTPUT: br_397 
* OUTPUT: bl_398 
* OUTPUT: br_398 
* OUTPUT: bl_399 
* OUTPUT: br_399 
* OUTPUT: bl_400 
* OUTPUT: br_400 
* OUTPUT: bl_401 
* OUTPUT: br_401 
* OUTPUT: bl_402 
* OUTPUT: br_402 
* OUTPUT: bl_403 
* OUTPUT: br_403 
* OUTPUT: bl_404 
* OUTPUT: br_404 
* OUTPUT: bl_405 
* OUTPUT: br_405 
* OUTPUT: bl_406 
* OUTPUT: br_406 
* OUTPUT: bl_407 
* OUTPUT: br_407 
* OUTPUT: bl_408 
* OUTPUT: br_408 
* OUTPUT: bl_409 
* OUTPUT: br_409 
* OUTPUT: bl_410 
* OUTPUT: br_410 
* OUTPUT: bl_411 
* OUTPUT: br_411 
* OUTPUT: bl_412 
* OUTPUT: br_412 
* OUTPUT: bl_413 
* OUTPUT: br_413 
* OUTPUT: bl_414 
* OUTPUT: br_414 
* OUTPUT: bl_415 
* OUTPUT: br_415 
* OUTPUT: bl_416 
* OUTPUT: br_416 
* OUTPUT: bl_417 
* OUTPUT: br_417 
* OUTPUT: bl_418 
* OUTPUT: br_418 
* OUTPUT: bl_419 
* OUTPUT: br_419 
* OUTPUT: bl_420 
* OUTPUT: br_420 
* OUTPUT: bl_421 
* OUTPUT: br_421 
* OUTPUT: bl_422 
* OUTPUT: br_422 
* OUTPUT: bl_423 
* OUTPUT: br_423 
* OUTPUT: bl_424 
* OUTPUT: br_424 
* OUTPUT: bl_425 
* OUTPUT: br_425 
* OUTPUT: bl_426 
* OUTPUT: br_426 
* OUTPUT: bl_427 
* OUTPUT: br_427 
* OUTPUT: bl_428 
* OUTPUT: br_428 
* OUTPUT: bl_429 
* OUTPUT: br_429 
* OUTPUT: bl_430 
* OUTPUT: br_430 
* OUTPUT: bl_431 
* OUTPUT: br_431 
* OUTPUT: bl_432 
* OUTPUT: br_432 
* OUTPUT: bl_433 
* OUTPUT: br_433 
* OUTPUT: bl_434 
* OUTPUT: br_434 
* OUTPUT: bl_435 
* OUTPUT: br_435 
* OUTPUT: bl_436 
* OUTPUT: br_436 
* OUTPUT: bl_437 
* OUTPUT: br_437 
* OUTPUT: bl_438 
* OUTPUT: br_438 
* OUTPUT: bl_439 
* OUTPUT: br_439 
* OUTPUT: bl_440 
* OUTPUT: br_440 
* OUTPUT: bl_441 
* OUTPUT: br_441 
* OUTPUT: bl_442 
* OUTPUT: br_442 
* OUTPUT: bl_443 
* OUTPUT: br_443 
* OUTPUT: bl_444 
* OUTPUT: br_444 
* OUTPUT: bl_445 
* OUTPUT: br_445 
* OUTPUT: bl_446 
* OUTPUT: br_446 
* OUTPUT: bl_447 
* OUTPUT: br_447 
* OUTPUT: bl_448 
* OUTPUT: br_448 
* OUTPUT: bl_449 
* OUTPUT: br_449 
* OUTPUT: bl_450 
* OUTPUT: br_450 
* OUTPUT: bl_451 
* OUTPUT: br_451 
* OUTPUT: bl_452 
* OUTPUT: br_452 
* OUTPUT: bl_453 
* OUTPUT: br_453 
* OUTPUT: bl_454 
* OUTPUT: br_454 
* OUTPUT: bl_455 
* OUTPUT: br_455 
* OUTPUT: bl_456 
* OUTPUT: br_456 
* OUTPUT: bl_457 
* OUTPUT: br_457 
* OUTPUT: bl_458 
* OUTPUT: br_458 
* OUTPUT: bl_459 
* OUTPUT: br_459 
* OUTPUT: bl_460 
* OUTPUT: br_460 
* OUTPUT: bl_461 
* OUTPUT: br_461 
* OUTPUT: bl_462 
* OUTPUT: br_462 
* OUTPUT: bl_463 
* OUTPUT: br_463 
* OUTPUT: bl_464 
* OUTPUT: br_464 
* OUTPUT: bl_465 
* OUTPUT: br_465 
* OUTPUT: bl_466 
* OUTPUT: br_466 
* OUTPUT: bl_467 
* OUTPUT: br_467 
* OUTPUT: bl_468 
* OUTPUT: br_468 
* OUTPUT: bl_469 
* OUTPUT: br_469 
* OUTPUT: bl_470 
* OUTPUT: br_470 
* OUTPUT: bl_471 
* OUTPUT: br_471 
* OUTPUT: bl_472 
* OUTPUT: br_472 
* OUTPUT: bl_473 
* OUTPUT: br_473 
* OUTPUT: bl_474 
* OUTPUT: br_474 
* OUTPUT: bl_475 
* OUTPUT: br_475 
* OUTPUT: bl_476 
* OUTPUT: br_476 
* OUTPUT: bl_477 
* OUTPUT: br_477 
* OUTPUT: bl_478 
* OUTPUT: br_478 
* OUTPUT: bl_479 
* OUTPUT: br_479 
* OUTPUT: bl_480 
* OUTPUT: br_480 
* OUTPUT: bl_481 
* OUTPUT: br_481 
* OUTPUT: bl_482 
* OUTPUT: br_482 
* OUTPUT: bl_483 
* OUTPUT: br_483 
* OUTPUT: bl_484 
* OUTPUT: br_484 
* OUTPUT: bl_485 
* OUTPUT: br_485 
* OUTPUT: bl_486 
* OUTPUT: br_486 
* OUTPUT: bl_487 
* OUTPUT: br_487 
* OUTPUT: bl_488 
* OUTPUT: br_488 
* OUTPUT: bl_489 
* OUTPUT: br_489 
* OUTPUT: bl_490 
* OUTPUT: br_490 
* OUTPUT: bl_491 
* OUTPUT: br_491 
* OUTPUT: bl_492 
* OUTPUT: br_492 
* OUTPUT: bl_493 
* OUTPUT: br_493 
* OUTPUT: bl_494 
* OUTPUT: br_494 
* OUTPUT: bl_495 
* OUTPUT: br_495 
* OUTPUT: bl_496 
* OUTPUT: br_496 
* OUTPUT: bl_497 
* OUTPUT: br_497 
* OUTPUT: bl_498 
* OUTPUT: br_498 
* OUTPUT: bl_499 
* OUTPUT: br_499 
* OUTPUT: bl_500 
* OUTPUT: br_500 
* OUTPUT: bl_501 
* OUTPUT: br_501 
* OUTPUT: bl_502 
* OUTPUT: br_502 
* OUTPUT: bl_503 
* OUTPUT: br_503 
* OUTPUT: bl_504 
* OUTPUT: br_504 
* OUTPUT: bl_505 
* OUTPUT: br_505 
* OUTPUT: bl_506 
* OUTPUT: br_506 
* OUTPUT: bl_507 
* OUTPUT: br_507 
* OUTPUT: bl_508 
* OUTPUT: br_508 
* OUTPUT: bl_509 
* OUTPUT: br_509 
* OUTPUT: bl_510 
* OUTPUT: br_510 
* OUTPUT: bl_511 
* OUTPUT: br_511 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* word_size 512
Xwrite_driver0
+ data_0 bl_0 br_0 en vdd gnd
+ write_driver
Xwrite_driver1
+ data_1 bl_1 br_1 en vdd gnd
+ write_driver
Xwrite_driver2
+ data_2 bl_2 br_2 en vdd gnd
+ write_driver
Xwrite_driver3
+ data_3 bl_3 br_3 en vdd gnd
+ write_driver
Xwrite_driver4
+ data_4 bl_4 br_4 en vdd gnd
+ write_driver
Xwrite_driver5
+ data_5 bl_5 br_5 en vdd gnd
+ write_driver
Xwrite_driver6
+ data_6 bl_6 br_6 en vdd gnd
+ write_driver
Xwrite_driver7
+ data_7 bl_7 br_7 en vdd gnd
+ write_driver
Xwrite_driver8
+ data_8 bl_8 br_8 en vdd gnd
+ write_driver
Xwrite_driver9
+ data_9 bl_9 br_9 en vdd gnd
+ write_driver
Xwrite_driver10
+ data_10 bl_10 br_10 en vdd gnd
+ write_driver
Xwrite_driver11
+ data_11 bl_11 br_11 en vdd gnd
+ write_driver
Xwrite_driver12
+ data_12 bl_12 br_12 en vdd gnd
+ write_driver
Xwrite_driver13
+ data_13 bl_13 br_13 en vdd gnd
+ write_driver
Xwrite_driver14
+ data_14 bl_14 br_14 en vdd gnd
+ write_driver
Xwrite_driver15
+ data_15 bl_15 br_15 en vdd gnd
+ write_driver
Xwrite_driver16
+ data_16 bl_16 br_16 en vdd gnd
+ write_driver
Xwrite_driver17
+ data_17 bl_17 br_17 en vdd gnd
+ write_driver
Xwrite_driver18
+ data_18 bl_18 br_18 en vdd gnd
+ write_driver
Xwrite_driver19
+ data_19 bl_19 br_19 en vdd gnd
+ write_driver
Xwrite_driver20
+ data_20 bl_20 br_20 en vdd gnd
+ write_driver
Xwrite_driver21
+ data_21 bl_21 br_21 en vdd gnd
+ write_driver
Xwrite_driver22
+ data_22 bl_22 br_22 en vdd gnd
+ write_driver
Xwrite_driver23
+ data_23 bl_23 br_23 en vdd gnd
+ write_driver
Xwrite_driver24
+ data_24 bl_24 br_24 en vdd gnd
+ write_driver
Xwrite_driver25
+ data_25 bl_25 br_25 en vdd gnd
+ write_driver
Xwrite_driver26
+ data_26 bl_26 br_26 en vdd gnd
+ write_driver
Xwrite_driver27
+ data_27 bl_27 br_27 en vdd gnd
+ write_driver
Xwrite_driver28
+ data_28 bl_28 br_28 en vdd gnd
+ write_driver
Xwrite_driver29
+ data_29 bl_29 br_29 en vdd gnd
+ write_driver
Xwrite_driver30
+ data_30 bl_30 br_30 en vdd gnd
+ write_driver
Xwrite_driver31
+ data_31 bl_31 br_31 en vdd gnd
+ write_driver
Xwrite_driver32
+ data_32 bl_32 br_32 en vdd gnd
+ write_driver
Xwrite_driver33
+ data_33 bl_33 br_33 en vdd gnd
+ write_driver
Xwrite_driver34
+ data_34 bl_34 br_34 en vdd gnd
+ write_driver
Xwrite_driver35
+ data_35 bl_35 br_35 en vdd gnd
+ write_driver
Xwrite_driver36
+ data_36 bl_36 br_36 en vdd gnd
+ write_driver
Xwrite_driver37
+ data_37 bl_37 br_37 en vdd gnd
+ write_driver
Xwrite_driver38
+ data_38 bl_38 br_38 en vdd gnd
+ write_driver
Xwrite_driver39
+ data_39 bl_39 br_39 en vdd gnd
+ write_driver
Xwrite_driver40
+ data_40 bl_40 br_40 en vdd gnd
+ write_driver
Xwrite_driver41
+ data_41 bl_41 br_41 en vdd gnd
+ write_driver
Xwrite_driver42
+ data_42 bl_42 br_42 en vdd gnd
+ write_driver
Xwrite_driver43
+ data_43 bl_43 br_43 en vdd gnd
+ write_driver
Xwrite_driver44
+ data_44 bl_44 br_44 en vdd gnd
+ write_driver
Xwrite_driver45
+ data_45 bl_45 br_45 en vdd gnd
+ write_driver
Xwrite_driver46
+ data_46 bl_46 br_46 en vdd gnd
+ write_driver
Xwrite_driver47
+ data_47 bl_47 br_47 en vdd gnd
+ write_driver
Xwrite_driver48
+ data_48 bl_48 br_48 en vdd gnd
+ write_driver
Xwrite_driver49
+ data_49 bl_49 br_49 en vdd gnd
+ write_driver
Xwrite_driver50
+ data_50 bl_50 br_50 en vdd gnd
+ write_driver
Xwrite_driver51
+ data_51 bl_51 br_51 en vdd gnd
+ write_driver
Xwrite_driver52
+ data_52 bl_52 br_52 en vdd gnd
+ write_driver
Xwrite_driver53
+ data_53 bl_53 br_53 en vdd gnd
+ write_driver
Xwrite_driver54
+ data_54 bl_54 br_54 en vdd gnd
+ write_driver
Xwrite_driver55
+ data_55 bl_55 br_55 en vdd gnd
+ write_driver
Xwrite_driver56
+ data_56 bl_56 br_56 en vdd gnd
+ write_driver
Xwrite_driver57
+ data_57 bl_57 br_57 en vdd gnd
+ write_driver
Xwrite_driver58
+ data_58 bl_58 br_58 en vdd gnd
+ write_driver
Xwrite_driver59
+ data_59 bl_59 br_59 en vdd gnd
+ write_driver
Xwrite_driver60
+ data_60 bl_60 br_60 en vdd gnd
+ write_driver
Xwrite_driver61
+ data_61 bl_61 br_61 en vdd gnd
+ write_driver
Xwrite_driver62
+ data_62 bl_62 br_62 en vdd gnd
+ write_driver
Xwrite_driver63
+ data_63 bl_63 br_63 en vdd gnd
+ write_driver
Xwrite_driver64
+ data_64 bl_64 br_64 en vdd gnd
+ write_driver
Xwrite_driver65
+ data_65 bl_65 br_65 en vdd gnd
+ write_driver
Xwrite_driver66
+ data_66 bl_66 br_66 en vdd gnd
+ write_driver
Xwrite_driver67
+ data_67 bl_67 br_67 en vdd gnd
+ write_driver
Xwrite_driver68
+ data_68 bl_68 br_68 en vdd gnd
+ write_driver
Xwrite_driver69
+ data_69 bl_69 br_69 en vdd gnd
+ write_driver
Xwrite_driver70
+ data_70 bl_70 br_70 en vdd gnd
+ write_driver
Xwrite_driver71
+ data_71 bl_71 br_71 en vdd gnd
+ write_driver
Xwrite_driver72
+ data_72 bl_72 br_72 en vdd gnd
+ write_driver
Xwrite_driver73
+ data_73 bl_73 br_73 en vdd gnd
+ write_driver
Xwrite_driver74
+ data_74 bl_74 br_74 en vdd gnd
+ write_driver
Xwrite_driver75
+ data_75 bl_75 br_75 en vdd gnd
+ write_driver
Xwrite_driver76
+ data_76 bl_76 br_76 en vdd gnd
+ write_driver
Xwrite_driver77
+ data_77 bl_77 br_77 en vdd gnd
+ write_driver
Xwrite_driver78
+ data_78 bl_78 br_78 en vdd gnd
+ write_driver
Xwrite_driver79
+ data_79 bl_79 br_79 en vdd gnd
+ write_driver
Xwrite_driver80
+ data_80 bl_80 br_80 en vdd gnd
+ write_driver
Xwrite_driver81
+ data_81 bl_81 br_81 en vdd gnd
+ write_driver
Xwrite_driver82
+ data_82 bl_82 br_82 en vdd gnd
+ write_driver
Xwrite_driver83
+ data_83 bl_83 br_83 en vdd gnd
+ write_driver
Xwrite_driver84
+ data_84 bl_84 br_84 en vdd gnd
+ write_driver
Xwrite_driver85
+ data_85 bl_85 br_85 en vdd gnd
+ write_driver
Xwrite_driver86
+ data_86 bl_86 br_86 en vdd gnd
+ write_driver
Xwrite_driver87
+ data_87 bl_87 br_87 en vdd gnd
+ write_driver
Xwrite_driver88
+ data_88 bl_88 br_88 en vdd gnd
+ write_driver
Xwrite_driver89
+ data_89 bl_89 br_89 en vdd gnd
+ write_driver
Xwrite_driver90
+ data_90 bl_90 br_90 en vdd gnd
+ write_driver
Xwrite_driver91
+ data_91 bl_91 br_91 en vdd gnd
+ write_driver
Xwrite_driver92
+ data_92 bl_92 br_92 en vdd gnd
+ write_driver
Xwrite_driver93
+ data_93 bl_93 br_93 en vdd gnd
+ write_driver
Xwrite_driver94
+ data_94 bl_94 br_94 en vdd gnd
+ write_driver
Xwrite_driver95
+ data_95 bl_95 br_95 en vdd gnd
+ write_driver
Xwrite_driver96
+ data_96 bl_96 br_96 en vdd gnd
+ write_driver
Xwrite_driver97
+ data_97 bl_97 br_97 en vdd gnd
+ write_driver
Xwrite_driver98
+ data_98 bl_98 br_98 en vdd gnd
+ write_driver
Xwrite_driver99
+ data_99 bl_99 br_99 en vdd gnd
+ write_driver
Xwrite_driver100
+ data_100 bl_100 br_100 en vdd gnd
+ write_driver
Xwrite_driver101
+ data_101 bl_101 br_101 en vdd gnd
+ write_driver
Xwrite_driver102
+ data_102 bl_102 br_102 en vdd gnd
+ write_driver
Xwrite_driver103
+ data_103 bl_103 br_103 en vdd gnd
+ write_driver
Xwrite_driver104
+ data_104 bl_104 br_104 en vdd gnd
+ write_driver
Xwrite_driver105
+ data_105 bl_105 br_105 en vdd gnd
+ write_driver
Xwrite_driver106
+ data_106 bl_106 br_106 en vdd gnd
+ write_driver
Xwrite_driver107
+ data_107 bl_107 br_107 en vdd gnd
+ write_driver
Xwrite_driver108
+ data_108 bl_108 br_108 en vdd gnd
+ write_driver
Xwrite_driver109
+ data_109 bl_109 br_109 en vdd gnd
+ write_driver
Xwrite_driver110
+ data_110 bl_110 br_110 en vdd gnd
+ write_driver
Xwrite_driver111
+ data_111 bl_111 br_111 en vdd gnd
+ write_driver
Xwrite_driver112
+ data_112 bl_112 br_112 en vdd gnd
+ write_driver
Xwrite_driver113
+ data_113 bl_113 br_113 en vdd gnd
+ write_driver
Xwrite_driver114
+ data_114 bl_114 br_114 en vdd gnd
+ write_driver
Xwrite_driver115
+ data_115 bl_115 br_115 en vdd gnd
+ write_driver
Xwrite_driver116
+ data_116 bl_116 br_116 en vdd gnd
+ write_driver
Xwrite_driver117
+ data_117 bl_117 br_117 en vdd gnd
+ write_driver
Xwrite_driver118
+ data_118 bl_118 br_118 en vdd gnd
+ write_driver
Xwrite_driver119
+ data_119 bl_119 br_119 en vdd gnd
+ write_driver
Xwrite_driver120
+ data_120 bl_120 br_120 en vdd gnd
+ write_driver
Xwrite_driver121
+ data_121 bl_121 br_121 en vdd gnd
+ write_driver
Xwrite_driver122
+ data_122 bl_122 br_122 en vdd gnd
+ write_driver
Xwrite_driver123
+ data_123 bl_123 br_123 en vdd gnd
+ write_driver
Xwrite_driver124
+ data_124 bl_124 br_124 en vdd gnd
+ write_driver
Xwrite_driver125
+ data_125 bl_125 br_125 en vdd gnd
+ write_driver
Xwrite_driver126
+ data_126 bl_126 br_126 en vdd gnd
+ write_driver
Xwrite_driver127
+ data_127 bl_127 br_127 en vdd gnd
+ write_driver
Xwrite_driver128
+ data_128 bl_128 br_128 en vdd gnd
+ write_driver
Xwrite_driver129
+ data_129 bl_129 br_129 en vdd gnd
+ write_driver
Xwrite_driver130
+ data_130 bl_130 br_130 en vdd gnd
+ write_driver
Xwrite_driver131
+ data_131 bl_131 br_131 en vdd gnd
+ write_driver
Xwrite_driver132
+ data_132 bl_132 br_132 en vdd gnd
+ write_driver
Xwrite_driver133
+ data_133 bl_133 br_133 en vdd gnd
+ write_driver
Xwrite_driver134
+ data_134 bl_134 br_134 en vdd gnd
+ write_driver
Xwrite_driver135
+ data_135 bl_135 br_135 en vdd gnd
+ write_driver
Xwrite_driver136
+ data_136 bl_136 br_136 en vdd gnd
+ write_driver
Xwrite_driver137
+ data_137 bl_137 br_137 en vdd gnd
+ write_driver
Xwrite_driver138
+ data_138 bl_138 br_138 en vdd gnd
+ write_driver
Xwrite_driver139
+ data_139 bl_139 br_139 en vdd gnd
+ write_driver
Xwrite_driver140
+ data_140 bl_140 br_140 en vdd gnd
+ write_driver
Xwrite_driver141
+ data_141 bl_141 br_141 en vdd gnd
+ write_driver
Xwrite_driver142
+ data_142 bl_142 br_142 en vdd gnd
+ write_driver
Xwrite_driver143
+ data_143 bl_143 br_143 en vdd gnd
+ write_driver
Xwrite_driver144
+ data_144 bl_144 br_144 en vdd gnd
+ write_driver
Xwrite_driver145
+ data_145 bl_145 br_145 en vdd gnd
+ write_driver
Xwrite_driver146
+ data_146 bl_146 br_146 en vdd gnd
+ write_driver
Xwrite_driver147
+ data_147 bl_147 br_147 en vdd gnd
+ write_driver
Xwrite_driver148
+ data_148 bl_148 br_148 en vdd gnd
+ write_driver
Xwrite_driver149
+ data_149 bl_149 br_149 en vdd gnd
+ write_driver
Xwrite_driver150
+ data_150 bl_150 br_150 en vdd gnd
+ write_driver
Xwrite_driver151
+ data_151 bl_151 br_151 en vdd gnd
+ write_driver
Xwrite_driver152
+ data_152 bl_152 br_152 en vdd gnd
+ write_driver
Xwrite_driver153
+ data_153 bl_153 br_153 en vdd gnd
+ write_driver
Xwrite_driver154
+ data_154 bl_154 br_154 en vdd gnd
+ write_driver
Xwrite_driver155
+ data_155 bl_155 br_155 en vdd gnd
+ write_driver
Xwrite_driver156
+ data_156 bl_156 br_156 en vdd gnd
+ write_driver
Xwrite_driver157
+ data_157 bl_157 br_157 en vdd gnd
+ write_driver
Xwrite_driver158
+ data_158 bl_158 br_158 en vdd gnd
+ write_driver
Xwrite_driver159
+ data_159 bl_159 br_159 en vdd gnd
+ write_driver
Xwrite_driver160
+ data_160 bl_160 br_160 en vdd gnd
+ write_driver
Xwrite_driver161
+ data_161 bl_161 br_161 en vdd gnd
+ write_driver
Xwrite_driver162
+ data_162 bl_162 br_162 en vdd gnd
+ write_driver
Xwrite_driver163
+ data_163 bl_163 br_163 en vdd gnd
+ write_driver
Xwrite_driver164
+ data_164 bl_164 br_164 en vdd gnd
+ write_driver
Xwrite_driver165
+ data_165 bl_165 br_165 en vdd gnd
+ write_driver
Xwrite_driver166
+ data_166 bl_166 br_166 en vdd gnd
+ write_driver
Xwrite_driver167
+ data_167 bl_167 br_167 en vdd gnd
+ write_driver
Xwrite_driver168
+ data_168 bl_168 br_168 en vdd gnd
+ write_driver
Xwrite_driver169
+ data_169 bl_169 br_169 en vdd gnd
+ write_driver
Xwrite_driver170
+ data_170 bl_170 br_170 en vdd gnd
+ write_driver
Xwrite_driver171
+ data_171 bl_171 br_171 en vdd gnd
+ write_driver
Xwrite_driver172
+ data_172 bl_172 br_172 en vdd gnd
+ write_driver
Xwrite_driver173
+ data_173 bl_173 br_173 en vdd gnd
+ write_driver
Xwrite_driver174
+ data_174 bl_174 br_174 en vdd gnd
+ write_driver
Xwrite_driver175
+ data_175 bl_175 br_175 en vdd gnd
+ write_driver
Xwrite_driver176
+ data_176 bl_176 br_176 en vdd gnd
+ write_driver
Xwrite_driver177
+ data_177 bl_177 br_177 en vdd gnd
+ write_driver
Xwrite_driver178
+ data_178 bl_178 br_178 en vdd gnd
+ write_driver
Xwrite_driver179
+ data_179 bl_179 br_179 en vdd gnd
+ write_driver
Xwrite_driver180
+ data_180 bl_180 br_180 en vdd gnd
+ write_driver
Xwrite_driver181
+ data_181 bl_181 br_181 en vdd gnd
+ write_driver
Xwrite_driver182
+ data_182 bl_182 br_182 en vdd gnd
+ write_driver
Xwrite_driver183
+ data_183 bl_183 br_183 en vdd gnd
+ write_driver
Xwrite_driver184
+ data_184 bl_184 br_184 en vdd gnd
+ write_driver
Xwrite_driver185
+ data_185 bl_185 br_185 en vdd gnd
+ write_driver
Xwrite_driver186
+ data_186 bl_186 br_186 en vdd gnd
+ write_driver
Xwrite_driver187
+ data_187 bl_187 br_187 en vdd gnd
+ write_driver
Xwrite_driver188
+ data_188 bl_188 br_188 en vdd gnd
+ write_driver
Xwrite_driver189
+ data_189 bl_189 br_189 en vdd gnd
+ write_driver
Xwrite_driver190
+ data_190 bl_190 br_190 en vdd gnd
+ write_driver
Xwrite_driver191
+ data_191 bl_191 br_191 en vdd gnd
+ write_driver
Xwrite_driver192
+ data_192 bl_192 br_192 en vdd gnd
+ write_driver
Xwrite_driver193
+ data_193 bl_193 br_193 en vdd gnd
+ write_driver
Xwrite_driver194
+ data_194 bl_194 br_194 en vdd gnd
+ write_driver
Xwrite_driver195
+ data_195 bl_195 br_195 en vdd gnd
+ write_driver
Xwrite_driver196
+ data_196 bl_196 br_196 en vdd gnd
+ write_driver
Xwrite_driver197
+ data_197 bl_197 br_197 en vdd gnd
+ write_driver
Xwrite_driver198
+ data_198 bl_198 br_198 en vdd gnd
+ write_driver
Xwrite_driver199
+ data_199 bl_199 br_199 en vdd gnd
+ write_driver
Xwrite_driver200
+ data_200 bl_200 br_200 en vdd gnd
+ write_driver
Xwrite_driver201
+ data_201 bl_201 br_201 en vdd gnd
+ write_driver
Xwrite_driver202
+ data_202 bl_202 br_202 en vdd gnd
+ write_driver
Xwrite_driver203
+ data_203 bl_203 br_203 en vdd gnd
+ write_driver
Xwrite_driver204
+ data_204 bl_204 br_204 en vdd gnd
+ write_driver
Xwrite_driver205
+ data_205 bl_205 br_205 en vdd gnd
+ write_driver
Xwrite_driver206
+ data_206 bl_206 br_206 en vdd gnd
+ write_driver
Xwrite_driver207
+ data_207 bl_207 br_207 en vdd gnd
+ write_driver
Xwrite_driver208
+ data_208 bl_208 br_208 en vdd gnd
+ write_driver
Xwrite_driver209
+ data_209 bl_209 br_209 en vdd gnd
+ write_driver
Xwrite_driver210
+ data_210 bl_210 br_210 en vdd gnd
+ write_driver
Xwrite_driver211
+ data_211 bl_211 br_211 en vdd gnd
+ write_driver
Xwrite_driver212
+ data_212 bl_212 br_212 en vdd gnd
+ write_driver
Xwrite_driver213
+ data_213 bl_213 br_213 en vdd gnd
+ write_driver
Xwrite_driver214
+ data_214 bl_214 br_214 en vdd gnd
+ write_driver
Xwrite_driver215
+ data_215 bl_215 br_215 en vdd gnd
+ write_driver
Xwrite_driver216
+ data_216 bl_216 br_216 en vdd gnd
+ write_driver
Xwrite_driver217
+ data_217 bl_217 br_217 en vdd gnd
+ write_driver
Xwrite_driver218
+ data_218 bl_218 br_218 en vdd gnd
+ write_driver
Xwrite_driver219
+ data_219 bl_219 br_219 en vdd gnd
+ write_driver
Xwrite_driver220
+ data_220 bl_220 br_220 en vdd gnd
+ write_driver
Xwrite_driver221
+ data_221 bl_221 br_221 en vdd gnd
+ write_driver
Xwrite_driver222
+ data_222 bl_222 br_222 en vdd gnd
+ write_driver
Xwrite_driver223
+ data_223 bl_223 br_223 en vdd gnd
+ write_driver
Xwrite_driver224
+ data_224 bl_224 br_224 en vdd gnd
+ write_driver
Xwrite_driver225
+ data_225 bl_225 br_225 en vdd gnd
+ write_driver
Xwrite_driver226
+ data_226 bl_226 br_226 en vdd gnd
+ write_driver
Xwrite_driver227
+ data_227 bl_227 br_227 en vdd gnd
+ write_driver
Xwrite_driver228
+ data_228 bl_228 br_228 en vdd gnd
+ write_driver
Xwrite_driver229
+ data_229 bl_229 br_229 en vdd gnd
+ write_driver
Xwrite_driver230
+ data_230 bl_230 br_230 en vdd gnd
+ write_driver
Xwrite_driver231
+ data_231 bl_231 br_231 en vdd gnd
+ write_driver
Xwrite_driver232
+ data_232 bl_232 br_232 en vdd gnd
+ write_driver
Xwrite_driver233
+ data_233 bl_233 br_233 en vdd gnd
+ write_driver
Xwrite_driver234
+ data_234 bl_234 br_234 en vdd gnd
+ write_driver
Xwrite_driver235
+ data_235 bl_235 br_235 en vdd gnd
+ write_driver
Xwrite_driver236
+ data_236 bl_236 br_236 en vdd gnd
+ write_driver
Xwrite_driver237
+ data_237 bl_237 br_237 en vdd gnd
+ write_driver
Xwrite_driver238
+ data_238 bl_238 br_238 en vdd gnd
+ write_driver
Xwrite_driver239
+ data_239 bl_239 br_239 en vdd gnd
+ write_driver
Xwrite_driver240
+ data_240 bl_240 br_240 en vdd gnd
+ write_driver
Xwrite_driver241
+ data_241 bl_241 br_241 en vdd gnd
+ write_driver
Xwrite_driver242
+ data_242 bl_242 br_242 en vdd gnd
+ write_driver
Xwrite_driver243
+ data_243 bl_243 br_243 en vdd gnd
+ write_driver
Xwrite_driver244
+ data_244 bl_244 br_244 en vdd gnd
+ write_driver
Xwrite_driver245
+ data_245 bl_245 br_245 en vdd gnd
+ write_driver
Xwrite_driver246
+ data_246 bl_246 br_246 en vdd gnd
+ write_driver
Xwrite_driver247
+ data_247 bl_247 br_247 en vdd gnd
+ write_driver
Xwrite_driver248
+ data_248 bl_248 br_248 en vdd gnd
+ write_driver
Xwrite_driver249
+ data_249 bl_249 br_249 en vdd gnd
+ write_driver
Xwrite_driver250
+ data_250 bl_250 br_250 en vdd gnd
+ write_driver
Xwrite_driver251
+ data_251 bl_251 br_251 en vdd gnd
+ write_driver
Xwrite_driver252
+ data_252 bl_252 br_252 en vdd gnd
+ write_driver
Xwrite_driver253
+ data_253 bl_253 br_253 en vdd gnd
+ write_driver
Xwrite_driver254
+ data_254 bl_254 br_254 en vdd gnd
+ write_driver
Xwrite_driver255
+ data_255 bl_255 br_255 en vdd gnd
+ write_driver
Xwrite_driver256
+ data_256 bl_256 br_256 en vdd gnd
+ write_driver
Xwrite_driver257
+ data_257 bl_257 br_257 en vdd gnd
+ write_driver
Xwrite_driver258
+ data_258 bl_258 br_258 en vdd gnd
+ write_driver
Xwrite_driver259
+ data_259 bl_259 br_259 en vdd gnd
+ write_driver
Xwrite_driver260
+ data_260 bl_260 br_260 en vdd gnd
+ write_driver
Xwrite_driver261
+ data_261 bl_261 br_261 en vdd gnd
+ write_driver
Xwrite_driver262
+ data_262 bl_262 br_262 en vdd gnd
+ write_driver
Xwrite_driver263
+ data_263 bl_263 br_263 en vdd gnd
+ write_driver
Xwrite_driver264
+ data_264 bl_264 br_264 en vdd gnd
+ write_driver
Xwrite_driver265
+ data_265 bl_265 br_265 en vdd gnd
+ write_driver
Xwrite_driver266
+ data_266 bl_266 br_266 en vdd gnd
+ write_driver
Xwrite_driver267
+ data_267 bl_267 br_267 en vdd gnd
+ write_driver
Xwrite_driver268
+ data_268 bl_268 br_268 en vdd gnd
+ write_driver
Xwrite_driver269
+ data_269 bl_269 br_269 en vdd gnd
+ write_driver
Xwrite_driver270
+ data_270 bl_270 br_270 en vdd gnd
+ write_driver
Xwrite_driver271
+ data_271 bl_271 br_271 en vdd gnd
+ write_driver
Xwrite_driver272
+ data_272 bl_272 br_272 en vdd gnd
+ write_driver
Xwrite_driver273
+ data_273 bl_273 br_273 en vdd gnd
+ write_driver
Xwrite_driver274
+ data_274 bl_274 br_274 en vdd gnd
+ write_driver
Xwrite_driver275
+ data_275 bl_275 br_275 en vdd gnd
+ write_driver
Xwrite_driver276
+ data_276 bl_276 br_276 en vdd gnd
+ write_driver
Xwrite_driver277
+ data_277 bl_277 br_277 en vdd gnd
+ write_driver
Xwrite_driver278
+ data_278 bl_278 br_278 en vdd gnd
+ write_driver
Xwrite_driver279
+ data_279 bl_279 br_279 en vdd gnd
+ write_driver
Xwrite_driver280
+ data_280 bl_280 br_280 en vdd gnd
+ write_driver
Xwrite_driver281
+ data_281 bl_281 br_281 en vdd gnd
+ write_driver
Xwrite_driver282
+ data_282 bl_282 br_282 en vdd gnd
+ write_driver
Xwrite_driver283
+ data_283 bl_283 br_283 en vdd gnd
+ write_driver
Xwrite_driver284
+ data_284 bl_284 br_284 en vdd gnd
+ write_driver
Xwrite_driver285
+ data_285 bl_285 br_285 en vdd gnd
+ write_driver
Xwrite_driver286
+ data_286 bl_286 br_286 en vdd gnd
+ write_driver
Xwrite_driver287
+ data_287 bl_287 br_287 en vdd gnd
+ write_driver
Xwrite_driver288
+ data_288 bl_288 br_288 en vdd gnd
+ write_driver
Xwrite_driver289
+ data_289 bl_289 br_289 en vdd gnd
+ write_driver
Xwrite_driver290
+ data_290 bl_290 br_290 en vdd gnd
+ write_driver
Xwrite_driver291
+ data_291 bl_291 br_291 en vdd gnd
+ write_driver
Xwrite_driver292
+ data_292 bl_292 br_292 en vdd gnd
+ write_driver
Xwrite_driver293
+ data_293 bl_293 br_293 en vdd gnd
+ write_driver
Xwrite_driver294
+ data_294 bl_294 br_294 en vdd gnd
+ write_driver
Xwrite_driver295
+ data_295 bl_295 br_295 en vdd gnd
+ write_driver
Xwrite_driver296
+ data_296 bl_296 br_296 en vdd gnd
+ write_driver
Xwrite_driver297
+ data_297 bl_297 br_297 en vdd gnd
+ write_driver
Xwrite_driver298
+ data_298 bl_298 br_298 en vdd gnd
+ write_driver
Xwrite_driver299
+ data_299 bl_299 br_299 en vdd gnd
+ write_driver
Xwrite_driver300
+ data_300 bl_300 br_300 en vdd gnd
+ write_driver
Xwrite_driver301
+ data_301 bl_301 br_301 en vdd gnd
+ write_driver
Xwrite_driver302
+ data_302 bl_302 br_302 en vdd gnd
+ write_driver
Xwrite_driver303
+ data_303 bl_303 br_303 en vdd gnd
+ write_driver
Xwrite_driver304
+ data_304 bl_304 br_304 en vdd gnd
+ write_driver
Xwrite_driver305
+ data_305 bl_305 br_305 en vdd gnd
+ write_driver
Xwrite_driver306
+ data_306 bl_306 br_306 en vdd gnd
+ write_driver
Xwrite_driver307
+ data_307 bl_307 br_307 en vdd gnd
+ write_driver
Xwrite_driver308
+ data_308 bl_308 br_308 en vdd gnd
+ write_driver
Xwrite_driver309
+ data_309 bl_309 br_309 en vdd gnd
+ write_driver
Xwrite_driver310
+ data_310 bl_310 br_310 en vdd gnd
+ write_driver
Xwrite_driver311
+ data_311 bl_311 br_311 en vdd gnd
+ write_driver
Xwrite_driver312
+ data_312 bl_312 br_312 en vdd gnd
+ write_driver
Xwrite_driver313
+ data_313 bl_313 br_313 en vdd gnd
+ write_driver
Xwrite_driver314
+ data_314 bl_314 br_314 en vdd gnd
+ write_driver
Xwrite_driver315
+ data_315 bl_315 br_315 en vdd gnd
+ write_driver
Xwrite_driver316
+ data_316 bl_316 br_316 en vdd gnd
+ write_driver
Xwrite_driver317
+ data_317 bl_317 br_317 en vdd gnd
+ write_driver
Xwrite_driver318
+ data_318 bl_318 br_318 en vdd gnd
+ write_driver
Xwrite_driver319
+ data_319 bl_319 br_319 en vdd gnd
+ write_driver
Xwrite_driver320
+ data_320 bl_320 br_320 en vdd gnd
+ write_driver
Xwrite_driver321
+ data_321 bl_321 br_321 en vdd gnd
+ write_driver
Xwrite_driver322
+ data_322 bl_322 br_322 en vdd gnd
+ write_driver
Xwrite_driver323
+ data_323 bl_323 br_323 en vdd gnd
+ write_driver
Xwrite_driver324
+ data_324 bl_324 br_324 en vdd gnd
+ write_driver
Xwrite_driver325
+ data_325 bl_325 br_325 en vdd gnd
+ write_driver
Xwrite_driver326
+ data_326 bl_326 br_326 en vdd gnd
+ write_driver
Xwrite_driver327
+ data_327 bl_327 br_327 en vdd gnd
+ write_driver
Xwrite_driver328
+ data_328 bl_328 br_328 en vdd gnd
+ write_driver
Xwrite_driver329
+ data_329 bl_329 br_329 en vdd gnd
+ write_driver
Xwrite_driver330
+ data_330 bl_330 br_330 en vdd gnd
+ write_driver
Xwrite_driver331
+ data_331 bl_331 br_331 en vdd gnd
+ write_driver
Xwrite_driver332
+ data_332 bl_332 br_332 en vdd gnd
+ write_driver
Xwrite_driver333
+ data_333 bl_333 br_333 en vdd gnd
+ write_driver
Xwrite_driver334
+ data_334 bl_334 br_334 en vdd gnd
+ write_driver
Xwrite_driver335
+ data_335 bl_335 br_335 en vdd gnd
+ write_driver
Xwrite_driver336
+ data_336 bl_336 br_336 en vdd gnd
+ write_driver
Xwrite_driver337
+ data_337 bl_337 br_337 en vdd gnd
+ write_driver
Xwrite_driver338
+ data_338 bl_338 br_338 en vdd gnd
+ write_driver
Xwrite_driver339
+ data_339 bl_339 br_339 en vdd gnd
+ write_driver
Xwrite_driver340
+ data_340 bl_340 br_340 en vdd gnd
+ write_driver
Xwrite_driver341
+ data_341 bl_341 br_341 en vdd gnd
+ write_driver
Xwrite_driver342
+ data_342 bl_342 br_342 en vdd gnd
+ write_driver
Xwrite_driver343
+ data_343 bl_343 br_343 en vdd gnd
+ write_driver
Xwrite_driver344
+ data_344 bl_344 br_344 en vdd gnd
+ write_driver
Xwrite_driver345
+ data_345 bl_345 br_345 en vdd gnd
+ write_driver
Xwrite_driver346
+ data_346 bl_346 br_346 en vdd gnd
+ write_driver
Xwrite_driver347
+ data_347 bl_347 br_347 en vdd gnd
+ write_driver
Xwrite_driver348
+ data_348 bl_348 br_348 en vdd gnd
+ write_driver
Xwrite_driver349
+ data_349 bl_349 br_349 en vdd gnd
+ write_driver
Xwrite_driver350
+ data_350 bl_350 br_350 en vdd gnd
+ write_driver
Xwrite_driver351
+ data_351 bl_351 br_351 en vdd gnd
+ write_driver
Xwrite_driver352
+ data_352 bl_352 br_352 en vdd gnd
+ write_driver
Xwrite_driver353
+ data_353 bl_353 br_353 en vdd gnd
+ write_driver
Xwrite_driver354
+ data_354 bl_354 br_354 en vdd gnd
+ write_driver
Xwrite_driver355
+ data_355 bl_355 br_355 en vdd gnd
+ write_driver
Xwrite_driver356
+ data_356 bl_356 br_356 en vdd gnd
+ write_driver
Xwrite_driver357
+ data_357 bl_357 br_357 en vdd gnd
+ write_driver
Xwrite_driver358
+ data_358 bl_358 br_358 en vdd gnd
+ write_driver
Xwrite_driver359
+ data_359 bl_359 br_359 en vdd gnd
+ write_driver
Xwrite_driver360
+ data_360 bl_360 br_360 en vdd gnd
+ write_driver
Xwrite_driver361
+ data_361 bl_361 br_361 en vdd gnd
+ write_driver
Xwrite_driver362
+ data_362 bl_362 br_362 en vdd gnd
+ write_driver
Xwrite_driver363
+ data_363 bl_363 br_363 en vdd gnd
+ write_driver
Xwrite_driver364
+ data_364 bl_364 br_364 en vdd gnd
+ write_driver
Xwrite_driver365
+ data_365 bl_365 br_365 en vdd gnd
+ write_driver
Xwrite_driver366
+ data_366 bl_366 br_366 en vdd gnd
+ write_driver
Xwrite_driver367
+ data_367 bl_367 br_367 en vdd gnd
+ write_driver
Xwrite_driver368
+ data_368 bl_368 br_368 en vdd gnd
+ write_driver
Xwrite_driver369
+ data_369 bl_369 br_369 en vdd gnd
+ write_driver
Xwrite_driver370
+ data_370 bl_370 br_370 en vdd gnd
+ write_driver
Xwrite_driver371
+ data_371 bl_371 br_371 en vdd gnd
+ write_driver
Xwrite_driver372
+ data_372 bl_372 br_372 en vdd gnd
+ write_driver
Xwrite_driver373
+ data_373 bl_373 br_373 en vdd gnd
+ write_driver
Xwrite_driver374
+ data_374 bl_374 br_374 en vdd gnd
+ write_driver
Xwrite_driver375
+ data_375 bl_375 br_375 en vdd gnd
+ write_driver
Xwrite_driver376
+ data_376 bl_376 br_376 en vdd gnd
+ write_driver
Xwrite_driver377
+ data_377 bl_377 br_377 en vdd gnd
+ write_driver
Xwrite_driver378
+ data_378 bl_378 br_378 en vdd gnd
+ write_driver
Xwrite_driver379
+ data_379 bl_379 br_379 en vdd gnd
+ write_driver
Xwrite_driver380
+ data_380 bl_380 br_380 en vdd gnd
+ write_driver
Xwrite_driver381
+ data_381 bl_381 br_381 en vdd gnd
+ write_driver
Xwrite_driver382
+ data_382 bl_382 br_382 en vdd gnd
+ write_driver
Xwrite_driver383
+ data_383 bl_383 br_383 en vdd gnd
+ write_driver
Xwrite_driver384
+ data_384 bl_384 br_384 en vdd gnd
+ write_driver
Xwrite_driver385
+ data_385 bl_385 br_385 en vdd gnd
+ write_driver
Xwrite_driver386
+ data_386 bl_386 br_386 en vdd gnd
+ write_driver
Xwrite_driver387
+ data_387 bl_387 br_387 en vdd gnd
+ write_driver
Xwrite_driver388
+ data_388 bl_388 br_388 en vdd gnd
+ write_driver
Xwrite_driver389
+ data_389 bl_389 br_389 en vdd gnd
+ write_driver
Xwrite_driver390
+ data_390 bl_390 br_390 en vdd gnd
+ write_driver
Xwrite_driver391
+ data_391 bl_391 br_391 en vdd gnd
+ write_driver
Xwrite_driver392
+ data_392 bl_392 br_392 en vdd gnd
+ write_driver
Xwrite_driver393
+ data_393 bl_393 br_393 en vdd gnd
+ write_driver
Xwrite_driver394
+ data_394 bl_394 br_394 en vdd gnd
+ write_driver
Xwrite_driver395
+ data_395 bl_395 br_395 en vdd gnd
+ write_driver
Xwrite_driver396
+ data_396 bl_396 br_396 en vdd gnd
+ write_driver
Xwrite_driver397
+ data_397 bl_397 br_397 en vdd gnd
+ write_driver
Xwrite_driver398
+ data_398 bl_398 br_398 en vdd gnd
+ write_driver
Xwrite_driver399
+ data_399 bl_399 br_399 en vdd gnd
+ write_driver
Xwrite_driver400
+ data_400 bl_400 br_400 en vdd gnd
+ write_driver
Xwrite_driver401
+ data_401 bl_401 br_401 en vdd gnd
+ write_driver
Xwrite_driver402
+ data_402 bl_402 br_402 en vdd gnd
+ write_driver
Xwrite_driver403
+ data_403 bl_403 br_403 en vdd gnd
+ write_driver
Xwrite_driver404
+ data_404 bl_404 br_404 en vdd gnd
+ write_driver
Xwrite_driver405
+ data_405 bl_405 br_405 en vdd gnd
+ write_driver
Xwrite_driver406
+ data_406 bl_406 br_406 en vdd gnd
+ write_driver
Xwrite_driver407
+ data_407 bl_407 br_407 en vdd gnd
+ write_driver
Xwrite_driver408
+ data_408 bl_408 br_408 en vdd gnd
+ write_driver
Xwrite_driver409
+ data_409 bl_409 br_409 en vdd gnd
+ write_driver
Xwrite_driver410
+ data_410 bl_410 br_410 en vdd gnd
+ write_driver
Xwrite_driver411
+ data_411 bl_411 br_411 en vdd gnd
+ write_driver
Xwrite_driver412
+ data_412 bl_412 br_412 en vdd gnd
+ write_driver
Xwrite_driver413
+ data_413 bl_413 br_413 en vdd gnd
+ write_driver
Xwrite_driver414
+ data_414 bl_414 br_414 en vdd gnd
+ write_driver
Xwrite_driver415
+ data_415 bl_415 br_415 en vdd gnd
+ write_driver
Xwrite_driver416
+ data_416 bl_416 br_416 en vdd gnd
+ write_driver
Xwrite_driver417
+ data_417 bl_417 br_417 en vdd gnd
+ write_driver
Xwrite_driver418
+ data_418 bl_418 br_418 en vdd gnd
+ write_driver
Xwrite_driver419
+ data_419 bl_419 br_419 en vdd gnd
+ write_driver
Xwrite_driver420
+ data_420 bl_420 br_420 en vdd gnd
+ write_driver
Xwrite_driver421
+ data_421 bl_421 br_421 en vdd gnd
+ write_driver
Xwrite_driver422
+ data_422 bl_422 br_422 en vdd gnd
+ write_driver
Xwrite_driver423
+ data_423 bl_423 br_423 en vdd gnd
+ write_driver
Xwrite_driver424
+ data_424 bl_424 br_424 en vdd gnd
+ write_driver
Xwrite_driver425
+ data_425 bl_425 br_425 en vdd gnd
+ write_driver
Xwrite_driver426
+ data_426 bl_426 br_426 en vdd gnd
+ write_driver
Xwrite_driver427
+ data_427 bl_427 br_427 en vdd gnd
+ write_driver
Xwrite_driver428
+ data_428 bl_428 br_428 en vdd gnd
+ write_driver
Xwrite_driver429
+ data_429 bl_429 br_429 en vdd gnd
+ write_driver
Xwrite_driver430
+ data_430 bl_430 br_430 en vdd gnd
+ write_driver
Xwrite_driver431
+ data_431 bl_431 br_431 en vdd gnd
+ write_driver
Xwrite_driver432
+ data_432 bl_432 br_432 en vdd gnd
+ write_driver
Xwrite_driver433
+ data_433 bl_433 br_433 en vdd gnd
+ write_driver
Xwrite_driver434
+ data_434 bl_434 br_434 en vdd gnd
+ write_driver
Xwrite_driver435
+ data_435 bl_435 br_435 en vdd gnd
+ write_driver
Xwrite_driver436
+ data_436 bl_436 br_436 en vdd gnd
+ write_driver
Xwrite_driver437
+ data_437 bl_437 br_437 en vdd gnd
+ write_driver
Xwrite_driver438
+ data_438 bl_438 br_438 en vdd gnd
+ write_driver
Xwrite_driver439
+ data_439 bl_439 br_439 en vdd gnd
+ write_driver
Xwrite_driver440
+ data_440 bl_440 br_440 en vdd gnd
+ write_driver
Xwrite_driver441
+ data_441 bl_441 br_441 en vdd gnd
+ write_driver
Xwrite_driver442
+ data_442 bl_442 br_442 en vdd gnd
+ write_driver
Xwrite_driver443
+ data_443 bl_443 br_443 en vdd gnd
+ write_driver
Xwrite_driver444
+ data_444 bl_444 br_444 en vdd gnd
+ write_driver
Xwrite_driver445
+ data_445 bl_445 br_445 en vdd gnd
+ write_driver
Xwrite_driver446
+ data_446 bl_446 br_446 en vdd gnd
+ write_driver
Xwrite_driver447
+ data_447 bl_447 br_447 en vdd gnd
+ write_driver
Xwrite_driver448
+ data_448 bl_448 br_448 en vdd gnd
+ write_driver
Xwrite_driver449
+ data_449 bl_449 br_449 en vdd gnd
+ write_driver
Xwrite_driver450
+ data_450 bl_450 br_450 en vdd gnd
+ write_driver
Xwrite_driver451
+ data_451 bl_451 br_451 en vdd gnd
+ write_driver
Xwrite_driver452
+ data_452 bl_452 br_452 en vdd gnd
+ write_driver
Xwrite_driver453
+ data_453 bl_453 br_453 en vdd gnd
+ write_driver
Xwrite_driver454
+ data_454 bl_454 br_454 en vdd gnd
+ write_driver
Xwrite_driver455
+ data_455 bl_455 br_455 en vdd gnd
+ write_driver
Xwrite_driver456
+ data_456 bl_456 br_456 en vdd gnd
+ write_driver
Xwrite_driver457
+ data_457 bl_457 br_457 en vdd gnd
+ write_driver
Xwrite_driver458
+ data_458 bl_458 br_458 en vdd gnd
+ write_driver
Xwrite_driver459
+ data_459 bl_459 br_459 en vdd gnd
+ write_driver
Xwrite_driver460
+ data_460 bl_460 br_460 en vdd gnd
+ write_driver
Xwrite_driver461
+ data_461 bl_461 br_461 en vdd gnd
+ write_driver
Xwrite_driver462
+ data_462 bl_462 br_462 en vdd gnd
+ write_driver
Xwrite_driver463
+ data_463 bl_463 br_463 en vdd gnd
+ write_driver
Xwrite_driver464
+ data_464 bl_464 br_464 en vdd gnd
+ write_driver
Xwrite_driver465
+ data_465 bl_465 br_465 en vdd gnd
+ write_driver
Xwrite_driver466
+ data_466 bl_466 br_466 en vdd gnd
+ write_driver
Xwrite_driver467
+ data_467 bl_467 br_467 en vdd gnd
+ write_driver
Xwrite_driver468
+ data_468 bl_468 br_468 en vdd gnd
+ write_driver
Xwrite_driver469
+ data_469 bl_469 br_469 en vdd gnd
+ write_driver
Xwrite_driver470
+ data_470 bl_470 br_470 en vdd gnd
+ write_driver
Xwrite_driver471
+ data_471 bl_471 br_471 en vdd gnd
+ write_driver
Xwrite_driver472
+ data_472 bl_472 br_472 en vdd gnd
+ write_driver
Xwrite_driver473
+ data_473 bl_473 br_473 en vdd gnd
+ write_driver
Xwrite_driver474
+ data_474 bl_474 br_474 en vdd gnd
+ write_driver
Xwrite_driver475
+ data_475 bl_475 br_475 en vdd gnd
+ write_driver
Xwrite_driver476
+ data_476 bl_476 br_476 en vdd gnd
+ write_driver
Xwrite_driver477
+ data_477 bl_477 br_477 en vdd gnd
+ write_driver
Xwrite_driver478
+ data_478 bl_478 br_478 en vdd gnd
+ write_driver
Xwrite_driver479
+ data_479 bl_479 br_479 en vdd gnd
+ write_driver
Xwrite_driver480
+ data_480 bl_480 br_480 en vdd gnd
+ write_driver
Xwrite_driver481
+ data_481 bl_481 br_481 en vdd gnd
+ write_driver
Xwrite_driver482
+ data_482 bl_482 br_482 en vdd gnd
+ write_driver
Xwrite_driver483
+ data_483 bl_483 br_483 en vdd gnd
+ write_driver
Xwrite_driver484
+ data_484 bl_484 br_484 en vdd gnd
+ write_driver
Xwrite_driver485
+ data_485 bl_485 br_485 en vdd gnd
+ write_driver
Xwrite_driver486
+ data_486 bl_486 br_486 en vdd gnd
+ write_driver
Xwrite_driver487
+ data_487 bl_487 br_487 en vdd gnd
+ write_driver
Xwrite_driver488
+ data_488 bl_488 br_488 en vdd gnd
+ write_driver
Xwrite_driver489
+ data_489 bl_489 br_489 en vdd gnd
+ write_driver
Xwrite_driver490
+ data_490 bl_490 br_490 en vdd gnd
+ write_driver
Xwrite_driver491
+ data_491 bl_491 br_491 en vdd gnd
+ write_driver
Xwrite_driver492
+ data_492 bl_492 br_492 en vdd gnd
+ write_driver
Xwrite_driver493
+ data_493 bl_493 br_493 en vdd gnd
+ write_driver
Xwrite_driver494
+ data_494 bl_494 br_494 en vdd gnd
+ write_driver
Xwrite_driver495
+ data_495 bl_495 br_495 en vdd gnd
+ write_driver
Xwrite_driver496
+ data_496 bl_496 br_496 en vdd gnd
+ write_driver
Xwrite_driver497
+ data_497 bl_497 br_497 en vdd gnd
+ write_driver
Xwrite_driver498
+ data_498 bl_498 br_498 en vdd gnd
+ write_driver
Xwrite_driver499
+ data_499 bl_499 br_499 en vdd gnd
+ write_driver
Xwrite_driver500
+ data_500 bl_500 br_500 en vdd gnd
+ write_driver
Xwrite_driver501
+ data_501 bl_501 br_501 en vdd gnd
+ write_driver
Xwrite_driver502
+ data_502 bl_502 br_502 en vdd gnd
+ write_driver
Xwrite_driver503
+ data_503 bl_503 br_503 en vdd gnd
+ write_driver
Xwrite_driver504
+ data_504 bl_504 br_504 en vdd gnd
+ write_driver
Xwrite_driver505
+ data_505 bl_505 br_505 en vdd gnd
+ write_driver
Xwrite_driver506
+ data_506 bl_506 br_506 en vdd gnd
+ write_driver
Xwrite_driver507
+ data_507 bl_507 br_507 en vdd gnd
+ write_driver
Xwrite_driver508
+ data_508 bl_508 br_508 en vdd gnd
+ write_driver
Xwrite_driver509
+ data_509 bl_509 br_509 en vdd gnd
+ write_driver
Xwrite_driver510
+ data_510 bl_510 br_510 en vdd gnd
+ write_driver
Xwrite_driver511
+ data_511 bl_511 br_511 en vdd gnd
+ write_driver
.ENDS freepdk45_sram_1rw0r_45x512_write_driver_array

.SUBCKT freepdk45_sram_1rw0r_45x512_port_data
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66
+ bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72
+ br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77
+ bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83
+ br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88
+ bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94
+ br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99
+ bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104
+ bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109
+ bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114
+ bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119
+ bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124
+ bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129
+ bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134
+ bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139
+ bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144
+ bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149
+ bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154
+ bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159
+ bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164
+ bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169
+ bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174
+ bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179
+ bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184
+ bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189
+ bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194
+ bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199
+ bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204
+ bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209
+ bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214
+ bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219
+ bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224
+ bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229
+ bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234
+ bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239
+ bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244
+ bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249
+ bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254
+ bl_255 br_255 bl_256 br_256 bl_257 br_257 bl_258 br_258 bl_259 br_259
+ bl_260 br_260 bl_261 br_261 bl_262 br_262 bl_263 br_263 bl_264 br_264
+ bl_265 br_265 bl_266 br_266 bl_267 br_267 bl_268 br_268 bl_269 br_269
+ bl_270 br_270 bl_271 br_271 bl_272 br_272 bl_273 br_273 bl_274 br_274
+ bl_275 br_275 bl_276 br_276 bl_277 br_277 bl_278 br_278 bl_279 br_279
+ bl_280 br_280 bl_281 br_281 bl_282 br_282 bl_283 br_283 bl_284 br_284
+ bl_285 br_285 bl_286 br_286 bl_287 br_287 bl_288 br_288 bl_289 br_289
+ bl_290 br_290 bl_291 br_291 bl_292 br_292 bl_293 br_293 bl_294 br_294
+ bl_295 br_295 bl_296 br_296 bl_297 br_297 bl_298 br_298 bl_299 br_299
+ bl_300 br_300 bl_301 br_301 bl_302 br_302 bl_303 br_303 bl_304 br_304
+ bl_305 br_305 bl_306 br_306 bl_307 br_307 bl_308 br_308 bl_309 br_309
+ bl_310 br_310 bl_311 br_311 bl_312 br_312 bl_313 br_313 bl_314 br_314
+ bl_315 br_315 bl_316 br_316 bl_317 br_317 bl_318 br_318 bl_319 br_319
+ bl_320 br_320 bl_321 br_321 bl_322 br_322 bl_323 br_323 bl_324 br_324
+ bl_325 br_325 bl_326 br_326 bl_327 br_327 bl_328 br_328 bl_329 br_329
+ bl_330 br_330 bl_331 br_331 bl_332 br_332 bl_333 br_333 bl_334 br_334
+ bl_335 br_335 bl_336 br_336 bl_337 br_337 bl_338 br_338 bl_339 br_339
+ bl_340 br_340 bl_341 br_341 bl_342 br_342 bl_343 br_343 bl_344 br_344
+ bl_345 br_345 bl_346 br_346 bl_347 br_347 bl_348 br_348 bl_349 br_349
+ bl_350 br_350 bl_351 br_351 bl_352 br_352 bl_353 br_353 bl_354 br_354
+ bl_355 br_355 bl_356 br_356 bl_357 br_357 bl_358 br_358 bl_359 br_359
+ bl_360 br_360 bl_361 br_361 bl_362 br_362 bl_363 br_363 bl_364 br_364
+ bl_365 br_365 bl_366 br_366 bl_367 br_367 bl_368 br_368 bl_369 br_369
+ bl_370 br_370 bl_371 br_371 bl_372 br_372 bl_373 br_373 bl_374 br_374
+ bl_375 br_375 bl_376 br_376 bl_377 br_377 bl_378 br_378 bl_379 br_379
+ bl_380 br_380 bl_381 br_381 bl_382 br_382 bl_383 br_383 bl_384 br_384
+ bl_385 br_385 bl_386 br_386 bl_387 br_387 bl_388 br_388 bl_389 br_389
+ bl_390 br_390 bl_391 br_391 bl_392 br_392 bl_393 br_393 bl_394 br_394
+ bl_395 br_395 bl_396 br_396 bl_397 br_397 bl_398 br_398 bl_399 br_399
+ bl_400 br_400 bl_401 br_401 bl_402 br_402 bl_403 br_403 bl_404 br_404
+ bl_405 br_405 bl_406 br_406 bl_407 br_407 bl_408 br_408 bl_409 br_409
+ bl_410 br_410 bl_411 br_411 bl_412 br_412 bl_413 br_413 bl_414 br_414
+ bl_415 br_415 bl_416 br_416 bl_417 br_417 bl_418 br_418 bl_419 br_419
+ bl_420 br_420 bl_421 br_421 bl_422 br_422 bl_423 br_423 bl_424 br_424
+ bl_425 br_425 bl_426 br_426 bl_427 br_427 bl_428 br_428 bl_429 br_429
+ bl_430 br_430 bl_431 br_431 bl_432 br_432 bl_433 br_433 bl_434 br_434
+ bl_435 br_435 bl_436 br_436 bl_437 br_437 bl_438 br_438 bl_439 br_439
+ bl_440 br_440 bl_441 br_441 bl_442 br_442 bl_443 br_443 bl_444 br_444
+ bl_445 br_445 bl_446 br_446 bl_447 br_447 bl_448 br_448 bl_449 br_449
+ bl_450 br_450 bl_451 br_451 bl_452 br_452 bl_453 br_453 bl_454 br_454
+ bl_455 br_455 bl_456 br_456 bl_457 br_457 bl_458 br_458 bl_459 br_459
+ bl_460 br_460 bl_461 br_461 bl_462 br_462 bl_463 br_463 bl_464 br_464
+ bl_465 br_465 bl_466 br_466 bl_467 br_467 bl_468 br_468 bl_469 br_469
+ bl_470 br_470 bl_471 br_471 bl_472 br_472 bl_473 br_473 bl_474 br_474
+ bl_475 br_475 bl_476 br_476 bl_477 br_477 bl_478 br_478 bl_479 br_479
+ bl_480 br_480 bl_481 br_481 bl_482 br_482 bl_483 br_483 bl_484 br_484
+ bl_485 br_485 bl_486 br_486 bl_487 br_487 bl_488 br_488 bl_489 br_489
+ bl_490 br_490 bl_491 br_491 bl_492 br_492 bl_493 br_493 bl_494 br_494
+ bl_495 br_495 bl_496 br_496 bl_497 br_497 bl_498 br_498 bl_499 br_499
+ bl_500 br_500 bl_501 br_501 bl_502 br_502 bl_503 br_503 bl_504 br_504
+ bl_505 br_505 bl_506 br_506 bl_507 br_507 bl_508 br_508 bl_509 br_509
+ bl_510 br_510 bl_511 br_511 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5
+ dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14
+ dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22
+ dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30
+ dout_31 dout_32 dout_33 dout_34 dout_35 dout_36 dout_37 dout_38
+ dout_39 dout_40 dout_41 dout_42 dout_43 dout_44 dout_45 dout_46
+ dout_47 dout_48 dout_49 dout_50 dout_51 dout_52 dout_53 dout_54
+ dout_55 dout_56 dout_57 dout_58 dout_59 dout_60 dout_61 dout_62
+ dout_63 dout_64 dout_65 dout_66 dout_67 dout_68 dout_69 dout_70
+ dout_71 dout_72 dout_73 dout_74 dout_75 dout_76 dout_77 dout_78
+ dout_79 dout_80 dout_81 dout_82 dout_83 dout_84 dout_85 dout_86
+ dout_87 dout_88 dout_89 dout_90 dout_91 dout_92 dout_93 dout_94
+ dout_95 dout_96 dout_97 dout_98 dout_99 dout_100 dout_101 dout_102
+ dout_103 dout_104 dout_105 dout_106 dout_107 dout_108 dout_109
+ dout_110 dout_111 dout_112 dout_113 dout_114 dout_115 dout_116
+ dout_117 dout_118 dout_119 dout_120 dout_121 dout_122 dout_123
+ dout_124 dout_125 dout_126 dout_127 dout_128 dout_129 dout_130
+ dout_131 dout_132 dout_133 dout_134 dout_135 dout_136 dout_137
+ dout_138 dout_139 dout_140 dout_141 dout_142 dout_143 dout_144
+ dout_145 dout_146 dout_147 dout_148 dout_149 dout_150 dout_151
+ dout_152 dout_153 dout_154 dout_155 dout_156 dout_157 dout_158
+ dout_159 dout_160 dout_161 dout_162 dout_163 dout_164 dout_165
+ dout_166 dout_167 dout_168 dout_169 dout_170 dout_171 dout_172
+ dout_173 dout_174 dout_175 dout_176 dout_177 dout_178 dout_179
+ dout_180 dout_181 dout_182 dout_183 dout_184 dout_185 dout_186
+ dout_187 dout_188 dout_189 dout_190 dout_191 dout_192 dout_193
+ dout_194 dout_195 dout_196 dout_197 dout_198 dout_199 dout_200
+ dout_201 dout_202 dout_203 dout_204 dout_205 dout_206 dout_207
+ dout_208 dout_209 dout_210 dout_211 dout_212 dout_213 dout_214
+ dout_215 dout_216 dout_217 dout_218 dout_219 dout_220 dout_221
+ dout_222 dout_223 dout_224 dout_225 dout_226 dout_227 dout_228
+ dout_229 dout_230 dout_231 dout_232 dout_233 dout_234 dout_235
+ dout_236 dout_237 dout_238 dout_239 dout_240 dout_241 dout_242
+ dout_243 dout_244 dout_245 dout_246 dout_247 dout_248 dout_249
+ dout_250 dout_251 dout_252 dout_253 dout_254 dout_255 dout_256
+ dout_257 dout_258 dout_259 dout_260 dout_261 dout_262 dout_263
+ dout_264 dout_265 dout_266 dout_267 dout_268 dout_269 dout_270
+ dout_271 dout_272 dout_273 dout_274 dout_275 dout_276 dout_277
+ dout_278 dout_279 dout_280 dout_281 dout_282 dout_283 dout_284
+ dout_285 dout_286 dout_287 dout_288 dout_289 dout_290 dout_291
+ dout_292 dout_293 dout_294 dout_295 dout_296 dout_297 dout_298
+ dout_299 dout_300 dout_301 dout_302 dout_303 dout_304 dout_305
+ dout_306 dout_307 dout_308 dout_309 dout_310 dout_311 dout_312
+ dout_313 dout_314 dout_315 dout_316 dout_317 dout_318 dout_319
+ dout_320 dout_321 dout_322 dout_323 dout_324 dout_325 dout_326
+ dout_327 dout_328 dout_329 dout_330 dout_331 dout_332 dout_333
+ dout_334 dout_335 dout_336 dout_337 dout_338 dout_339 dout_340
+ dout_341 dout_342 dout_343 dout_344 dout_345 dout_346 dout_347
+ dout_348 dout_349 dout_350 dout_351 dout_352 dout_353 dout_354
+ dout_355 dout_356 dout_357 dout_358 dout_359 dout_360 dout_361
+ dout_362 dout_363 dout_364 dout_365 dout_366 dout_367 dout_368
+ dout_369 dout_370 dout_371 dout_372 dout_373 dout_374 dout_375
+ dout_376 dout_377 dout_378 dout_379 dout_380 dout_381 dout_382
+ dout_383 dout_384 dout_385 dout_386 dout_387 dout_388 dout_389
+ dout_390 dout_391 dout_392 dout_393 dout_394 dout_395 dout_396
+ dout_397 dout_398 dout_399 dout_400 dout_401 dout_402 dout_403
+ dout_404 dout_405 dout_406 dout_407 dout_408 dout_409 dout_410
+ dout_411 dout_412 dout_413 dout_414 dout_415 dout_416 dout_417
+ dout_418 dout_419 dout_420 dout_421 dout_422 dout_423 dout_424
+ dout_425 dout_426 dout_427 dout_428 dout_429 dout_430 dout_431
+ dout_432 dout_433 dout_434 dout_435 dout_436 dout_437 dout_438
+ dout_439 dout_440 dout_441 dout_442 dout_443 dout_444 dout_445
+ dout_446 dout_447 dout_448 dout_449 dout_450 dout_451 dout_452
+ dout_453 dout_454 dout_455 dout_456 dout_457 dout_458 dout_459
+ dout_460 dout_461 dout_462 dout_463 dout_464 dout_465 dout_466
+ dout_467 dout_468 dout_469 dout_470 dout_471 dout_472 dout_473
+ dout_474 dout_475 dout_476 dout_477 dout_478 dout_479 dout_480
+ dout_481 dout_482 dout_483 dout_484 dout_485 dout_486 dout_487
+ dout_488 dout_489 dout_490 dout_491 dout_492 dout_493 dout_494
+ dout_495 dout_496 dout_497 dout_498 dout_499 dout_500 dout_501
+ dout_502 dout_503 dout_504 dout_505 dout_506 dout_507 dout_508
+ dout_509 dout_510 dout_511 din_0 din_1 din_2 din_3 din_4 din_5 din_6
+ din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16
+ din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26
+ din_27 din_28 din_29 din_30 din_31 din_32 din_33 din_34 din_35 din_36
+ din_37 din_38 din_39 din_40 din_41 din_42 din_43 din_44 din_45 din_46
+ din_47 din_48 din_49 din_50 din_51 din_52 din_53 din_54 din_55 din_56
+ din_57 din_58 din_59 din_60 din_61 din_62 din_63 din_64 din_65 din_66
+ din_67 din_68 din_69 din_70 din_71 din_72 din_73 din_74 din_75 din_76
+ din_77 din_78 din_79 din_80 din_81 din_82 din_83 din_84 din_85 din_86
+ din_87 din_88 din_89 din_90 din_91 din_92 din_93 din_94 din_95 din_96
+ din_97 din_98 din_99 din_100 din_101 din_102 din_103 din_104 din_105
+ din_106 din_107 din_108 din_109 din_110 din_111 din_112 din_113
+ din_114 din_115 din_116 din_117 din_118 din_119 din_120 din_121
+ din_122 din_123 din_124 din_125 din_126 din_127 din_128 din_129
+ din_130 din_131 din_132 din_133 din_134 din_135 din_136 din_137
+ din_138 din_139 din_140 din_141 din_142 din_143 din_144 din_145
+ din_146 din_147 din_148 din_149 din_150 din_151 din_152 din_153
+ din_154 din_155 din_156 din_157 din_158 din_159 din_160 din_161
+ din_162 din_163 din_164 din_165 din_166 din_167 din_168 din_169
+ din_170 din_171 din_172 din_173 din_174 din_175 din_176 din_177
+ din_178 din_179 din_180 din_181 din_182 din_183 din_184 din_185
+ din_186 din_187 din_188 din_189 din_190 din_191 din_192 din_193
+ din_194 din_195 din_196 din_197 din_198 din_199 din_200 din_201
+ din_202 din_203 din_204 din_205 din_206 din_207 din_208 din_209
+ din_210 din_211 din_212 din_213 din_214 din_215 din_216 din_217
+ din_218 din_219 din_220 din_221 din_222 din_223 din_224 din_225
+ din_226 din_227 din_228 din_229 din_230 din_231 din_232 din_233
+ din_234 din_235 din_236 din_237 din_238 din_239 din_240 din_241
+ din_242 din_243 din_244 din_245 din_246 din_247 din_248 din_249
+ din_250 din_251 din_252 din_253 din_254 din_255 din_256 din_257
+ din_258 din_259 din_260 din_261 din_262 din_263 din_264 din_265
+ din_266 din_267 din_268 din_269 din_270 din_271 din_272 din_273
+ din_274 din_275 din_276 din_277 din_278 din_279 din_280 din_281
+ din_282 din_283 din_284 din_285 din_286 din_287 din_288 din_289
+ din_290 din_291 din_292 din_293 din_294 din_295 din_296 din_297
+ din_298 din_299 din_300 din_301 din_302 din_303 din_304 din_305
+ din_306 din_307 din_308 din_309 din_310 din_311 din_312 din_313
+ din_314 din_315 din_316 din_317 din_318 din_319 din_320 din_321
+ din_322 din_323 din_324 din_325 din_326 din_327 din_328 din_329
+ din_330 din_331 din_332 din_333 din_334 din_335 din_336 din_337
+ din_338 din_339 din_340 din_341 din_342 din_343 din_344 din_345
+ din_346 din_347 din_348 din_349 din_350 din_351 din_352 din_353
+ din_354 din_355 din_356 din_357 din_358 din_359 din_360 din_361
+ din_362 din_363 din_364 din_365 din_366 din_367 din_368 din_369
+ din_370 din_371 din_372 din_373 din_374 din_375 din_376 din_377
+ din_378 din_379 din_380 din_381 din_382 din_383 din_384 din_385
+ din_386 din_387 din_388 din_389 din_390 din_391 din_392 din_393
+ din_394 din_395 din_396 din_397 din_398 din_399 din_400 din_401
+ din_402 din_403 din_404 din_405 din_406 din_407 din_408 din_409
+ din_410 din_411 din_412 din_413 din_414 din_415 din_416 din_417
+ din_418 din_419 din_420 din_421 din_422 din_423 din_424 din_425
+ din_426 din_427 din_428 din_429 din_430 din_431 din_432 din_433
+ din_434 din_435 din_436 din_437 din_438 din_439 din_440 din_441
+ din_442 din_443 din_444 din_445 din_446 din_447 din_448 din_449
+ din_450 din_451 din_452 din_453 din_454 din_455 din_456 din_457
+ din_458 din_459 din_460 din_461 din_462 din_463 din_464 din_465
+ din_466 din_467 din_468 din_469 din_470 din_471 din_472 din_473
+ din_474 din_475 din_476 din_477 din_478 din_479 din_480 din_481
+ din_482 din_483 din_484 din_485 din_486 din_487 din_488 din_489
+ din_490 din_491 din_492 din_493 din_494 din_495 din_496 din_497
+ din_498 din_499 din_500 din_501 din_502 din_503 din_504 din_505
+ din_506 din_507 din_508 din_509 din_510 din_511 s_en p_en_bar w_en vdd
+ gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INOUT : bl_256 
* INOUT : br_256 
* INOUT : bl_257 
* INOUT : br_257 
* INOUT : bl_258 
* INOUT : br_258 
* INOUT : bl_259 
* INOUT : br_259 
* INOUT : bl_260 
* INOUT : br_260 
* INOUT : bl_261 
* INOUT : br_261 
* INOUT : bl_262 
* INOUT : br_262 
* INOUT : bl_263 
* INOUT : br_263 
* INOUT : bl_264 
* INOUT : br_264 
* INOUT : bl_265 
* INOUT : br_265 
* INOUT : bl_266 
* INOUT : br_266 
* INOUT : bl_267 
* INOUT : br_267 
* INOUT : bl_268 
* INOUT : br_268 
* INOUT : bl_269 
* INOUT : br_269 
* INOUT : bl_270 
* INOUT : br_270 
* INOUT : bl_271 
* INOUT : br_271 
* INOUT : bl_272 
* INOUT : br_272 
* INOUT : bl_273 
* INOUT : br_273 
* INOUT : bl_274 
* INOUT : br_274 
* INOUT : bl_275 
* INOUT : br_275 
* INOUT : bl_276 
* INOUT : br_276 
* INOUT : bl_277 
* INOUT : br_277 
* INOUT : bl_278 
* INOUT : br_278 
* INOUT : bl_279 
* INOUT : br_279 
* INOUT : bl_280 
* INOUT : br_280 
* INOUT : bl_281 
* INOUT : br_281 
* INOUT : bl_282 
* INOUT : br_282 
* INOUT : bl_283 
* INOUT : br_283 
* INOUT : bl_284 
* INOUT : br_284 
* INOUT : bl_285 
* INOUT : br_285 
* INOUT : bl_286 
* INOUT : br_286 
* INOUT : bl_287 
* INOUT : br_287 
* INOUT : bl_288 
* INOUT : br_288 
* INOUT : bl_289 
* INOUT : br_289 
* INOUT : bl_290 
* INOUT : br_290 
* INOUT : bl_291 
* INOUT : br_291 
* INOUT : bl_292 
* INOUT : br_292 
* INOUT : bl_293 
* INOUT : br_293 
* INOUT : bl_294 
* INOUT : br_294 
* INOUT : bl_295 
* INOUT : br_295 
* INOUT : bl_296 
* INOUT : br_296 
* INOUT : bl_297 
* INOUT : br_297 
* INOUT : bl_298 
* INOUT : br_298 
* INOUT : bl_299 
* INOUT : br_299 
* INOUT : bl_300 
* INOUT : br_300 
* INOUT : bl_301 
* INOUT : br_301 
* INOUT : bl_302 
* INOUT : br_302 
* INOUT : bl_303 
* INOUT : br_303 
* INOUT : bl_304 
* INOUT : br_304 
* INOUT : bl_305 
* INOUT : br_305 
* INOUT : bl_306 
* INOUT : br_306 
* INOUT : bl_307 
* INOUT : br_307 
* INOUT : bl_308 
* INOUT : br_308 
* INOUT : bl_309 
* INOUT : br_309 
* INOUT : bl_310 
* INOUT : br_310 
* INOUT : bl_311 
* INOUT : br_311 
* INOUT : bl_312 
* INOUT : br_312 
* INOUT : bl_313 
* INOUT : br_313 
* INOUT : bl_314 
* INOUT : br_314 
* INOUT : bl_315 
* INOUT : br_315 
* INOUT : bl_316 
* INOUT : br_316 
* INOUT : bl_317 
* INOUT : br_317 
* INOUT : bl_318 
* INOUT : br_318 
* INOUT : bl_319 
* INOUT : br_319 
* INOUT : bl_320 
* INOUT : br_320 
* INOUT : bl_321 
* INOUT : br_321 
* INOUT : bl_322 
* INOUT : br_322 
* INOUT : bl_323 
* INOUT : br_323 
* INOUT : bl_324 
* INOUT : br_324 
* INOUT : bl_325 
* INOUT : br_325 
* INOUT : bl_326 
* INOUT : br_326 
* INOUT : bl_327 
* INOUT : br_327 
* INOUT : bl_328 
* INOUT : br_328 
* INOUT : bl_329 
* INOUT : br_329 
* INOUT : bl_330 
* INOUT : br_330 
* INOUT : bl_331 
* INOUT : br_331 
* INOUT : bl_332 
* INOUT : br_332 
* INOUT : bl_333 
* INOUT : br_333 
* INOUT : bl_334 
* INOUT : br_334 
* INOUT : bl_335 
* INOUT : br_335 
* INOUT : bl_336 
* INOUT : br_336 
* INOUT : bl_337 
* INOUT : br_337 
* INOUT : bl_338 
* INOUT : br_338 
* INOUT : bl_339 
* INOUT : br_339 
* INOUT : bl_340 
* INOUT : br_340 
* INOUT : bl_341 
* INOUT : br_341 
* INOUT : bl_342 
* INOUT : br_342 
* INOUT : bl_343 
* INOUT : br_343 
* INOUT : bl_344 
* INOUT : br_344 
* INOUT : bl_345 
* INOUT : br_345 
* INOUT : bl_346 
* INOUT : br_346 
* INOUT : bl_347 
* INOUT : br_347 
* INOUT : bl_348 
* INOUT : br_348 
* INOUT : bl_349 
* INOUT : br_349 
* INOUT : bl_350 
* INOUT : br_350 
* INOUT : bl_351 
* INOUT : br_351 
* INOUT : bl_352 
* INOUT : br_352 
* INOUT : bl_353 
* INOUT : br_353 
* INOUT : bl_354 
* INOUT : br_354 
* INOUT : bl_355 
* INOUT : br_355 
* INOUT : bl_356 
* INOUT : br_356 
* INOUT : bl_357 
* INOUT : br_357 
* INOUT : bl_358 
* INOUT : br_358 
* INOUT : bl_359 
* INOUT : br_359 
* INOUT : bl_360 
* INOUT : br_360 
* INOUT : bl_361 
* INOUT : br_361 
* INOUT : bl_362 
* INOUT : br_362 
* INOUT : bl_363 
* INOUT : br_363 
* INOUT : bl_364 
* INOUT : br_364 
* INOUT : bl_365 
* INOUT : br_365 
* INOUT : bl_366 
* INOUT : br_366 
* INOUT : bl_367 
* INOUT : br_367 
* INOUT : bl_368 
* INOUT : br_368 
* INOUT : bl_369 
* INOUT : br_369 
* INOUT : bl_370 
* INOUT : br_370 
* INOUT : bl_371 
* INOUT : br_371 
* INOUT : bl_372 
* INOUT : br_372 
* INOUT : bl_373 
* INOUT : br_373 
* INOUT : bl_374 
* INOUT : br_374 
* INOUT : bl_375 
* INOUT : br_375 
* INOUT : bl_376 
* INOUT : br_376 
* INOUT : bl_377 
* INOUT : br_377 
* INOUT : bl_378 
* INOUT : br_378 
* INOUT : bl_379 
* INOUT : br_379 
* INOUT : bl_380 
* INOUT : br_380 
* INOUT : bl_381 
* INOUT : br_381 
* INOUT : bl_382 
* INOUT : br_382 
* INOUT : bl_383 
* INOUT : br_383 
* INOUT : bl_384 
* INOUT : br_384 
* INOUT : bl_385 
* INOUT : br_385 
* INOUT : bl_386 
* INOUT : br_386 
* INOUT : bl_387 
* INOUT : br_387 
* INOUT : bl_388 
* INOUT : br_388 
* INOUT : bl_389 
* INOUT : br_389 
* INOUT : bl_390 
* INOUT : br_390 
* INOUT : bl_391 
* INOUT : br_391 
* INOUT : bl_392 
* INOUT : br_392 
* INOUT : bl_393 
* INOUT : br_393 
* INOUT : bl_394 
* INOUT : br_394 
* INOUT : bl_395 
* INOUT : br_395 
* INOUT : bl_396 
* INOUT : br_396 
* INOUT : bl_397 
* INOUT : br_397 
* INOUT : bl_398 
* INOUT : br_398 
* INOUT : bl_399 
* INOUT : br_399 
* INOUT : bl_400 
* INOUT : br_400 
* INOUT : bl_401 
* INOUT : br_401 
* INOUT : bl_402 
* INOUT : br_402 
* INOUT : bl_403 
* INOUT : br_403 
* INOUT : bl_404 
* INOUT : br_404 
* INOUT : bl_405 
* INOUT : br_405 
* INOUT : bl_406 
* INOUT : br_406 
* INOUT : bl_407 
* INOUT : br_407 
* INOUT : bl_408 
* INOUT : br_408 
* INOUT : bl_409 
* INOUT : br_409 
* INOUT : bl_410 
* INOUT : br_410 
* INOUT : bl_411 
* INOUT : br_411 
* INOUT : bl_412 
* INOUT : br_412 
* INOUT : bl_413 
* INOUT : br_413 
* INOUT : bl_414 
* INOUT : br_414 
* INOUT : bl_415 
* INOUT : br_415 
* INOUT : bl_416 
* INOUT : br_416 
* INOUT : bl_417 
* INOUT : br_417 
* INOUT : bl_418 
* INOUT : br_418 
* INOUT : bl_419 
* INOUT : br_419 
* INOUT : bl_420 
* INOUT : br_420 
* INOUT : bl_421 
* INOUT : br_421 
* INOUT : bl_422 
* INOUT : br_422 
* INOUT : bl_423 
* INOUT : br_423 
* INOUT : bl_424 
* INOUT : br_424 
* INOUT : bl_425 
* INOUT : br_425 
* INOUT : bl_426 
* INOUT : br_426 
* INOUT : bl_427 
* INOUT : br_427 
* INOUT : bl_428 
* INOUT : br_428 
* INOUT : bl_429 
* INOUT : br_429 
* INOUT : bl_430 
* INOUT : br_430 
* INOUT : bl_431 
* INOUT : br_431 
* INOUT : bl_432 
* INOUT : br_432 
* INOUT : bl_433 
* INOUT : br_433 
* INOUT : bl_434 
* INOUT : br_434 
* INOUT : bl_435 
* INOUT : br_435 
* INOUT : bl_436 
* INOUT : br_436 
* INOUT : bl_437 
* INOUT : br_437 
* INOUT : bl_438 
* INOUT : br_438 
* INOUT : bl_439 
* INOUT : br_439 
* INOUT : bl_440 
* INOUT : br_440 
* INOUT : bl_441 
* INOUT : br_441 
* INOUT : bl_442 
* INOUT : br_442 
* INOUT : bl_443 
* INOUT : br_443 
* INOUT : bl_444 
* INOUT : br_444 
* INOUT : bl_445 
* INOUT : br_445 
* INOUT : bl_446 
* INOUT : br_446 
* INOUT : bl_447 
* INOUT : br_447 
* INOUT : bl_448 
* INOUT : br_448 
* INOUT : bl_449 
* INOUT : br_449 
* INOUT : bl_450 
* INOUT : br_450 
* INOUT : bl_451 
* INOUT : br_451 
* INOUT : bl_452 
* INOUT : br_452 
* INOUT : bl_453 
* INOUT : br_453 
* INOUT : bl_454 
* INOUT : br_454 
* INOUT : bl_455 
* INOUT : br_455 
* INOUT : bl_456 
* INOUT : br_456 
* INOUT : bl_457 
* INOUT : br_457 
* INOUT : bl_458 
* INOUT : br_458 
* INOUT : bl_459 
* INOUT : br_459 
* INOUT : bl_460 
* INOUT : br_460 
* INOUT : bl_461 
* INOUT : br_461 
* INOUT : bl_462 
* INOUT : br_462 
* INOUT : bl_463 
* INOUT : br_463 
* INOUT : bl_464 
* INOUT : br_464 
* INOUT : bl_465 
* INOUT : br_465 
* INOUT : bl_466 
* INOUT : br_466 
* INOUT : bl_467 
* INOUT : br_467 
* INOUT : bl_468 
* INOUT : br_468 
* INOUT : bl_469 
* INOUT : br_469 
* INOUT : bl_470 
* INOUT : br_470 
* INOUT : bl_471 
* INOUT : br_471 
* INOUT : bl_472 
* INOUT : br_472 
* INOUT : bl_473 
* INOUT : br_473 
* INOUT : bl_474 
* INOUT : br_474 
* INOUT : bl_475 
* INOUT : br_475 
* INOUT : bl_476 
* INOUT : br_476 
* INOUT : bl_477 
* INOUT : br_477 
* INOUT : bl_478 
* INOUT : br_478 
* INOUT : bl_479 
* INOUT : br_479 
* INOUT : bl_480 
* INOUT : br_480 
* INOUT : bl_481 
* INOUT : br_481 
* INOUT : bl_482 
* INOUT : br_482 
* INOUT : bl_483 
* INOUT : br_483 
* INOUT : bl_484 
* INOUT : br_484 
* INOUT : bl_485 
* INOUT : br_485 
* INOUT : bl_486 
* INOUT : br_486 
* INOUT : bl_487 
* INOUT : br_487 
* INOUT : bl_488 
* INOUT : br_488 
* INOUT : bl_489 
* INOUT : br_489 
* INOUT : bl_490 
* INOUT : br_490 
* INOUT : bl_491 
* INOUT : br_491 
* INOUT : bl_492 
* INOUT : br_492 
* INOUT : bl_493 
* INOUT : br_493 
* INOUT : bl_494 
* INOUT : br_494 
* INOUT : bl_495 
* INOUT : br_495 
* INOUT : bl_496 
* INOUT : br_496 
* INOUT : bl_497 
* INOUT : br_497 
* INOUT : bl_498 
* INOUT : br_498 
* INOUT : bl_499 
* INOUT : br_499 
* INOUT : bl_500 
* INOUT : br_500 
* INOUT : bl_501 
* INOUT : br_501 
* INOUT : bl_502 
* INOUT : br_502 
* INOUT : bl_503 
* INOUT : br_503 
* INOUT : bl_504 
* INOUT : br_504 
* INOUT : bl_505 
* INOUT : br_505 
* INOUT : bl_506 
* INOUT : br_506 
* INOUT : bl_507 
* INOUT : br_507 
* INOUT : bl_508 
* INOUT : br_508 
* INOUT : bl_509 
* INOUT : br_509 
* INOUT : bl_510 
* INOUT : br_510 
* INOUT : bl_511 
* INOUT : br_511 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* OUTPUT: dout_33 
* OUTPUT: dout_34 
* OUTPUT: dout_35 
* OUTPUT: dout_36 
* OUTPUT: dout_37 
* OUTPUT: dout_38 
* OUTPUT: dout_39 
* OUTPUT: dout_40 
* OUTPUT: dout_41 
* OUTPUT: dout_42 
* OUTPUT: dout_43 
* OUTPUT: dout_44 
* OUTPUT: dout_45 
* OUTPUT: dout_46 
* OUTPUT: dout_47 
* OUTPUT: dout_48 
* OUTPUT: dout_49 
* OUTPUT: dout_50 
* OUTPUT: dout_51 
* OUTPUT: dout_52 
* OUTPUT: dout_53 
* OUTPUT: dout_54 
* OUTPUT: dout_55 
* OUTPUT: dout_56 
* OUTPUT: dout_57 
* OUTPUT: dout_58 
* OUTPUT: dout_59 
* OUTPUT: dout_60 
* OUTPUT: dout_61 
* OUTPUT: dout_62 
* OUTPUT: dout_63 
* OUTPUT: dout_64 
* OUTPUT: dout_65 
* OUTPUT: dout_66 
* OUTPUT: dout_67 
* OUTPUT: dout_68 
* OUTPUT: dout_69 
* OUTPUT: dout_70 
* OUTPUT: dout_71 
* OUTPUT: dout_72 
* OUTPUT: dout_73 
* OUTPUT: dout_74 
* OUTPUT: dout_75 
* OUTPUT: dout_76 
* OUTPUT: dout_77 
* OUTPUT: dout_78 
* OUTPUT: dout_79 
* OUTPUT: dout_80 
* OUTPUT: dout_81 
* OUTPUT: dout_82 
* OUTPUT: dout_83 
* OUTPUT: dout_84 
* OUTPUT: dout_85 
* OUTPUT: dout_86 
* OUTPUT: dout_87 
* OUTPUT: dout_88 
* OUTPUT: dout_89 
* OUTPUT: dout_90 
* OUTPUT: dout_91 
* OUTPUT: dout_92 
* OUTPUT: dout_93 
* OUTPUT: dout_94 
* OUTPUT: dout_95 
* OUTPUT: dout_96 
* OUTPUT: dout_97 
* OUTPUT: dout_98 
* OUTPUT: dout_99 
* OUTPUT: dout_100 
* OUTPUT: dout_101 
* OUTPUT: dout_102 
* OUTPUT: dout_103 
* OUTPUT: dout_104 
* OUTPUT: dout_105 
* OUTPUT: dout_106 
* OUTPUT: dout_107 
* OUTPUT: dout_108 
* OUTPUT: dout_109 
* OUTPUT: dout_110 
* OUTPUT: dout_111 
* OUTPUT: dout_112 
* OUTPUT: dout_113 
* OUTPUT: dout_114 
* OUTPUT: dout_115 
* OUTPUT: dout_116 
* OUTPUT: dout_117 
* OUTPUT: dout_118 
* OUTPUT: dout_119 
* OUTPUT: dout_120 
* OUTPUT: dout_121 
* OUTPUT: dout_122 
* OUTPUT: dout_123 
* OUTPUT: dout_124 
* OUTPUT: dout_125 
* OUTPUT: dout_126 
* OUTPUT: dout_127 
* OUTPUT: dout_128 
* OUTPUT: dout_129 
* OUTPUT: dout_130 
* OUTPUT: dout_131 
* OUTPUT: dout_132 
* OUTPUT: dout_133 
* OUTPUT: dout_134 
* OUTPUT: dout_135 
* OUTPUT: dout_136 
* OUTPUT: dout_137 
* OUTPUT: dout_138 
* OUTPUT: dout_139 
* OUTPUT: dout_140 
* OUTPUT: dout_141 
* OUTPUT: dout_142 
* OUTPUT: dout_143 
* OUTPUT: dout_144 
* OUTPUT: dout_145 
* OUTPUT: dout_146 
* OUTPUT: dout_147 
* OUTPUT: dout_148 
* OUTPUT: dout_149 
* OUTPUT: dout_150 
* OUTPUT: dout_151 
* OUTPUT: dout_152 
* OUTPUT: dout_153 
* OUTPUT: dout_154 
* OUTPUT: dout_155 
* OUTPUT: dout_156 
* OUTPUT: dout_157 
* OUTPUT: dout_158 
* OUTPUT: dout_159 
* OUTPUT: dout_160 
* OUTPUT: dout_161 
* OUTPUT: dout_162 
* OUTPUT: dout_163 
* OUTPUT: dout_164 
* OUTPUT: dout_165 
* OUTPUT: dout_166 
* OUTPUT: dout_167 
* OUTPUT: dout_168 
* OUTPUT: dout_169 
* OUTPUT: dout_170 
* OUTPUT: dout_171 
* OUTPUT: dout_172 
* OUTPUT: dout_173 
* OUTPUT: dout_174 
* OUTPUT: dout_175 
* OUTPUT: dout_176 
* OUTPUT: dout_177 
* OUTPUT: dout_178 
* OUTPUT: dout_179 
* OUTPUT: dout_180 
* OUTPUT: dout_181 
* OUTPUT: dout_182 
* OUTPUT: dout_183 
* OUTPUT: dout_184 
* OUTPUT: dout_185 
* OUTPUT: dout_186 
* OUTPUT: dout_187 
* OUTPUT: dout_188 
* OUTPUT: dout_189 
* OUTPUT: dout_190 
* OUTPUT: dout_191 
* OUTPUT: dout_192 
* OUTPUT: dout_193 
* OUTPUT: dout_194 
* OUTPUT: dout_195 
* OUTPUT: dout_196 
* OUTPUT: dout_197 
* OUTPUT: dout_198 
* OUTPUT: dout_199 
* OUTPUT: dout_200 
* OUTPUT: dout_201 
* OUTPUT: dout_202 
* OUTPUT: dout_203 
* OUTPUT: dout_204 
* OUTPUT: dout_205 
* OUTPUT: dout_206 
* OUTPUT: dout_207 
* OUTPUT: dout_208 
* OUTPUT: dout_209 
* OUTPUT: dout_210 
* OUTPUT: dout_211 
* OUTPUT: dout_212 
* OUTPUT: dout_213 
* OUTPUT: dout_214 
* OUTPUT: dout_215 
* OUTPUT: dout_216 
* OUTPUT: dout_217 
* OUTPUT: dout_218 
* OUTPUT: dout_219 
* OUTPUT: dout_220 
* OUTPUT: dout_221 
* OUTPUT: dout_222 
* OUTPUT: dout_223 
* OUTPUT: dout_224 
* OUTPUT: dout_225 
* OUTPUT: dout_226 
* OUTPUT: dout_227 
* OUTPUT: dout_228 
* OUTPUT: dout_229 
* OUTPUT: dout_230 
* OUTPUT: dout_231 
* OUTPUT: dout_232 
* OUTPUT: dout_233 
* OUTPUT: dout_234 
* OUTPUT: dout_235 
* OUTPUT: dout_236 
* OUTPUT: dout_237 
* OUTPUT: dout_238 
* OUTPUT: dout_239 
* OUTPUT: dout_240 
* OUTPUT: dout_241 
* OUTPUT: dout_242 
* OUTPUT: dout_243 
* OUTPUT: dout_244 
* OUTPUT: dout_245 
* OUTPUT: dout_246 
* OUTPUT: dout_247 
* OUTPUT: dout_248 
* OUTPUT: dout_249 
* OUTPUT: dout_250 
* OUTPUT: dout_251 
* OUTPUT: dout_252 
* OUTPUT: dout_253 
* OUTPUT: dout_254 
* OUTPUT: dout_255 
* OUTPUT: dout_256 
* OUTPUT: dout_257 
* OUTPUT: dout_258 
* OUTPUT: dout_259 
* OUTPUT: dout_260 
* OUTPUT: dout_261 
* OUTPUT: dout_262 
* OUTPUT: dout_263 
* OUTPUT: dout_264 
* OUTPUT: dout_265 
* OUTPUT: dout_266 
* OUTPUT: dout_267 
* OUTPUT: dout_268 
* OUTPUT: dout_269 
* OUTPUT: dout_270 
* OUTPUT: dout_271 
* OUTPUT: dout_272 
* OUTPUT: dout_273 
* OUTPUT: dout_274 
* OUTPUT: dout_275 
* OUTPUT: dout_276 
* OUTPUT: dout_277 
* OUTPUT: dout_278 
* OUTPUT: dout_279 
* OUTPUT: dout_280 
* OUTPUT: dout_281 
* OUTPUT: dout_282 
* OUTPUT: dout_283 
* OUTPUT: dout_284 
* OUTPUT: dout_285 
* OUTPUT: dout_286 
* OUTPUT: dout_287 
* OUTPUT: dout_288 
* OUTPUT: dout_289 
* OUTPUT: dout_290 
* OUTPUT: dout_291 
* OUTPUT: dout_292 
* OUTPUT: dout_293 
* OUTPUT: dout_294 
* OUTPUT: dout_295 
* OUTPUT: dout_296 
* OUTPUT: dout_297 
* OUTPUT: dout_298 
* OUTPUT: dout_299 
* OUTPUT: dout_300 
* OUTPUT: dout_301 
* OUTPUT: dout_302 
* OUTPUT: dout_303 
* OUTPUT: dout_304 
* OUTPUT: dout_305 
* OUTPUT: dout_306 
* OUTPUT: dout_307 
* OUTPUT: dout_308 
* OUTPUT: dout_309 
* OUTPUT: dout_310 
* OUTPUT: dout_311 
* OUTPUT: dout_312 
* OUTPUT: dout_313 
* OUTPUT: dout_314 
* OUTPUT: dout_315 
* OUTPUT: dout_316 
* OUTPUT: dout_317 
* OUTPUT: dout_318 
* OUTPUT: dout_319 
* OUTPUT: dout_320 
* OUTPUT: dout_321 
* OUTPUT: dout_322 
* OUTPUT: dout_323 
* OUTPUT: dout_324 
* OUTPUT: dout_325 
* OUTPUT: dout_326 
* OUTPUT: dout_327 
* OUTPUT: dout_328 
* OUTPUT: dout_329 
* OUTPUT: dout_330 
* OUTPUT: dout_331 
* OUTPUT: dout_332 
* OUTPUT: dout_333 
* OUTPUT: dout_334 
* OUTPUT: dout_335 
* OUTPUT: dout_336 
* OUTPUT: dout_337 
* OUTPUT: dout_338 
* OUTPUT: dout_339 
* OUTPUT: dout_340 
* OUTPUT: dout_341 
* OUTPUT: dout_342 
* OUTPUT: dout_343 
* OUTPUT: dout_344 
* OUTPUT: dout_345 
* OUTPUT: dout_346 
* OUTPUT: dout_347 
* OUTPUT: dout_348 
* OUTPUT: dout_349 
* OUTPUT: dout_350 
* OUTPUT: dout_351 
* OUTPUT: dout_352 
* OUTPUT: dout_353 
* OUTPUT: dout_354 
* OUTPUT: dout_355 
* OUTPUT: dout_356 
* OUTPUT: dout_357 
* OUTPUT: dout_358 
* OUTPUT: dout_359 
* OUTPUT: dout_360 
* OUTPUT: dout_361 
* OUTPUT: dout_362 
* OUTPUT: dout_363 
* OUTPUT: dout_364 
* OUTPUT: dout_365 
* OUTPUT: dout_366 
* OUTPUT: dout_367 
* OUTPUT: dout_368 
* OUTPUT: dout_369 
* OUTPUT: dout_370 
* OUTPUT: dout_371 
* OUTPUT: dout_372 
* OUTPUT: dout_373 
* OUTPUT: dout_374 
* OUTPUT: dout_375 
* OUTPUT: dout_376 
* OUTPUT: dout_377 
* OUTPUT: dout_378 
* OUTPUT: dout_379 
* OUTPUT: dout_380 
* OUTPUT: dout_381 
* OUTPUT: dout_382 
* OUTPUT: dout_383 
* OUTPUT: dout_384 
* OUTPUT: dout_385 
* OUTPUT: dout_386 
* OUTPUT: dout_387 
* OUTPUT: dout_388 
* OUTPUT: dout_389 
* OUTPUT: dout_390 
* OUTPUT: dout_391 
* OUTPUT: dout_392 
* OUTPUT: dout_393 
* OUTPUT: dout_394 
* OUTPUT: dout_395 
* OUTPUT: dout_396 
* OUTPUT: dout_397 
* OUTPUT: dout_398 
* OUTPUT: dout_399 
* OUTPUT: dout_400 
* OUTPUT: dout_401 
* OUTPUT: dout_402 
* OUTPUT: dout_403 
* OUTPUT: dout_404 
* OUTPUT: dout_405 
* OUTPUT: dout_406 
* OUTPUT: dout_407 
* OUTPUT: dout_408 
* OUTPUT: dout_409 
* OUTPUT: dout_410 
* OUTPUT: dout_411 
* OUTPUT: dout_412 
* OUTPUT: dout_413 
* OUTPUT: dout_414 
* OUTPUT: dout_415 
* OUTPUT: dout_416 
* OUTPUT: dout_417 
* OUTPUT: dout_418 
* OUTPUT: dout_419 
* OUTPUT: dout_420 
* OUTPUT: dout_421 
* OUTPUT: dout_422 
* OUTPUT: dout_423 
* OUTPUT: dout_424 
* OUTPUT: dout_425 
* OUTPUT: dout_426 
* OUTPUT: dout_427 
* OUTPUT: dout_428 
* OUTPUT: dout_429 
* OUTPUT: dout_430 
* OUTPUT: dout_431 
* OUTPUT: dout_432 
* OUTPUT: dout_433 
* OUTPUT: dout_434 
* OUTPUT: dout_435 
* OUTPUT: dout_436 
* OUTPUT: dout_437 
* OUTPUT: dout_438 
* OUTPUT: dout_439 
* OUTPUT: dout_440 
* OUTPUT: dout_441 
* OUTPUT: dout_442 
* OUTPUT: dout_443 
* OUTPUT: dout_444 
* OUTPUT: dout_445 
* OUTPUT: dout_446 
* OUTPUT: dout_447 
* OUTPUT: dout_448 
* OUTPUT: dout_449 
* OUTPUT: dout_450 
* OUTPUT: dout_451 
* OUTPUT: dout_452 
* OUTPUT: dout_453 
* OUTPUT: dout_454 
* OUTPUT: dout_455 
* OUTPUT: dout_456 
* OUTPUT: dout_457 
* OUTPUT: dout_458 
* OUTPUT: dout_459 
* OUTPUT: dout_460 
* OUTPUT: dout_461 
* OUTPUT: dout_462 
* OUTPUT: dout_463 
* OUTPUT: dout_464 
* OUTPUT: dout_465 
* OUTPUT: dout_466 
* OUTPUT: dout_467 
* OUTPUT: dout_468 
* OUTPUT: dout_469 
* OUTPUT: dout_470 
* OUTPUT: dout_471 
* OUTPUT: dout_472 
* OUTPUT: dout_473 
* OUTPUT: dout_474 
* OUTPUT: dout_475 
* OUTPUT: dout_476 
* OUTPUT: dout_477 
* OUTPUT: dout_478 
* OUTPUT: dout_479 
* OUTPUT: dout_480 
* OUTPUT: dout_481 
* OUTPUT: dout_482 
* OUTPUT: dout_483 
* OUTPUT: dout_484 
* OUTPUT: dout_485 
* OUTPUT: dout_486 
* OUTPUT: dout_487 
* OUTPUT: dout_488 
* OUTPUT: dout_489 
* OUTPUT: dout_490 
* OUTPUT: dout_491 
* OUTPUT: dout_492 
* OUTPUT: dout_493 
* OUTPUT: dout_494 
* OUTPUT: dout_495 
* OUTPUT: dout_496 
* OUTPUT: dout_497 
* OUTPUT: dout_498 
* OUTPUT: dout_499 
* OUTPUT: dout_500 
* OUTPUT: dout_501 
* OUTPUT: dout_502 
* OUTPUT: dout_503 
* OUTPUT: dout_504 
* OUTPUT: dout_505 
* OUTPUT: dout_506 
* OUTPUT: dout_507 
* OUTPUT: dout_508 
* OUTPUT: dout_509 
* OUTPUT: dout_510 
* OUTPUT: dout_511 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : din_33 
* INPUT : din_34 
* INPUT : din_35 
* INPUT : din_36 
* INPUT : din_37 
* INPUT : din_38 
* INPUT : din_39 
* INPUT : din_40 
* INPUT : din_41 
* INPUT : din_42 
* INPUT : din_43 
* INPUT : din_44 
* INPUT : din_45 
* INPUT : din_46 
* INPUT : din_47 
* INPUT : din_48 
* INPUT : din_49 
* INPUT : din_50 
* INPUT : din_51 
* INPUT : din_52 
* INPUT : din_53 
* INPUT : din_54 
* INPUT : din_55 
* INPUT : din_56 
* INPUT : din_57 
* INPUT : din_58 
* INPUT : din_59 
* INPUT : din_60 
* INPUT : din_61 
* INPUT : din_62 
* INPUT : din_63 
* INPUT : din_64 
* INPUT : din_65 
* INPUT : din_66 
* INPUT : din_67 
* INPUT : din_68 
* INPUT : din_69 
* INPUT : din_70 
* INPUT : din_71 
* INPUT : din_72 
* INPUT : din_73 
* INPUT : din_74 
* INPUT : din_75 
* INPUT : din_76 
* INPUT : din_77 
* INPUT : din_78 
* INPUT : din_79 
* INPUT : din_80 
* INPUT : din_81 
* INPUT : din_82 
* INPUT : din_83 
* INPUT : din_84 
* INPUT : din_85 
* INPUT : din_86 
* INPUT : din_87 
* INPUT : din_88 
* INPUT : din_89 
* INPUT : din_90 
* INPUT : din_91 
* INPUT : din_92 
* INPUT : din_93 
* INPUT : din_94 
* INPUT : din_95 
* INPUT : din_96 
* INPUT : din_97 
* INPUT : din_98 
* INPUT : din_99 
* INPUT : din_100 
* INPUT : din_101 
* INPUT : din_102 
* INPUT : din_103 
* INPUT : din_104 
* INPUT : din_105 
* INPUT : din_106 
* INPUT : din_107 
* INPUT : din_108 
* INPUT : din_109 
* INPUT : din_110 
* INPUT : din_111 
* INPUT : din_112 
* INPUT : din_113 
* INPUT : din_114 
* INPUT : din_115 
* INPUT : din_116 
* INPUT : din_117 
* INPUT : din_118 
* INPUT : din_119 
* INPUT : din_120 
* INPUT : din_121 
* INPUT : din_122 
* INPUT : din_123 
* INPUT : din_124 
* INPUT : din_125 
* INPUT : din_126 
* INPUT : din_127 
* INPUT : din_128 
* INPUT : din_129 
* INPUT : din_130 
* INPUT : din_131 
* INPUT : din_132 
* INPUT : din_133 
* INPUT : din_134 
* INPUT : din_135 
* INPUT : din_136 
* INPUT : din_137 
* INPUT : din_138 
* INPUT : din_139 
* INPUT : din_140 
* INPUT : din_141 
* INPUT : din_142 
* INPUT : din_143 
* INPUT : din_144 
* INPUT : din_145 
* INPUT : din_146 
* INPUT : din_147 
* INPUT : din_148 
* INPUT : din_149 
* INPUT : din_150 
* INPUT : din_151 
* INPUT : din_152 
* INPUT : din_153 
* INPUT : din_154 
* INPUT : din_155 
* INPUT : din_156 
* INPUT : din_157 
* INPUT : din_158 
* INPUT : din_159 
* INPUT : din_160 
* INPUT : din_161 
* INPUT : din_162 
* INPUT : din_163 
* INPUT : din_164 
* INPUT : din_165 
* INPUT : din_166 
* INPUT : din_167 
* INPUT : din_168 
* INPUT : din_169 
* INPUT : din_170 
* INPUT : din_171 
* INPUT : din_172 
* INPUT : din_173 
* INPUT : din_174 
* INPUT : din_175 
* INPUT : din_176 
* INPUT : din_177 
* INPUT : din_178 
* INPUT : din_179 
* INPUT : din_180 
* INPUT : din_181 
* INPUT : din_182 
* INPUT : din_183 
* INPUT : din_184 
* INPUT : din_185 
* INPUT : din_186 
* INPUT : din_187 
* INPUT : din_188 
* INPUT : din_189 
* INPUT : din_190 
* INPUT : din_191 
* INPUT : din_192 
* INPUT : din_193 
* INPUT : din_194 
* INPUT : din_195 
* INPUT : din_196 
* INPUT : din_197 
* INPUT : din_198 
* INPUT : din_199 
* INPUT : din_200 
* INPUT : din_201 
* INPUT : din_202 
* INPUT : din_203 
* INPUT : din_204 
* INPUT : din_205 
* INPUT : din_206 
* INPUT : din_207 
* INPUT : din_208 
* INPUT : din_209 
* INPUT : din_210 
* INPUT : din_211 
* INPUT : din_212 
* INPUT : din_213 
* INPUT : din_214 
* INPUT : din_215 
* INPUT : din_216 
* INPUT : din_217 
* INPUT : din_218 
* INPUT : din_219 
* INPUT : din_220 
* INPUT : din_221 
* INPUT : din_222 
* INPUT : din_223 
* INPUT : din_224 
* INPUT : din_225 
* INPUT : din_226 
* INPUT : din_227 
* INPUT : din_228 
* INPUT : din_229 
* INPUT : din_230 
* INPUT : din_231 
* INPUT : din_232 
* INPUT : din_233 
* INPUT : din_234 
* INPUT : din_235 
* INPUT : din_236 
* INPUT : din_237 
* INPUT : din_238 
* INPUT : din_239 
* INPUT : din_240 
* INPUT : din_241 
* INPUT : din_242 
* INPUT : din_243 
* INPUT : din_244 
* INPUT : din_245 
* INPUT : din_246 
* INPUT : din_247 
* INPUT : din_248 
* INPUT : din_249 
* INPUT : din_250 
* INPUT : din_251 
* INPUT : din_252 
* INPUT : din_253 
* INPUT : din_254 
* INPUT : din_255 
* INPUT : din_256 
* INPUT : din_257 
* INPUT : din_258 
* INPUT : din_259 
* INPUT : din_260 
* INPUT : din_261 
* INPUT : din_262 
* INPUT : din_263 
* INPUT : din_264 
* INPUT : din_265 
* INPUT : din_266 
* INPUT : din_267 
* INPUT : din_268 
* INPUT : din_269 
* INPUT : din_270 
* INPUT : din_271 
* INPUT : din_272 
* INPUT : din_273 
* INPUT : din_274 
* INPUT : din_275 
* INPUT : din_276 
* INPUT : din_277 
* INPUT : din_278 
* INPUT : din_279 
* INPUT : din_280 
* INPUT : din_281 
* INPUT : din_282 
* INPUT : din_283 
* INPUT : din_284 
* INPUT : din_285 
* INPUT : din_286 
* INPUT : din_287 
* INPUT : din_288 
* INPUT : din_289 
* INPUT : din_290 
* INPUT : din_291 
* INPUT : din_292 
* INPUT : din_293 
* INPUT : din_294 
* INPUT : din_295 
* INPUT : din_296 
* INPUT : din_297 
* INPUT : din_298 
* INPUT : din_299 
* INPUT : din_300 
* INPUT : din_301 
* INPUT : din_302 
* INPUT : din_303 
* INPUT : din_304 
* INPUT : din_305 
* INPUT : din_306 
* INPUT : din_307 
* INPUT : din_308 
* INPUT : din_309 
* INPUT : din_310 
* INPUT : din_311 
* INPUT : din_312 
* INPUT : din_313 
* INPUT : din_314 
* INPUT : din_315 
* INPUT : din_316 
* INPUT : din_317 
* INPUT : din_318 
* INPUT : din_319 
* INPUT : din_320 
* INPUT : din_321 
* INPUT : din_322 
* INPUT : din_323 
* INPUT : din_324 
* INPUT : din_325 
* INPUT : din_326 
* INPUT : din_327 
* INPUT : din_328 
* INPUT : din_329 
* INPUT : din_330 
* INPUT : din_331 
* INPUT : din_332 
* INPUT : din_333 
* INPUT : din_334 
* INPUT : din_335 
* INPUT : din_336 
* INPUT : din_337 
* INPUT : din_338 
* INPUT : din_339 
* INPUT : din_340 
* INPUT : din_341 
* INPUT : din_342 
* INPUT : din_343 
* INPUT : din_344 
* INPUT : din_345 
* INPUT : din_346 
* INPUT : din_347 
* INPUT : din_348 
* INPUT : din_349 
* INPUT : din_350 
* INPUT : din_351 
* INPUT : din_352 
* INPUT : din_353 
* INPUT : din_354 
* INPUT : din_355 
* INPUT : din_356 
* INPUT : din_357 
* INPUT : din_358 
* INPUT : din_359 
* INPUT : din_360 
* INPUT : din_361 
* INPUT : din_362 
* INPUT : din_363 
* INPUT : din_364 
* INPUT : din_365 
* INPUT : din_366 
* INPUT : din_367 
* INPUT : din_368 
* INPUT : din_369 
* INPUT : din_370 
* INPUT : din_371 
* INPUT : din_372 
* INPUT : din_373 
* INPUT : din_374 
* INPUT : din_375 
* INPUT : din_376 
* INPUT : din_377 
* INPUT : din_378 
* INPUT : din_379 
* INPUT : din_380 
* INPUT : din_381 
* INPUT : din_382 
* INPUT : din_383 
* INPUT : din_384 
* INPUT : din_385 
* INPUT : din_386 
* INPUT : din_387 
* INPUT : din_388 
* INPUT : din_389 
* INPUT : din_390 
* INPUT : din_391 
* INPUT : din_392 
* INPUT : din_393 
* INPUT : din_394 
* INPUT : din_395 
* INPUT : din_396 
* INPUT : din_397 
* INPUT : din_398 
* INPUT : din_399 
* INPUT : din_400 
* INPUT : din_401 
* INPUT : din_402 
* INPUT : din_403 
* INPUT : din_404 
* INPUT : din_405 
* INPUT : din_406 
* INPUT : din_407 
* INPUT : din_408 
* INPUT : din_409 
* INPUT : din_410 
* INPUT : din_411 
* INPUT : din_412 
* INPUT : din_413 
* INPUT : din_414 
* INPUT : din_415 
* INPUT : din_416 
* INPUT : din_417 
* INPUT : din_418 
* INPUT : din_419 
* INPUT : din_420 
* INPUT : din_421 
* INPUT : din_422 
* INPUT : din_423 
* INPUT : din_424 
* INPUT : din_425 
* INPUT : din_426 
* INPUT : din_427 
* INPUT : din_428 
* INPUT : din_429 
* INPUT : din_430 
* INPUT : din_431 
* INPUT : din_432 
* INPUT : din_433 
* INPUT : din_434 
* INPUT : din_435 
* INPUT : din_436 
* INPUT : din_437 
* INPUT : din_438 
* INPUT : din_439 
* INPUT : din_440 
* INPUT : din_441 
* INPUT : din_442 
* INPUT : din_443 
* INPUT : din_444 
* INPUT : din_445 
* INPUT : din_446 
* INPUT : din_447 
* INPUT : din_448 
* INPUT : din_449 
* INPUT : din_450 
* INPUT : din_451 
* INPUT : din_452 
* INPUT : din_453 
* INPUT : din_454 
* INPUT : din_455 
* INPUT : din_456 
* INPUT : din_457 
* INPUT : din_458 
* INPUT : din_459 
* INPUT : din_460 
* INPUT : din_461 
* INPUT : din_462 
* INPUT : din_463 
* INPUT : din_464 
* INPUT : din_465 
* INPUT : din_466 
* INPUT : din_467 
* INPUT : din_468 
* INPUT : din_469 
* INPUT : din_470 
* INPUT : din_471 
* INPUT : din_472 
* INPUT : din_473 
* INPUT : din_474 
* INPUT : din_475 
* INPUT : din_476 
* INPUT : din_477 
* INPUT : din_478 
* INPUT : din_479 
* INPUT : din_480 
* INPUT : din_481 
* INPUT : din_482 
* INPUT : din_483 
* INPUT : din_484 
* INPUT : din_485 
* INPUT : din_486 
* INPUT : din_487 
* INPUT : din_488 
* INPUT : din_489 
* INPUT : din_490 
* INPUT : din_491 
* INPUT : din_492 
* INPUT : din_493 
* INPUT : din_494 
* INPUT : din_495 
* INPUT : din_496 
* INPUT : din_497 
* INPUT : din_498 
* INPUT : din_499 
* INPUT : din_500 
* INPUT : din_501 
* INPUT : din_502 
* INPUT : din_503 
* INPUT : din_504 
* INPUT : din_505 
* INPUT : din_506 
* INPUT : din_507 
* INPUT : din_508 
* INPUT : din_509 
* INPUT : din_510 
* INPUT : din_511 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66
+ bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72
+ br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77
+ bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83
+ br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88
+ bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94
+ br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99
+ bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104
+ bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109
+ bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114
+ bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119
+ bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124
+ bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129
+ bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134
+ bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139
+ bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144
+ bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149
+ bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154
+ bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159
+ bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164
+ bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169
+ bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174
+ bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179
+ bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184
+ bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189
+ bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194
+ bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199
+ bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204
+ bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209
+ bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214
+ bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219
+ bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224
+ bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229
+ bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234
+ bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239
+ bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244
+ bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249
+ bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254
+ bl_255 br_255 bl_256 br_256 bl_257 br_257 bl_258 br_258 bl_259 br_259
+ bl_260 br_260 bl_261 br_261 bl_262 br_262 bl_263 br_263 bl_264 br_264
+ bl_265 br_265 bl_266 br_266 bl_267 br_267 bl_268 br_268 bl_269 br_269
+ bl_270 br_270 bl_271 br_271 bl_272 br_272 bl_273 br_273 bl_274 br_274
+ bl_275 br_275 bl_276 br_276 bl_277 br_277 bl_278 br_278 bl_279 br_279
+ bl_280 br_280 bl_281 br_281 bl_282 br_282 bl_283 br_283 bl_284 br_284
+ bl_285 br_285 bl_286 br_286 bl_287 br_287 bl_288 br_288 bl_289 br_289
+ bl_290 br_290 bl_291 br_291 bl_292 br_292 bl_293 br_293 bl_294 br_294
+ bl_295 br_295 bl_296 br_296 bl_297 br_297 bl_298 br_298 bl_299 br_299
+ bl_300 br_300 bl_301 br_301 bl_302 br_302 bl_303 br_303 bl_304 br_304
+ bl_305 br_305 bl_306 br_306 bl_307 br_307 bl_308 br_308 bl_309 br_309
+ bl_310 br_310 bl_311 br_311 bl_312 br_312 bl_313 br_313 bl_314 br_314
+ bl_315 br_315 bl_316 br_316 bl_317 br_317 bl_318 br_318 bl_319 br_319
+ bl_320 br_320 bl_321 br_321 bl_322 br_322 bl_323 br_323 bl_324 br_324
+ bl_325 br_325 bl_326 br_326 bl_327 br_327 bl_328 br_328 bl_329 br_329
+ bl_330 br_330 bl_331 br_331 bl_332 br_332 bl_333 br_333 bl_334 br_334
+ bl_335 br_335 bl_336 br_336 bl_337 br_337 bl_338 br_338 bl_339 br_339
+ bl_340 br_340 bl_341 br_341 bl_342 br_342 bl_343 br_343 bl_344 br_344
+ bl_345 br_345 bl_346 br_346 bl_347 br_347 bl_348 br_348 bl_349 br_349
+ bl_350 br_350 bl_351 br_351 bl_352 br_352 bl_353 br_353 bl_354 br_354
+ bl_355 br_355 bl_356 br_356 bl_357 br_357 bl_358 br_358 bl_359 br_359
+ bl_360 br_360 bl_361 br_361 bl_362 br_362 bl_363 br_363 bl_364 br_364
+ bl_365 br_365 bl_366 br_366 bl_367 br_367 bl_368 br_368 bl_369 br_369
+ bl_370 br_370 bl_371 br_371 bl_372 br_372 bl_373 br_373 bl_374 br_374
+ bl_375 br_375 bl_376 br_376 bl_377 br_377 bl_378 br_378 bl_379 br_379
+ bl_380 br_380 bl_381 br_381 bl_382 br_382 bl_383 br_383 bl_384 br_384
+ bl_385 br_385 bl_386 br_386 bl_387 br_387 bl_388 br_388 bl_389 br_389
+ bl_390 br_390 bl_391 br_391 bl_392 br_392 bl_393 br_393 bl_394 br_394
+ bl_395 br_395 bl_396 br_396 bl_397 br_397 bl_398 br_398 bl_399 br_399
+ bl_400 br_400 bl_401 br_401 bl_402 br_402 bl_403 br_403 bl_404 br_404
+ bl_405 br_405 bl_406 br_406 bl_407 br_407 bl_408 br_408 bl_409 br_409
+ bl_410 br_410 bl_411 br_411 bl_412 br_412 bl_413 br_413 bl_414 br_414
+ bl_415 br_415 bl_416 br_416 bl_417 br_417 bl_418 br_418 bl_419 br_419
+ bl_420 br_420 bl_421 br_421 bl_422 br_422 bl_423 br_423 bl_424 br_424
+ bl_425 br_425 bl_426 br_426 bl_427 br_427 bl_428 br_428 bl_429 br_429
+ bl_430 br_430 bl_431 br_431 bl_432 br_432 bl_433 br_433 bl_434 br_434
+ bl_435 br_435 bl_436 br_436 bl_437 br_437 bl_438 br_438 bl_439 br_439
+ bl_440 br_440 bl_441 br_441 bl_442 br_442 bl_443 br_443 bl_444 br_444
+ bl_445 br_445 bl_446 br_446 bl_447 br_447 bl_448 br_448 bl_449 br_449
+ bl_450 br_450 bl_451 br_451 bl_452 br_452 bl_453 br_453 bl_454 br_454
+ bl_455 br_455 bl_456 br_456 bl_457 br_457 bl_458 br_458 bl_459 br_459
+ bl_460 br_460 bl_461 br_461 bl_462 br_462 bl_463 br_463 bl_464 br_464
+ bl_465 br_465 bl_466 br_466 bl_467 br_467 bl_468 br_468 bl_469 br_469
+ bl_470 br_470 bl_471 br_471 bl_472 br_472 bl_473 br_473 bl_474 br_474
+ bl_475 br_475 bl_476 br_476 bl_477 br_477 bl_478 br_478 bl_479 br_479
+ bl_480 br_480 bl_481 br_481 bl_482 br_482 bl_483 br_483 bl_484 br_484
+ bl_485 br_485 bl_486 br_486 bl_487 br_487 bl_488 br_488 bl_489 br_489
+ bl_490 br_490 bl_491 br_491 bl_492 br_492 bl_493 br_493 bl_494 br_494
+ bl_495 br_495 bl_496 br_496 bl_497 br_497 bl_498 br_498 bl_499 br_499
+ bl_500 br_500 bl_501 br_501 bl_502 br_502 bl_503 br_503 bl_504 br_504
+ bl_505 br_505 bl_506 br_506 bl_507 br_507 bl_508 br_508 bl_509 br_509
+ bl_510 br_510 bl_511 br_511 p_en_bar vdd
+ freepdk45_sram_1rw0r_45x512_precharge_array
Xsense_amp_array0
+ dout_0 bl_0 br_0 dout_1 bl_1 br_1 dout_2 bl_2 br_2 dout_3 bl_3 br_3
+ dout_4 bl_4 br_4 dout_5 bl_5 br_5 dout_6 bl_6 br_6 dout_7 bl_7 br_7
+ dout_8 bl_8 br_8 dout_9 bl_9 br_9 dout_10 bl_10 br_10 dout_11 bl_11
+ br_11 dout_12 bl_12 br_12 dout_13 bl_13 br_13 dout_14 bl_14 br_14
+ dout_15 bl_15 br_15 dout_16 bl_16 br_16 dout_17 bl_17 br_17 dout_18
+ bl_18 br_18 dout_19 bl_19 br_19 dout_20 bl_20 br_20 dout_21 bl_21
+ br_21 dout_22 bl_22 br_22 dout_23 bl_23 br_23 dout_24 bl_24 br_24
+ dout_25 bl_25 br_25 dout_26 bl_26 br_26 dout_27 bl_27 br_27 dout_28
+ bl_28 br_28 dout_29 bl_29 br_29 dout_30 bl_30 br_30 dout_31 bl_31
+ br_31 dout_32 bl_32 br_32 dout_33 bl_33 br_33 dout_34 bl_34 br_34
+ dout_35 bl_35 br_35 dout_36 bl_36 br_36 dout_37 bl_37 br_37 dout_38
+ bl_38 br_38 dout_39 bl_39 br_39 dout_40 bl_40 br_40 dout_41 bl_41
+ br_41 dout_42 bl_42 br_42 dout_43 bl_43 br_43 dout_44 bl_44 br_44
+ dout_45 bl_45 br_45 dout_46 bl_46 br_46 dout_47 bl_47 br_47 dout_48
+ bl_48 br_48 dout_49 bl_49 br_49 dout_50 bl_50 br_50 dout_51 bl_51
+ br_51 dout_52 bl_52 br_52 dout_53 bl_53 br_53 dout_54 bl_54 br_54
+ dout_55 bl_55 br_55 dout_56 bl_56 br_56 dout_57 bl_57 br_57 dout_58
+ bl_58 br_58 dout_59 bl_59 br_59 dout_60 bl_60 br_60 dout_61 bl_61
+ br_61 dout_62 bl_62 br_62 dout_63 bl_63 br_63 dout_64 bl_64 br_64
+ dout_65 bl_65 br_65 dout_66 bl_66 br_66 dout_67 bl_67 br_67 dout_68
+ bl_68 br_68 dout_69 bl_69 br_69 dout_70 bl_70 br_70 dout_71 bl_71
+ br_71 dout_72 bl_72 br_72 dout_73 bl_73 br_73 dout_74 bl_74 br_74
+ dout_75 bl_75 br_75 dout_76 bl_76 br_76 dout_77 bl_77 br_77 dout_78
+ bl_78 br_78 dout_79 bl_79 br_79 dout_80 bl_80 br_80 dout_81 bl_81
+ br_81 dout_82 bl_82 br_82 dout_83 bl_83 br_83 dout_84 bl_84 br_84
+ dout_85 bl_85 br_85 dout_86 bl_86 br_86 dout_87 bl_87 br_87 dout_88
+ bl_88 br_88 dout_89 bl_89 br_89 dout_90 bl_90 br_90 dout_91 bl_91
+ br_91 dout_92 bl_92 br_92 dout_93 bl_93 br_93 dout_94 bl_94 br_94
+ dout_95 bl_95 br_95 dout_96 bl_96 br_96 dout_97 bl_97 br_97 dout_98
+ bl_98 br_98 dout_99 bl_99 br_99 dout_100 bl_100 br_100 dout_101 bl_101
+ br_101 dout_102 bl_102 br_102 dout_103 bl_103 br_103 dout_104 bl_104
+ br_104 dout_105 bl_105 br_105 dout_106 bl_106 br_106 dout_107 bl_107
+ br_107 dout_108 bl_108 br_108 dout_109 bl_109 br_109 dout_110 bl_110
+ br_110 dout_111 bl_111 br_111 dout_112 bl_112 br_112 dout_113 bl_113
+ br_113 dout_114 bl_114 br_114 dout_115 bl_115 br_115 dout_116 bl_116
+ br_116 dout_117 bl_117 br_117 dout_118 bl_118 br_118 dout_119 bl_119
+ br_119 dout_120 bl_120 br_120 dout_121 bl_121 br_121 dout_122 bl_122
+ br_122 dout_123 bl_123 br_123 dout_124 bl_124 br_124 dout_125 bl_125
+ br_125 dout_126 bl_126 br_126 dout_127 bl_127 br_127 dout_128 bl_128
+ br_128 dout_129 bl_129 br_129 dout_130 bl_130 br_130 dout_131 bl_131
+ br_131 dout_132 bl_132 br_132 dout_133 bl_133 br_133 dout_134 bl_134
+ br_134 dout_135 bl_135 br_135 dout_136 bl_136 br_136 dout_137 bl_137
+ br_137 dout_138 bl_138 br_138 dout_139 bl_139 br_139 dout_140 bl_140
+ br_140 dout_141 bl_141 br_141 dout_142 bl_142 br_142 dout_143 bl_143
+ br_143 dout_144 bl_144 br_144 dout_145 bl_145 br_145 dout_146 bl_146
+ br_146 dout_147 bl_147 br_147 dout_148 bl_148 br_148 dout_149 bl_149
+ br_149 dout_150 bl_150 br_150 dout_151 bl_151 br_151 dout_152 bl_152
+ br_152 dout_153 bl_153 br_153 dout_154 bl_154 br_154 dout_155 bl_155
+ br_155 dout_156 bl_156 br_156 dout_157 bl_157 br_157 dout_158 bl_158
+ br_158 dout_159 bl_159 br_159 dout_160 bl_160 br_160 dout_161 bl_161
+ br_161 dout_162 bl_162 br_162 dout_163 bl_163 br_163 dout_164 bl_164
+ br_164 dout_165 bl_165 br_165 dout_166 bl_166 br_166 dout_167 bl_167
+ br_167 dout_168 bl_168 br_168 dout_169 bl_169 br_169 dout_170 bl_170
+ br_170 dout_171 bl_171 br_171 dout_172 bl_172 br_172 dout_173 bl_173
+ br_173 dout_174 bl_174 br_174 dout_175 bl_175 br_175 dout_176 bl_176
+ br_176 dout_177 bl_177 br_177 dout_178 bl_178 br_178 dout_179 bl_179
+ br_179 dout_180 bl_180 br_180 dout_181 bl_181 br_181 dout_182 bl_182
+ br_182 dout_183 bl_183 br_183 dout_184 bl_184 br_184 dout_185 bl_185
+ br_185 dout_186 bl_186 br_186 dout_187 bl_187 br_187 dout_188 bl_188
+ br_188 dout_189 bl_189 br_189 dout_190 bl_190 br_190 dout_191 bl_191
+ br_191 dout_192 bl_192 br_192 dout_193 bl_193 br_193 dout_194 bl_194
+ br_194 dout_195 bl_195 br_195 dout_196 bl_196 br_196 dout_197 bl_197
+ br_197 dout_198 bl_198 br_198 dout_199 bl_199 br_199 dout_200 bl_200
+ br_200 dout_201 bl_201 br_201 dout_202 bl_202 br_202 dout_203 bl_203
+ br_203 dout_204 bl_204 br_204 dout_205 bl_205 br_205 dout_206 bl_206
+ br_206 dout_207 bl_207 br_207 dout_208 bl_208 br_208 dout_209 bl_209
+ br_209 dout_210 bl_210 br_210 dout_211 bl_211 br_211 dout_212 bl_212
+ br_212 dout_213 bl_213 br_213 dout_214 bl_214 br_214 dout_215 bl_215
+ br_215 dout_216 bl_216 br_216 dout_217 bl_217 br_217 dout_218 bl_218
+ br_218 dout_219 bl_219 br_219 dout_220 bl_220 br_220 dout_221 bl_221
+ br_221 dout_222 bl_222 br_222 dout_223 bl_223 br_223 dout_224 bl_224
+ br_224 dout_225 bl_225 br_225 dout_226 bl_226 br_226 dout_227 bl_227
+ br_227 dout_228 bl_228 br_228 dout_229 bl_229 br_229 dout_230 bl_230
+ br_230 dout_231 bl_231 br_231 dout_232 bl_232 br_232 dout_233 bl_233
+ br_233 dout_234 bl_234 br_234 dout_235 bl_235 br_235 dout_236 bl_236
+ br_236 dout_237 bl_237 br_237 dout_238 bl_238 br_238 dout_239 bl_239
+ br_239 dout_240 bl_240 br_240 dout_241 bl_241 br_241 dout_242 bl_242
+ br_242 dout_243 bl_243 br_243 dout_244 bl_244 br_244 dout_245 bl_245
+ br_245 dout_246 bl_246 br_246 dout_247 bl_247 br_247 dout_248 bl_248
+ br_248 dout_249 bl_249 br_249 dout_250 bl_250 br_250 dout_251 bl_251
+ br_251 dout_252 bl_252 br_252 dout_253 bl_253 br_253 dout_254 bl_254
+ br_254 dout_255 bl_255 br_255 dout_256 bl_256 br_256 dout_257 bl_257
+ br_257 dout_258 bl_258 br_258 dout_259 bl_259 br_259 dout_260 bl_260
+ br_260 dout_261 bl_261 br_261 dout_262 bl_262 br_262 dout_263 bl_263
+ br_263 dout_264 bl_264 br_264 dout_265 bl_265 br_265 dout_266 bl_266
+ br_266 dout_267 bl_267 br_267 dout_268 bl_268 br_268 dout_269 bl_269
+ br_269 dout_270 bl_270 br_270 dout_271 bl_271 br_271 dout_272 bl_272
+ br_272 dout_273 bl_273 br_273 dout_274 bl_274 br_274 dout_275 bl_275
+ br_275 dout_276 bl_276 br_276 dout_277 bl_277 br_277 dout_278 bl_278
+ br_278 dout_279 bl_279 br_279 dout_280 bl_280 br_280 dout_281 bl_281
+ br_281 dout_282 bl_282 br_282 dout_283 bl_283 br_283 dout_284 bl_284
+ br_284 dout_285 bl_285 br_285 dout_286 bl_286 br_286 dout_287 bl_287
+ br_287 dout_288 bl_288 br_288 dout_289 bl_289 br_289 dout_290 bl_290
+ br_290 dout_291 bl_291 br_291 dout_292 bl_292 br_292 dout_293 bl_293
+ br_293 dout_294 bl_294 br_294 dout_295 bl_295 br_295 dout_296 bl_296
+ br_296 dout_297 bl_297 br_297 dout_298 bl_298 br_298 dout_299 bl_299
+ br_299 dout_300 bl_300 br_300 dout_301 bl_301 br_301 dout_302 bl_302
+ br_302 dout_303 bl_303 br_303 dout_304 bl_304 br_304 dout_305 bl_305
+ br_305 dout_306 bl_306 br_306 dout_307 bl_307 br_307 dout_308 bl_308
+ br_308 dout_309 bl_309 br_309 dout_310 bl_310 br_310 dout_311 bl_311
+ br_311 dout_312 bl_312 br_312 dout_313 bl_313 br_313 dout_314 bl_314
+ br_314 dout_315 bl_315 br_315 dout_316 bl_316 br_316 dout_317 bl_317
+ br_317 dout_318 bl_318 br_318 dout_319 bl_319 br_319 dout_320 bl_320
+ br_320 dout_321 bl_321 br_321 dout_322 bl_322 br_322 dout_323 bl_323
+ br_323 dout_324 bl_324 br_324 dout_325 bl_325 br_325 dout_326 bl_326
+ br_326 dout_327 bl_327 br_327 dout_328 bl_328 br_328 dout_329 bl_329
+ br_329 dout_330 bl_330 br_330 dout_331 bl_331 br_331 dout_332 bl_332
+ br_332 dout_333 bl_333 br_333 dout_334 bl_334 br_334 dout_335 bl_335
+ br_335 dout_336 bl_336 br_336 dout_337 bl_337 br_337 dout_338 bl_338
+ br_338 dout_339 bl_339 br_339 dout_340 bl_340 br_340 dout_341 bl_341
+ br_341 dout_342 bl_342 br_342 dout_343 bl_343 br_343 dout_344 bl_344
+ br_344 dout_345 bl_345 br_345 dout_346 bl_346 br_346 dout_347 bl_347
+ br_347 dout_348 bl_348 br_348 dout_349 bl_349 br_349 dout_350 bl_350
+ br_350 dout_351 bl_351 br_351 dout_352 bl_352 br_352 dout_353 bl_353
+ br_353 dout_354 bl_354 br_354 dout_355 bl_355 br_355 dout_356 bl_356
+ br_356 dout_357 bl_357 br_357 dout_358 bl_358 br_358 dout_359 bl_359
+ br_359 dout_360 bl_360 br_360 dout_361 bl_361 br_361 dout_362 bl_362
+ br_362 dout_363 bl_363 br_363 dout_364 bl_364 br_364 dout_365 bl_365
+ br_365 dout_366 bl_366 br_366 dout_367 bl_367 br_367 dout_368 bl_368
+ br_368 dout_369 bl_369 br_369 dout_370 bl_370 br_370 dout_371 bl_371
+ br_371 dout_372 bl_372 br_372 dout_373 bl_373 br_373 dout_374 bl_374
+ br_374 dout_375 bl_375 br_375 dout_376 bl_376 br_376 dout_377 bl_377
+ br_377 dout_378 bl_378 br_378 dout_379 bl_379 br_379 dout_380 bl_380
+ br_380 dout_381 bl_381 br_381 dout_382 bl_382 br_382 dout_383 bl_383
+ br_383 dout_384 bl_384 br_384 dout_385 bl_385 br_385 dout_386 bl_386
+ br_386 dout_387 bl_387 br_387 dout_388 bl_388 br_388 dout_389 bl_389
+ br_389 dout_390 bl_390 br_390 dout_391 bl_391 br_391 dout_392 bl_392
+ br_392 dout_393 bl_393 br_393 dout_394 bl_394 br_394 dout_395 bl_395
+ br_395 dout_396 bl_396 br_396 dout_397 bl_397 br_397 dout_398 bl_398
+ br_398 dout_399 bl_399 br_399 dout_400 bl_400 br_400 dout_401 bl_401
+ br_401 dout_402 bl_402 br_402 dout_403 bl_403 br_403 dout_404 bl_404
+ br_404 dout_405 bl_405 br_405 dout_406 bl_406 br_406 dout_407 bl_407
+ br_407 dout_408 bl_408 br_408 dout_409 bl_409 br_409 dout_410 bl_410
+ br_410 dout_411 bl_411 br_411 dout_412 bl_412 br_412 dout_413 bl_413
+ br_413 dout_414 bl_414 br_414 dout_415 bl_415 br_415 dout_416 bl_416
+ br_416 dout_417 bl_417 br_417 dout_418 bl_418 br_418 dout_419 bl_419
+ br_419 dout_420 bl_420 br_420 dout_421 bl_421 br_421 dout_422 bl_422
+ br_422 dout_423 bl_423 br_423 dout_424 bl_424 br_424 dout_425 bl_425
+ br_425 dout_426 bl_426 br_426 dout_427 bl_427 br_427 dout_428 bl_428
+ br_428 dout_429 bl_429 br_429 dout_430 bl_430 br_430 dout_431 bl_431
+ br_431 dout_432 bl_432 br_432 dout_433 bl_433 br_433 dout_434 bl_434
+ br_434 dout_435 bl_435 br_435 dout_436 bl_436 br_436 dout_437 bl_437
+ br_437 dout_438 bl_438 br_438 dout_439 bl_439 br_439 dout_440 bl_440
+ br_440 dout_441 bl_441 br_441 dout_442 bl_442 br_442 dout_443 bl_443
+ br_443 dout_444 bl_444 br_444 dout_445 bl_445 br_445 dout_446 bl_446
+ br_446 dout_447 bl_447 br_447 dout_448 bl_448 br_448 dout_449 bl_449
+ br_449 dout_450 bl_450 br_450 dout_451 bl_451 br_451 dout_452 bl_452
+ br_452 dout_453 bl_453 br_453 dout_454 bl_454 br_454 dout_455 bl_455
+ br_455 dout_456 bl_456 br_456 dout_457 bl_457 br_457 dout_458 bl_458
+ br_458 dout_459 bl_459 br_459 dout_460 bl_460 br_460 dout_461 bl_461
+ br_461 dout_462 bl_462 br_462 dout_463 bl_463 br_463 dout_464 bl_464
+ br_464 dout_465 bl_465 br_465 dout_466 bl_466 br_466 dout_467 bl_467
+ br_467 dout_468 bl_468 br_468 dout_469 bl_469 br_469 dout_470 bl_470
+ br_470 dout_471 bl_471 br_471 dout_472 bl_472 br_472 dout_473 bl_473
+ br_473 dout_474 bl_474 br_474 dout_475 bl_475 br_475 dout_476 bl_476
+ br_476 dout_477 bl_477 br_477 dout_478 bl_478 br_478 dout_479 bl_479
+ br_479 dout_480 bl_480 br_480 dout_481 bl_481 br_481 dout_482 bl_482
+ br_482 dout_483 bl_483 br_483 dout_484 bl_484 br_484 dout_485 bl_485
+ br_485 dout_486 bl_486 br_486 dout_487 bl_487 br_487 dout_488 bl_488
+ br_488 dout_489 bl_489 br_489 dout_490 bl_490 br_490 dout_491 bl_491
+ br_491 dout_492 bl_492 br_492 dout_493 bl_493 br_493 dout_494 bl_494
+ br_494 dout_495 bl_495 br_495 dout_496 bl_496 br_496 dout_497 bl_497
+ br_497 dout_498 bl_498 br_498 dout_499 bl_499 br_499 dout_500 bl_500
+ br_500 dout_501 bl_501 br_501 dout_502 bl_502 br_502 dout_503 bl_503
+ br_503 dout_504 bl_504 br_504 dout_505 bl_505 br_505 dout_506 bl_506
+ br_506 dout_507 bl_507 br_507 dout_508 bl_508 br_508 dout_509 bl_509
+ br_509 dout_510 bl_510 br_510 dout_511 bl_511 br_511 s_en vdd gnd
+ freepdk45_sram_1rw0r_45x512_sense_amp_array
Xwrite_driver_array0
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10
+ din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20
+ din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30
+ din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40
+ din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50
+ din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60
+ din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70
+ din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80
+ din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90
+ din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100
+ din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108
+ din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116
+ din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124
+ din_125 din_126 din_127 din_128 din_129 din_130 din_131 din_132
+ din_133 din_134 din_135 din_136 din_137 din_138 din_139 din_140
+ din_141 din_142 din_143 din_144 din_145 din_146 din_147 din_148
+ din_149 din_150 din_151 din_152 din_153 din_154 din_155 din_156
+ din_157 din_158 din_159 din_160 din_161 din_162 din_163 din_164
+ din_165 din_166 din_167 din_168 din_169 din_170 din_171 din_172
+ din_173 din_174 din_175 din_176 din_177 din_178 din_179 din_180
+ din_181 din_182 din_183 din_184 din_185 din_186 din_187 din_188
+ din_189 din_190 din_191 din_192 din_193 din_194 din_195 din_196
+ din_197 din_198 din_199 din_200 din_201 din_202 din_203 din_204
+ din_205 din_206 din_207 din_208 din_209 din_210 din_211 din_212
+ din_213 din_214 din_215 din_216 din_217 din_218 din_219 din_220
+ din_221 din_222 din_223 din_224 din_225 din_226 din_227 din_228
+ din_229 din_230 din_231 din_232 din_233 din_234 din_235 din_236
+ din_237 din_238 din_239 din_240 din_241 din_242 din_243 din_244
+ din_245 din_246 din_247 din_248 din_249 din_250 din_251 din_252
+ din_253 din_254 din_255 din_256 din_257 din_258 din_259 din_260
+ din_261 din_262 din_263 din_264 din_265 din_266 din_267 din_268
+ din_269 din_270 din_271 din_272 din_273 din_274 din_275 din_276
+ din_277 din_278 din_279 din_280 din_281 din_282 din_283 din_284
+ din_285 din_286 din_287 din_288 din_289 din_290 din_291 din_292
+ din_293 din_294 din_295 din_296 din_297 din_298 din_299 din_300
+ din_301 din_302 din_303 din_304 din_305 din_306 din_307 din_308
+ din_309 din_310 din_311 din_312 din_313 din_314 din_315 din_316
+ din_317 din_318 din_319 din_320 din_321 din_322 din_323 din_324
+ din_325 din_326 din_327 din_328 din_329 din_330 din_331 din_332
+ din_333 din_334 din_335 din_336 din_337 din_338 din_339 din_340
+ din_341 din_342 din_343 din_344 din_345 din_346 din_347 din_348
+ din_349 din_350 din_351 din_352 din_353 din_354 din_355 din_356
+ din_357 din_358 din_359 din_360 din_361 din_362 din_363 din_364
+ din_365 din_366 din_367 din_368 din_369 din_370 din_371 din_372
+ din_373 din_374 din_375 din_376 din_377 din_378 din_379 din_380
+ din_381 din_382 din_383 din_384 din_385 din_386 din_387 din_388
+ din_389 din_390 din_391 din_392 din_393 din_394 din_395 din_396
+ din_397 din_398 din_399 din_400 din_401 din_402 din_403 din_404
+ din_405 din_406 din_407 din_408 din_409 din_410 din_411 din_412
+ din_413 din_414 din_415 din_416 din_417 din_418 din_419 din_420
+ din_421 din_422 din_423 din_424 din_425 din_426 din_427 din_428
+ din_429 din_430 din_431 din_432 din_433 din_434 din_435 din_436
+ din_437 din_438 din_439 din_440 din_441 din_442 din_443 din_444
+ din_445 din_446 din_447 din_448 din_449 din_450 din_451 din_452
+ din_453 din_454 din_455 din_456 din_457 din_458 din_459 din_460
+ din_461 din_462 din_463 din_464 din_465 din_466 din_467 din_468
+ din_469 din_470 din_471 din_472 din_473 din_474 din_475 din_476
+ din_477 din_478 din_479 din_480 din_481 din_482 din_483 din_484
+ din_485 din_486 din_487 din_488 din_489 din_490 din_491 din_492
+ din_493 din_494 din_495 din_496 din_497 din_498 din_499 din_500
+ din_501 din_502 din_503 din_504 din_505 din_506 din_507 din_508
+ din_509 din_510 din_511 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4
+ br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10
+ bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16
+ br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21
+ bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27
+ br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32
+ bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38
+ br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43
+ bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49
+ br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54
+ bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60
+ br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65
+ bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71
+ br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76
+ bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82
+ br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87
+ bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93
+ br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98
+ bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103
+ bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108
+ bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113
+ bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118
+ bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123
+ bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128
+ bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133
+ bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138
+ bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143
+ bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148
+ bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153
+ bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158
+ bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163
+ bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168
+ bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173
+ bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178
+ bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183
+ bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188
+ bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193
+ bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198
+ bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203
+ bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208
+ bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213
+ bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218
+ bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223
+ bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228
+ bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233
+ bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238
+ bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243
+ bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248
+ bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253
+ bl_254 br_254 bl_255 br_255 bl_256 br_256 bl_257 br_257 bl_258 br_258
+ bl_259 br_259 bl_260 br_260 bl_261 br_261 bl_262 br_262 bl_263 br_263
+ bl_264 br_264 bl_265 br_265 bl_266 br_266 bl_267 br_267 bl_268 br_268
+ bl_269 br_269 bl_270 br_270 bl_271 br_271 bl_272 br_272 bl_273 br_273
+ bl_274 br_274 bl_275 br_275 bl_276 br_276 bl_277 br_277 bl_278 br_278
+ bl_279 br_279 bl_280 br_280 bl_281 br_281 bl_282 br_282 bl_283 br_283
+ bl_284 br_284 bl_285 br_285 bl_286 br_286 bl_287 br_287 bl_288 br_288
+ bl_289 br_289 bl_290 br_290 bl_291 br_291 bl_292 br_292 bl_293 br_293
+ bl_294 br_294 bl_295 br_295 bl_296 br_296 bl_297 br_297 bl_298 br_298
+ bl_299 br_299 bl_300 br_300 bl_301 br_301 bl_302 br_302 bl_303 br_303
+ bl_304 br_304 bl_305 br_305 bl_306 br_306 bl_307 br_307 bl_308 br_308
+ bl_309 br_309 bl_310 br_310 bl_311 br_311 bl_312 br_312 bl_313 br_313
+ bl_314 br_314 bl_315 br_315 bl_316 br_316 bl_317 br_317 bl_318 br_318
+ bl_319 br_319 bl_320 br_320 bl_321 br_321 bl_322 br_322 bl_323 br_323
+ bl_324 br_324 bl_325 br_325 bl_326 br_326 bl_327 br_327 bl_328 br_328
+ bl_329 br_329 bl_330 br_330 bl_331 br_331 bl_332 br_332 bl_333 br_333
+ bl_334 br_334 bl_335 br_335 bl_336 br_336 bl_337 br_337 bl_338 br_338
+ bl_339 br_339 bl_340 br_340 bl_341 br_341 bl_342 br_342 bl_343 br_343
+ bl_344 br_344 bl_345 br_345 bl_346 br_346 bl_347 br_347 bl_348 br_348
+ bl_349 br_349 bl_350 br_350 bl_351 br_351 bl_352 br_352 bl_353 br_353
+ bl_354 br_354 bl_355 br_355 bl_356 br_356 bl_357 br_357 bl_358 br_358
+ bl_359 br_359 bl_360 br_360 bl_361 br_361 bl_362 br_362 bl_363 br_363
+ bl_364 br_364 bl_365 br_365 bl_366 br_366 bl_367 br_367 bl_368 br_368
+ bl_369 br_369 bl_370 br_370 bl_371 br_371 bl_372 br_372 bl_373 br_373
+ bl_374 br_374 bl_375 br_375 bl_376 br_376 bl_377 br_377 bl_378 br_378
+ bl_379 br_379 bl_380 br_380 bl_381 br_381 bl_382 br_382 bl_383 br_383
+ bl_384 br_384 bl_385 br_385 bl_386 br_386 bl_387 br_387 bl_388 br_388
+ bl_389 br_389 bl_390 br_390 bl_391 br_391 bl_392 br_392 bl_393 br_393
+ bl_394 br_394 bl_395 br_395 bl_396 br_396 bl_397 br_397 bl_398 br_398
+ bl_399 br_399 bl_400 br_400 bl_401 br_401 bl_402 br_402 bl_403 br_403
+ bl_404 br_404 bl_405 br_405 bl_406 br_406 bl_407 br_407 bl_408 br_408
+ bl_409 br_409 bl_410 br_410 bl_411 br_411 bl_412 br_412 bl_413 br_413
+ bl_414 br_414 bl_415 br_415 bl_416 br_416 bl_417 br_417 bl_418 br_418
+ bl_419 br_419 bl_420 br_420 bl_421 br_421 bl_422 br_422 bl_423 br_423
+ bl_424 br_424 bl_425 br_425 bl_426 br_426 bl_427 br_427 bl_428 br_428
+ bl_429 br_429 bl_430 br_430 bl_431 br_431 bl_432 br_432 bl_433 br_433
+ bl_434 br_434 bl_435 br_435 bl_436 br_436 bl_437 br_437 bl_438 br_438
+ bl_439 br_439 bl_440 br_440 bl_441 br_441 bl_442 br_442 bl_443 br_443
+ bl_444 br_444 bl_445 br_445 bl_446 br_446 bl_447 br_447 bl_448 br_448
+ bl_449 br_449 bl_450 br_450 bl_451 br_451 bl_452 br_452 bl_453 br_453
+ bl_454 br_454 bl_455 br_455 bl_456 br_456 bl_457 br_457 bl_458 br_458
+ bl_459 br_459 bl_460 br_460 bl_461 br_461 bl_462 br_462 bl_463 br_463
+ bl_464 br_464 bl_465 br_465 bl_466 br_466 bl_467 br_467 bl_468 br_468
+ bl_469 br_469 bl_470 br_470 bl_471 br_471 bl_472 br_472 bl_473 br_473
+ bl_474 br_474 bl_475 br_475 bl_476 br_476 bl_477 br_477 bl_478 br_478
+ bl_479 br_479 bl_480 br_480 bl_481 br_481 bl_482 br_482 bl_483 br_483
+ bl_484 br_484 bl_485 br_485 bl_486 br_486 bl_487 br_487 bl_488 br_488
+ bl_489 br_489 bl_490 br_490 bl_491 br_491 bl_492 br_492 bl_493 br_493
+ bl_494 br_494 bl_495 br_495 bl_496 br_496 bl_497 br_497 bl_498 br_498
+ bl_499 br_499 bl_500 br_500 bl_501 br_501 bl_502 br_502 bl_503 br_503
+ bl_504 br_504 bl_505 br_505 bl_506 br_506 bl_507 br_507 bl_508 br_508
+ bl_509 br_509 bl_510 br_510 bl_511 br_511 w_en vdd gnd
+ freepdk45_sram_1rw0r_45x512_write_driver_array
.ENDS freepdk45_sram_1rw0r_45x512_port_data

.SUBCKT cell_1rw bl br wl vdd gnd
* Inverter 1
MM0 Q_bar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Q_bar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Q_bar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Q_bar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl Q_bar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_1rw


.SUBCKT freepdk45_sram_1rw0r_45x512_bitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258 br_0_258 bl_0_259
+ br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261 bl_0_262 br_0_262
+ bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265 br_0_265 bl_0_266
+ br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268 bl_0_269 br_0_269
+ bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272 br_0_272 bl_0_273
+ br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275 bl_0_276 br_0_276
+ bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279 br_0_279 bl_0_280
+ br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282 bl_0_283 br_0_283
+ bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286 br_0_286 bl_0_287
+ br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289 bl_0_290 br_0_290
+ bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293 br_0_293 bl_0_294
+ br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296 bl_0_297 br_0_297
+ bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300 br_0_300 bl_0_301
+ br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303 bl_0_304 br_0_304
+ bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307 br_0_307 bl_0_308
+ br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310 bl_0_311 br_0_311
+ bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314 br_0_314 bl_0_315
+ br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317 bl_0_318 br_0_318
+ bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321 br_0_321 bl_0_322
+ br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324 bl_0_325 br_0_325
+ bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328 br_0_328 bl_0_329
+ br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331 bl_0_332 br_0_332
+ bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335 br_0_335 bl_0_336
+ br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338 bl_0_339 br_0_339
+ bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342 br_0_342 bl_0_343
+ br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345 bl_0_346 br_0_346
+ bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349 br_0_349 bl_0_350
+ br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352 bl_0_353 br_0_353
+ bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356 br_0_356 bl_0_357
+ br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359 bl_0_360 br_0_360
+ bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363 br_0_363 bl_0_364
+ br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366 bl_0_367 br_0_367
+ bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370 br_0_370 bl_0_371
+ br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373 bl_0_374 br_0_374
+ bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377 br_0_377 bl_0_378
+ br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380 bl_0_381 br_0_381
+ bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384 br_0_384 bl_0_385
+ br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387 bl_0_388 br_0_388
+ bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391 br_0_391 bl_0_392
+ br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394 bl_0_395 br_0_395
+ bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398 br_0_398 bl_0_399
+ br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401 bl_0_402 br_0_402
+ bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405 br_0_405 bl_0_406
+ br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408 bl_0_409 br_0_409
+ bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412 br_0_412 bl_0_413
+ br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415 bl_0_416 br_0_416
+ bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419 br_0_419 bl_0_420
+ br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422 bl_0_423 br_0_423
+ bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426 br_0_426 bl_0_427
+ br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429 bl_0_430 br_0_430
+ bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433 br_0_433 bl_0_434
+ br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436 bl_0_437 br_0_437
+ bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440 br_0_440 bl_0_441
+ br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443 bl_0_444 br_0_444
+ bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447 br_0_447 bl_0_448
+ br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450 bl_0_451 br_0_451
+ bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454 br_0_454 bl_0_455
+ br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457 bl_0_458 br_0_458
+ bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461 br_0_461 bl_0_462
+ br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464 bl_0_465 br_0_465
+ bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468 br_0_468 bl_0_469
+ br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471 bl_0_472 br_0_472
+ bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475 br_0_475 bl_0_476
+ br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478 bl_0_479 br_0_479
+ bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482 br_0_482 bl_0_483
+ br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485 bl_0_486 br_0_486
+ bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489 br_0_489 bl_0_490
+ br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492 bl_0_493 br_0_493
+ bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496 br_0_496 bl_0_497
+ br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499 bl_0_500 br_0_500
+ bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503 br_0_503 bl_0_504
+ br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506 bl_0_507 br_0_507
+ bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510 br_0_510 bl_0_511
+ br_0_511 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INOUT : bl_0_257 
* INOUT : br_0_257 
* INOUT : bl_0_258 
* INOUT : br_0_258 
* INOUT : bl_0_259 
* INOUT : br_0_259 
* INOUT : bl_0_260 
* INOUT : br_0_260 
* INOUT : bl_0_261 
* INOUT : br_0_261 
* INOUT : bl_0_262 
* INOUT : br_0_262 
* INOUT : bl_0_263 
* INOUT : br_0_263 
* INOUT : bl_0_264 
* INOUT : br_0_264 
* INOUT : bl_0_265 
* INOUT : br_0_265 
* INOUT : bl_0_266 
* INOUT : br_0_266 
* INOUT : bl_0_267 
* INOUT : br_0_267 
* INOUT : bl_0_268 
* INOUT : br_0_268 
* INOUT : bl_0_269 
* INOUT : br_0_269 
* INOUT : bl_0_270 
* INOUT : br_0_270 
* INOUT : bl_0_271 
* INOUT : br_0_271 
* INOUT : bl_0_272 
* INOUT : br_0_272 
* INOUT : bl_0_273 
* INOUT : br_0_273 
* INOUT : bl_0_274 
* INOUT : br_0_274 
* INOUT : bl_0_275 
* INOUT : br_0_275 
* INOUT : bl_0_276 
* INOUT : br_0_276 
* INOUT : bl_0_277 
* INOUT : br_0_277 
* INOUT : bl_0_278 
* INOUT : br_0_278 
* INOUT : bl_0_279 
* INOUT : br_0_279 
* INOUT : bl_0_280 
* INOUT : br_0_280 
* INOUT : bl_0_281 
* INOUT : br_0_281 
* INOUT : bl_0_282 
* INOUT : br_0_282 
* INOUT : bl_0_283 
* INOUT : br_0_283 
* INOUT : bl_0_284 
* INOUT : br_0_284 
* INOUT : bl_0_285 
* INOUT : br_0_285 
* INOUT : bl_0_286 
* INOUT : br_0_286 
* INOUT : bl_0_287 
* INOUT : br_0_287 
* INOUT : bl_0_288 
* INOUT : br_0_288 
* INOUT : bl_0_289 
* INOUT : br_0_289 
* INOUT : bl_0_290 
* INOUT : br_0_290 
* INOUT : bl_0_291 
* INOUT : br_0_291 
* INOUT : bl_0_292 
* INOUT : br_0_292 
* INOUT : bl_0_293 
* INOUT : br_0_293 
* INOUT : bl_0_294 
* INOUT : br_0_294 
* INOUT : bl_0_295 
* INOUT : br_0_295 
* INOUT : bl_0_296 
* INOUT : br_0_296 
* INOUT : bl_0_297 
* INOUT : br_0_297 
* INOUT : bl_0_298 
* INOUT : br_0_298 
* INOUT : bl_0_299 
* INOUT : br_0_299 
* INOUT : bl_0_300 
* INOUT : br_0_300 
* INOUT : bl_0_301 
* INOUT : br_0_301 
* INOUT : bl_0_302 
* INOUT : br_0_302 
* INOUT : bl_0_303 
* INOUT : br_0_303 
* INOUT : bl_0_304 
* INOUT : br_0_304 
* INOUT : bl_0_305 
* INOUT : br_0_305 
* INOUT : bl_0_306 
* INOUT : br_0_306 
* INOUT : bl_0_307 
* INOUT : br_0_307 
* INOUT : bl_0_308 
* INOUT : br_0_308 
* INOUT : bl_0_309 
* INOUT : br_0_309 
* INOUT : bl_0_310 
* INOUT : br_0_310 
* INOUT : bl_0_311 
* INOUT : br_0_311 
* INOUT : bl_0_312 
* INOUT : br_0_312 
* INOUT : bl_0_313 
* INOUT : br_0_313 
* INOUT : bl_0_314 
* INOUT : br_0_314 
* INOUT : bl_0_315 
* INOUT : br_0_315 
* INOUT : bl_0_316 
* INOUT : br_0_316 
* INOUT : bl_0_317 
* INOUT : br_0_317 
* INOUT : bl_0_318 
* INOUT : br_0_318 
* INOUT : bl_0_319 
* INOUT : br_0_319 
* INOUT : bl_0_320 
* INOUT : br_0_320 
* INOUT : bl_0_321 
* INOUT : br_0_321 
* INOUT : bl_0_322 
* INOUT : br_0_322 
* INOUT : bl_0_323 
* INOUT : br_0_323 
* INOUT : bl_0_324 
* INOUT : br_0_324 
* INOUT : bl_0_325 
* INOUT : br_0_325 
* INOUT : bl_0_326 
* INOUT : br_0_326 
* INOUT : bl_0_327 
* INOUT : br_0_327 
* INOUT : bl_0_328 
* INOUT : br_0_328 
* INOUT : bl_0_329 
* INOUT : br_0_329 
* INOUT : bl_0_330 
* INOUT : br_0_330 
* INOUT : bl_0_331 
* INOUT : br_0_331 
* INOUT : bl_0_332 
* INOUT : br_0_332 
* INOUT : bl_0_333 
* INOUT : br_0_333 
* INOUT : bl_0_334 
* INOUT : br_0_334 
* INOUT : bl_0_335 
* INOUT : br_0_335 
* INOUT : bl_0_336 
* INOUT : br_0_336 
* INOUT : bl_0_337 
* INOUT : br_0_337 
* INOUT : bl_0_338 
* INOUT : br_0_338 
* INOUT : bl_0_339 
* INOUT : br_0_339 
* INOUT : bl_0_340 
* INOUT : br_0_340 
* INOUT : bl_0_341 
* INOUT : br_0_341 
* INOUT : bl_0_342 
* INOUT : br_0_342 
* INOUT : bl_0_343 
* INOUT : br_0_343 
* INOUT : bl_0_344 
* INOUT : br_0_344 
* INOUT : bl_0_345 
* INOUT : br_0_345 
* INOUT : bl_0_346 
* INOUT : br_0_346 
* INOUT : bl_0_347 
* INOUT : br_0_347 
* INOUT : bl_0_348 
* INOUT : br_0_348 
* INOUT : bl_0_349 
* INOUT : br_0_349 
* INOUT : bl_0_350 
* INOUT : br_0_350 
* INOUT : bl_0_351 
* INOUT : br_0_351 
* INOUT : bl_0_352 
* INOUT : br_0_352 
* INOUT : bl_0_353 
* INOUT : br_0_353 
* INOUT : bl_0_354 
* INOUT : br_0_354 
* INOUT : bl_0_355 
* INOUT : br_0_355 
* INOUT : bl_0_356 
* INOUT : br_0_356 
* INOUT : bl_0_357 
* INOUT : br_0_357 
* INOUT : bl_0_358 
* INOUT : br_0_358 
* INOUT : bl_0_359 
* INOUT : br_0_359 
* INOUT : bl_0_360 
* INOUT : br_0_360 
* INOUT : bl_0_361 
* INOUT : br_0_361 
* INOUT : bl_0_362 
* INOUT : br_0_362 
* INOUT : bl_0_363 
* INOUT : br_0_363 
* INOUT : bl_0_364 
* INOUT : br_0_364 
* INOUT : bl_0_365 
* INOUT : br_0_365 
* INOUT : bl_0_366 
* INOUT : br_0_366 
* INOUT : bl_0_367 
* INOUT : br_0_367 
* INOUT : bl_0_368 
* INOUT : br_0_368 
* INOUT : bl_0_369 
* INOUT : br_0_369 
* INOUT : bl_0_370 
* INOUT : br_0_370 
* INOUT : bl_0_371 
* INOUT : br_0_371 
* INOUT : bl_0_372 
* INOUT : br_0_372 
* INOUT : bl_0_373 
* INOUT : br_0_373 
* INOUT : bl_0_374 
* INOUT : br_0_374 
* INOUT : bl_0_375 
* INOUT : br_0_375 
* INOUT : bl_0_376 
* INOUT : br_0_376 
* INOUT : bl_0_377 
* INOUT : br_0_377 
* INOUT : bl_0_378 
* INOUT : br_0_378 
* INOUT : bl_0_379 
* INOUT : br_0_379 
* INOUT : bl_0_380 
* INOUT : br_0_380 
* INOUT : bl_0_381 
* INOUT : br_0_381 
* INOUT : bl_0_382 
* INOUT : br_0_382 
* INOUT : bl_0_383 
* INOUT : br_0_383 
* INOUT : bl_0_384 
* INOUT : br_0_384 
* INOUT : bl_0_385 
* INOUT : br_0_385 
* INOUT : bl_0_386 
* INOUT : br_0_386 
* INOUT : bl_0_387 
* INOUT : br_0_387 
* INOUT : bl_0_388 
* INOUT : br_0_388 
* INOUT : bl_0_389 
* INOUT : br_0_389 
* INOUT : bl_0_390 
* INOUT : br_0_390 
* INOUT : bl_0_391 
* INOUT : br_0_391 
* INOUT : bl_0_392 
* INOUT : br_0_392 
* INOUT : bl_0_393 
* INOUT : br_0_393 
* INOUT : bl_0_394 
* INOUT : br_0_394 
* INOUT : bl_0_395 
* INOUT : br_0_395 
* INOUT : bl_0_396 
* INOUT : br_0_396 
* INOUT : bl_0_397 
* INOUT : br_0_397 
* INOUT : bl_0_398 
* INOUT : br_0_398 
* INOUT : bl_0_399 
* INOUT : br_0_399 
* INOUT : bl_0_400 
* INOUT : br_0_400 
* INOUT : bl_0_401 
* INOUT : br_0_401 
* INOUT : bl_0_402 
* INOUT : br_0_402 
* INOUT : bl_0_403 
* INOUT : br_0_403 
* INOUT : bl_0_404 
* INOUT : br_0_404 
* INOUT : bl_0_405 
* INOUT : br_0_405 
* INOUT : bl_0_406 
* INOUT : br_0_406 
* INOUT : bl_0_407 
* INOUT : br_0_407 
* INOUT : bl_0_408 
* INOUT : br_0_408 
* INOUT : bl_0_409 
* INOUT : br_0_409 
* INOUT : bl_0_410 
* INOUT : br_0_410 
* INOUT : bl_0_411 
* INOUT : br_0_411 
* INOUT : bl_0_412 
* INOUT : br_0_412 
* INOUT : bl_0_413 
* INOUT : br_0_413 
* INOUT : bl_0_414 
* INOUT : br_0_414 
* INOUT : bl_0_415 
* INOUT : br_0_415 
* INOUT : bl_0_416 
* INOUT : br_0_416 
* INOUT : bl_0_417 
* INOUT : br_0_417 
* INOUT : bl_0_418 
* INOUT : br_0_418 
* INOUT : bl_0_419 
* INOUT : br_0_419 
* INOUT : bl_0_420 
* INOUT : br_0_420 
* INOUT : bl_0_421 
* INOUT : br_0_421 
* INOUT : bl_0_422 
* INOUT : br_0_422 
* INOUT : bl_0_423 
* INOUT : br_0_423 
* INOUT : bl_0_424 
* INOUT : br_0_424 
* INOUT : bl_0_425 
* INOUT : br_0_425 
* INOUT : bl_0_426 
* INOUT : br_0_426 
* INOUT : bl_0_427 
* INOUT : br_0_427 
* INOUT : bl_0_428 
* INOUT : br_0_428 
* INOUT : bl_0_429 
* INOUT : br_0_429 
* INOUT : bl_0_430 
* INOUT : br_0_430 
* INOUT : bl_0_431 
* INOUT : br_0_431 
* INOUT : bl_0_432 
* INOUT : br_0_432 
* INOUT : bl_0_433 
* INOUT : br_0_433 
* INOUT : bl_0_434 
* INOUT : br_0_434 
* INOUT : bl_0_435 
* INOUT : br_0_435 
* INOUT : bl_0_436 
* INOUT : br_0_436 
* INOUT : bl_0_437 
* INOUT : br_0_437 
* INOUT : bl_0_438 
* INOUT : br_0_438 
* INOUT : bl_0_439 
* INOUT : br_0_439 
* INOUT : bl_0_440 
* INOUT : br_0_440 
* INOUT : bl_0_441 
* INOUT : br_0_441 
* INOUT : bl_0_442 
* INOUT : br_0_442 
* INOUT : bl_0_443 
* INOUT : br_0_443 
* INOUT : bl_0_444 
* INOUT : br_0_444 
* INOUT : bl_0_445 
* INOUT : br_0_445 
* INOUT : bl_0_446 
* INOUT : br_0_446 
* INOUT : bl_0_447 
* INOUT : br_0_447 
* INOUT : bl_0_448 
* INOUT : br_0_448 
* INOUT : bl_0_449 
* INOUT : br_0_449 
* INOUT : bl_0_450 
* INOUT : br_0_450 
* INOUT : bl_0_451 
* INOUT : br_0_451 
* INOUT : bl_0_452 
* INOUT : br_0_452 
* INOUT : bl_0_453 
* INOUT : br_0_453 
* INOUT : bl_0_454 
* INOUT : br_0_454 
* INOUT : bl_0_455 
* INOUT : br_0_455 
* INOUT : bl_0_456 
* INOUT : br_0_456 
* INOUT : bl_0_457 
* INOUT : br_0_457 
* INOUT : bl_0_458 
* INOUT : br_0_458 
* INOUT : bl_0_459 
* INOUT : br_0_459 
* INOUT : bl_0_460 
* INOUT : br_0_460 
* INOUT : bl_0_461 
* INOUT : br_0_461 
* INOUT : bl_0_462 
* INOUT : br_0_462 
* INOUT : bl_0_463 
* INOUT : br_0_463 
* INOUT : bl_0_464 
* INOUT : br_0_464 
* INOUT : bl_0_465 
* INOUT : br_0_465 
* INOUT : bl_0_466 
* INOUT : br_0_466 
* INOUT : bl_0_467 
* INOUT : br_0_467 
* INOUT : bl_0_468 
* INOUT : br_0_468 
* INOUT : bl_0_469 
* INOUT : br_0_469 
* INOUT : bl_0_470 
* INOUT : br_0_470 
* INOUT : bl_0_471 
* INOUT : br_0_471 
* INOUT : bl_0_472 
* INOUT : br_0_472 
* INOUT : bl_0_473 
* INOUT : br_0_473 
* INOUT : bl_0_474 
* INOUT : br_0_474 
* INOUT : bl_0_475 
* INOUT : br_0_475 
* INOUT : bl_0_476 
* INOUT : br_0_476 
* INOUT : bl_0_477 
* INOUT : br_0_477 
* INOUT : bl_0_478 
* INOUT : br_0_478 
* INOUT : bl_0_479 
* INOUT : br_0_479 
* INOUT : bl_0_480 
* INOUT : br_0_480 
* INOUT : bl_0_481 
* INOUT : br_0_481 
* INOUT : bl_0_482 
* INOUT : br_0_482 
* INOUT : bl_0_483 
* INOUT : br_0_483 
* INOUT : bl_0_484 
* INOUT : br_0_484 
* INOUT : bl_0_485 
* INOUT : br_0_485 
* INOUT : bl_0_486 
* INOUT : br_0_486 
* INOUT : bl_0_487 
* INOUT : br_0_487 
* INOUT : bl_0_488 
* INOUT : br_0_488 
* INOUT : bl_0_489 
* INOUT : br_0_489 
* INOUT : bl_0_490 
* INOUT : br_0_490 
* INOUT : bl_0_491 
* INOUT : br_0_491 
* INOUT : bl_0_492 
* INOUT : br_0_492 
* INOUT : bl_0_493 
* INOUT : br_0_493 
* INOUT : bl_0_494 
* INOUT : br_0_494 
* INOUT : bl_0_495 
* INOUT : br_0_495 
* INOUT : bl_0_496 
* INOUT : br_0_496 
* INOUT : bl_0_497 
* INOUT : br_0_497 
* INOUT : bl_0_498 
* INOUT : br_0_498 
* INOUT : bl_0_499 
* INOUT : br_0_499 
* INOUT : bl_0_500 
* INOUT : br_0_500 
* INOUT : bl_0_501 
* INOUT : br_0_501 
* INOUT : bl_0_502 
* INOUT : br_0_502 
* INOUT : bl_0_503 
* INOUT : br_0_503 
* INOUT : bl_0_504 
* INOUT : br_0_504 
* INOUT : bl_0_505 
* INOUT : br_0_505 
* INOUT : bl_0_506 
* INOUT : br_0_506 
* INOUT : bl_0_507 
* INOUT : br_0_507 
* INOUT : bl_0_508 
* INOUT : br_0_508 
* INOUT : bl_0_509 
* INOUT : br_0_509 
* INOUT : bl_0_510 
* INOUT : br_0_510 
* INOUT : bl_0_511 
* INOUT : br_0_511 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* POWER : vdd 
* GROUND: gnd 
* rows: 45 cols: 512
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c0
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c0
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c0
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c0
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c0
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c0
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c0
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c0
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c0
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c0
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c1
+ bl_0_1 br_0_1 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c1
+ bl_0_1 br_0_1 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c1
+ bl_0_1 br_0_1 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c1
+ bl_0_1 br_0_1 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c1
+ bl_0_1 br_0_1 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c1
+ bl_0_1 br_0_1 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c1
+ bl_0_1 br_0_1 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c1
+ bl_0_1 br_0_1 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c1
+ bl_0_1 br_0_1 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c1
+ bl_0_1 br_0_1 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c1
+ bl_0_1 br_0_1 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c1
+ bl_0_1 br_0_1 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c1
+ bl_0_1 br_0_1 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c1
+ bl_0_1 br_0_1 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c1
+ bl_0_1 br_0_1 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c1
+ bl_0_1 br_0_1 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c1
+ bl_0_1 br_0_1 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c1
+ bl_0_1 br_0_1 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c1
+ bl_0_1 br_0_1 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c1
+ bl_0_1 br_0_1 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c1
+ bl_0_1 br_0_1 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c1
+ bl_0_1 br_0_1 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c1
+ bl_0_1 br_0_1 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c1
+ bl_0_1 br_0_1 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c1
+ bl_0_1 br_0_1 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c1
+ bl_0_1 br_0_1 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c1
+ bl_0_1 br_0_1 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c1
+ bl_0_1 br_0_1 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c1
+ bl_0_1 br_0_1 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c1
+ bl_0_1 br_0_1 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c1
+ bl_0_1 br_0_1 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c1
+ bl_0_1 br_0_1 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c1
+ bl_0_1 br_0_1 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c1
+ bl_0_1 br_0_1 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c1
+ bl_0_1 br_0_1 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c1
+ bl_0_1 br_0_1 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c1
+ bl_0_1 br_0_1 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c1
+ bl_0_1 br_0_1 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c1
+ bl_0_1 br_0_1 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c1
+ bl_0_1 br_0_1 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c1
+ bl_0_1 br_0_1 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c1
+ bl_0_1 br_0_1 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c1
+ bl_0_1 br_0_1 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c1
+ bl_0_1 br_0_1 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c2
+ bl_0_2 br_0_2 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c2
+ bl_0_2 br_0_2 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c2
+ bl_0_2 br_0_2 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c2
+ bl_0_2 br_0_2 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c2
+ bl_0_2 br_0_2 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c2
+ bl_0_2 br_0_2 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c2
+ bl_0_2 br_0_2 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c2
+ bl_0_2 br_0_2 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c2
+ bl_0_2 br_0_2 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c2
+ bl_0_2 br_0_2 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c2
+ bl_0_2 br_0_2 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c2
+ bl_0_2 br_0_2 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c2
+ bl_0_2 br_0_2 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c2
+ bl_0_2 br_0_2 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c2
+ bl_0_2 br_0_2 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c2
+ bl_0_2 br_0_2 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c2
+ bl_0_2 br_0_2 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c2
+ bl_0_2 br_0_2 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c2
+ bl_0_2 br_0_2 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c2
+ bl_0_2 br_0_2 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c2
+ bl_0_2 br_0_2 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c2
+ bl_0_2 br_0_2 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c2
+ bl_0_2 br_0_2 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c2
+ bl_0_2 br_0_2 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c2
+ bl_0_2 br_0_2 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c2
+ bl_0_2 br_0_2 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c2
+ bl_0_2 br_0_2 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c2
+ bl_0_2 br_0_2 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c2
+ bl_0_2 br_0_2 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c2
+ bl_0_2 br_0_2 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c2
+ bl_0_2 br_0_2 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c2
+ bl_0_2 br_0_2 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c2
+ bl_0_2 br_0_2 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c2
+ bl_0_2 br_0_2 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c2
+ bl_0_2 br_0_2 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c2
+ bl_0_2 br_0_2 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c2
+ bl_0_2 br_0_2 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c2
+ bl_0_2 br_0_2 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c2
+ bl_0_2 br_0_2 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c2
+ bl_0_2 br_0_2 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c2
+ bl_0_2 br_0_2 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c2
+ bl_0_2 br_0_2 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c2
+ bl_0_2 br_0_2 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c2
+ bl_0_2 br_0_2 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c3
+ bl_0_3 br_0_3 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c3
+ bl_0_3 br_0_3 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c3
+ bl_0_3 br_0_3 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c3
+ bl_0_3 br_0_3 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c3
+ bl_0_3 br_0_3 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c3
+ bl_0_3 br_0_3 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c3
+ bl_0_3 br_0_3 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c3
+ bl_0_3 br_0_3 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c3
+ bl_0_3 br_0_3 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c3
+ bl_0_3 br_0_3 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c3
+ bl_0_3 br_0_3 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c3
+ bl_0_3 br_0_3 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c3
+ bl_0_3 br_0_3 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c3
+ bl_0_3 br_0_3 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c3
+ bl_0_3 br_0_3 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c3
+ bl_0_3 br_0_3 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c3
+ bl_0_3 br_0_3 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c3
+ bl_0_3 br_0_3 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c3
+ bl_0_3 br_0_3 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c3
+ bl_0_3 br_0_3 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c3
+ bl_0_3 br_0_3 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c3
+ bl_0_3 br_0_3 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c3
+ bl_0_3 br_0_3 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c3
+ bl_0_3 br_0_3 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c3
+ bl_0_3 br_0_3 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c3
+ bl_0_3 br_0_3 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c3
+ bl_0_3 br_0_3 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c3
+ bl_0_3 br_0_3 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c3
+ bl_0_3 br_0_3 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c3
+ bl_0_3 br_0_3 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c3
+ bl_0_3 br_0_3 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c3
+ bl_0_3 br_0_3 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c3
+ bl_0_3 br_0_3 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c3
+ bl_0_3 br_0_3 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c3
+ bl_0_3 br_0_3 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c3
+ bl_0_3 br_0_3 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c3
+ bl_0_3 br_0_3 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c3
+ bl_0_3 br_0_3 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c3
+ bl_0_3 br_0_3 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c3
+ bl_0_3 br_0_3 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c3
+ bl_0_3 br_0_3 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c3
+ bl_0_3 br_0_3 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c3
+ bl_0_3 br_0_3 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c3
+ bl_0_3 br_0_3 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c4
+ bl_0_4 br_0_4 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c4
+ bl_0_4 br_0_4 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c4
+ bl_0_4 br_0_4 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c4
+ bl_0_4 br_0_4 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c4
+ bl_0_4 br_0_4 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c4
+ bl_0_4 br_0_4 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c4
+ bl_0_4 br_0_4 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c4
+ bl_0_4 br_0_4 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c4
+ bl_0_4 br_0_4 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c4
+ bl_0_4 br_0_4 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c4
+ bl_0_4 br_0_4 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c4
+ bl_0_4 br_0_4 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c4
+ bl_0_4 br_0_4 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c4
+ bl_0_4 br_0_4 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c4
+ bl_0_4 br_0_4 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c4
+ bl_0_4 br_0_4 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c4
+ bl_0_4 br_0_4 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c4
+ bl_0_4 br_0_4 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c4
+ bl_0_4 br_0_4 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c4
+ bl_0_4 br_0_4 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c4
+ bl_0_4 br_0_4 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c4
+ bl_0_4 br_0_4 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c4
+ bl_0_4 br_0_4 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c4
+ bl_0_4 br_0_4 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c4
+ bl_0_4 br_0_4 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c4
+ bl_0_4 br_0_4 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c4
+ bl_0_4 br_0_4 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c4
+ bl_0_4 br_0_4 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c4
+ bl_0_4 br_0_4 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c4
+ bl_0_4 br_0_4 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c4
+ bl_0_4 br_0_4 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c4
+ bl_0_4 br_0_4 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c4
+ bl_0_4 br_0_4 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c4
+ bl_0_4 br_0_4 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c4
+ bl_0_4 br_0_4 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c4
+ bl_0_4 br_0_4 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c4
+ bl_0_4 br_0_4 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c4
+ bl_0_4 br_0_4 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c4
+ bl_0_4 br_0_4 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c4
+ bl_0_4 br_0_4 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c4
+ bl_0_4 br_0_4 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c4
+ bl_0_4 br_0_4 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c4
+ bl_0_4 br_0_4 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c4
+ bl_0_4 br_0_4 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c5
+ bl_0_5 br_0_5 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c5
+ bl_0_5 br_0_5 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c5
+ bl_0_5 br_0_5 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c5
+ bl_0_5 br_0_5 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c5
+ bl_0_5 br_0_5 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c5
+ bl_0_5 br_0_5 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c5
+ bl_0_5 br_0_5 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c5
+ bl_0_5 br_0_5 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c5
+ bl_0_5 br_0_5 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c5
+ bl_0_5 br_0_5 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c5
+ bl_0_5 br_0_5 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c5
+ bl_0_5 br_0_5 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c5
+ bl_0_5 br_0_5 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c5
+ bl_0_5 br_0_5 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c5
+ bl_0_5 br_0_5 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c5
+ bl_0_5 br_0_5 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c5
+ bl_0_5 br_0_5 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c5
+ bl_0_5 br_0_5 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c5
+ bl_0_5 br_0_5 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c5
+ bl_0_5 br_0_5 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c5
+ bl_0_5 br_0_5 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c5
+ bl_0_5 br_0_5 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c5
+ bl_0_5 br_0_5 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c5
+ bl_0_5 br_0_5 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c5
+ bl_0_5 br_0_5 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c5
+ bl_0_5 br_0_5 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c5
+ bl_0_5 br_0_5 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c5
+ bl_0_5 br_0_5 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c5
+ bl_0_5 br_0_5 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c5
+ bl_0_5 br_0_5 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c5
+ bl_0_5 br_0_5 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c5
+ bl_0_5 br_0_5 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c5
+ bl_0_5 br_0_5 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c5
+ bl_0_5 br_0_5 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c5
+ bl_0_5 br_0_5 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c5
+ bl_0_5 br_0_5 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c5
+ bl_0_5 br_0_5 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c5
+ bl_0_5 br_0_5 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c5
+ bl_0_5 br_0_5 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c5
+ bl_0_5 br_0_5 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c5
+ bl_0_5 br_0_5 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c5
+ bl_0_5 br_0_5 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c5
+ bl_0_5 br_0_5 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c5
+ bl_0_5 br_0_5 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c6
+ bl_0_6 br_0_6 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c6
+ bl_0_6 br_0_6 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c6
+ bl_0_6 br_0_6 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c6
+ bl_0_6 br_0_6 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c6
+ bl_0_6 br_0_6 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c6
+ bl_0_6 br_0_6 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c6
+ bl_0_6 br_0_6 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c6
+ bl_0_6 br_0_6 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c6
+ bl_0_6 br_0_6 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c6
+ bl_0_6 br_0_6 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c6
+ bl_0_6 br_0_6 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c6
+ bl_0_6 br_0_6 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c6
+ bl_0_6 br_0_6 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c6
+ bl_0_6 br_0_6 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c6
+ bl_0_6 br_0_6 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c6
+ bl_0_6 br_0_6 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c6
+ bl_0_6 br_0_6 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c6
+ bl_0_6 br_0_6 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c6
+ bl_0_6 br_0_6 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c6
+ bl_0_6 br_0_6 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c6
+ bl_0_6 br_0_6 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c6
+ bl_0_6 br_0_6 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c6
+ bl_0_6 br_0_6 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c6
+ bl_0_6 br_0_6 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c6
+ bl_0_6 br_0_6 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c6
+ bl_0_6 br_0_6 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c6
+ bl_0_6 br_0_6 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c6
+ bl_0_6 br_0_6 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c6
+ bl_0_6 br_0_6 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c6
+ bl_0_6 br_0_6 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c6
+ bl_0_6 br_0_6 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c6
+ bl_0_6 br_0_6 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c6
+ bl_0_6 br_0_6 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c6
+ bl_0_6 br_0_6 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c6
+ bl_0_6 br_0_6 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c6
+ bl_0_6 br_0_6 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c6
+ bl_0_6 br_0_6 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c6
+ bl_0_6 br_0_6 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c6
+ bl_0_6 br_0_6 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c6
+ bl_0_6 br_0_6 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c6
+ bl_0_6 br_0_6 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c6
+ bl_0_6 br_0_6 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c6
+ bl_0_6 br_0_6 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c6
+ bl_0_6 br_0_6 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c7
+ bl_0_7 br_0_7 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c7
+ bl_0_7 br_0_7 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c7
+ bl_0_7 br_0_7 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c7
+ bl_0_7 br_0_7 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c7
+ bl_0_7 br_0_7 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c7
+ bl_0_7 br_0_7 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c7
+ bl_0_7 br_0_7 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c7
+ bl_0_7 br_0_7 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c7
+ bl_0_7 br_0_7 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c7
+ bl_0_7 br_0_7 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c7
+ bl_0_7 br_0_7 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c7
+ bl_0_7 br_0_7 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c7
+ bl_0_7 br_0_7 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c7
+ bl_0_7 br_0_7 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c7
+ bl_0_7 br_0_7 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c7
+ bl_0_7 br_0_7 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c7
+ bl_0_7 br_0_7 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c7
+ bl_0_7 br_0_7 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c7
+ bl_0_7 br_0_7 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c7
+ bl_0_7 br_0_7 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c7
+ bl_0_7 br_0_7 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c7
+ bl_0_7 br_0_7 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c7
+ bl_0_7 br_0_7 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c7
+ bl_0_7 br_0_7 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c7
+ bl_0_7 br_0_7 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c7
+ bl_0_7 br_0_7 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c7
+ bl_0_7 br_0_7 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c7
+ bl_0_7 br_0_7 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c7
+ bl_0_7 br_0_7 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c7
+ bl_0_7 br_0_7 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c7
+ bl_0_7 br_0_7 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c7
+ bl_0_7 br_0_7 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c7
+ bl_0_7 br_0_7 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c7
+ bl_0_7 br_0_7 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c7
+ bl_0_7 br_0_7 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c7
+ bl_0_7 br_0_7 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c7
+ bl_0_7 br_0_7 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c7
+ bl_0_7 br_0_7 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c7
+ bl_0_7 br_0_7 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c7
+ bl_0_7 br_0_7 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c7
+ bl_0_7 br_0_7 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c7
+ bl_0_7 br_0_7 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c7
+ bl_0_7 br_0_7 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c7
+ bl_0_7 br_0_7 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c8
+ bl_0_8 br_0_8 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c8
+ bl_0_8 br_0_8 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c8
+ bl_0_8 br_0_8 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c8
+ bl_0_8 br_0_8 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c8
+ bl_0_8 br_0_8 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c8
+ bl_0_8 br_0_8 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c8
+ bl_0_8 br_0_8 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c8
+ bl_0_8 br_0_8 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c8
+ bl_0_8 br_0_8 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c8
+ bl_0_8 br_0_8 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c8
+ bl_0_8 br_0_8 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c8
+ bl_0_8 br_0_8 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c8
+ bl_0_8 br_0_8 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c8
+ bl_0_8 br_0_8 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c8
+ bl_0_8 br_0_8 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c8
+ bl_0_8 br_0_8 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c8
+ bl_0_8 br_0_8 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c8
+ bl_0_8 br_0_8 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c8
+ bl_0_8 br_0_8 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c8
+ bl_0_8 br_0_8 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c8
+ bl_0_8 br_0_8 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c8
+ bl_0_8 br_0_8 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c8
+ bl_0_8 br_0_8 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c8
+ bl_0_8 br_0_8 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c8
+ bl_0_8 br_0_8 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c8
+ bl_0_8 br_0_8 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c8
+ bl_0_8 br_0_8 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c8
+ bl_0_8 br_0_8 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c8
+ bl_0_8 br_0_8 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c8
+ bl_0_8 br_0_8 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c8
+ bl_0_8 br_0_8 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c8
+ bl_0_8 br_0_8 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c8
+ bl_0_8 br_0_8 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c8
+ bl_0_8 br_0_8 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c8
+ bl_0_8 br_0_8 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c8
+ bl_0_8 br_0_8 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c8
+ bl_0_8 br_0_8 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c8
+ bl_0_8 br_0_8 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c8
+ bl_0_8 br_0_8 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c8
+ bl_0_8 br_0_8 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c8
+ bl_0_8 br_0_8 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c8
+ bl_0_8 br_0_8 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c8
+ bl_0_8 br_0_8 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c8
+ bl_0_8 br_0_8 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c9
+ bl_0_9 br_0_9 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c9
+ bl_0_9 br_0_9 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c9
+ bl_0_9 br_0_9 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c9
+ bl_0_9 br_0_9 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c9
+ bl_0_9 br_0_9 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c9
+ bl_0_9 br_0_9 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c9
+ bl_0_9 br_0_9 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c9
+ bl_0_9 br_0_9 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c9
+ bl_0_9 br_0_9 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c9
+ bl_0_9 br_0_9 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c9
+ bl_0_9 br_0_9 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c9
+ bl_0_9 br_0_9 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c9
+ bl_0_9 br_0_9 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c9
+ bl_0_9 br_0_9 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c9
+ bl_0_9 br_0_9 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c9
+ bl_0_9 br_0_9 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c9
+ bl_0_9 br_0_9 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c9
+ bl_0_9 br_0_9 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c9
+ bl_0_9 br_0_9 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c9
+ bl_0_9 br_0_9 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c9
+ bl_0_9 br_0_9 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c9
+ bl_0_9 br_0_9 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c9
+ bl_0_9 br_0_9 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c9
+ bl_0_9 br_0_9 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c9
+ bl_0_9 br_0_9 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c9
+ bl_0_9 br_0_9 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c9
+ bl_0_9 br_0_9 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c9
+ bl_0_9 br_0_9 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c9
+ bl_0_9 br_0_9 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c9
+ bl_0_9 br_0_9 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c9
+ bl_0_9 br_0_9 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c9
+ bl_0_9 br_0_9 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c9
+ bl_0_9 br_0_9 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c9
+ bl_0_9 br_0_9 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c9
+ bl_0_9 br_0_9 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c9
+ bl_0_9 br_0_9 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c9
+ bl_0_9 br_0_9 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c9
+ bl_0_9 br_0_9 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c9
+ bl_0_9 br_0_9 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c9
+ bl_0_9 br_0_9 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c9
+ bl_0_9 br_0_9 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c9
+ bl_0_9 br_0_9 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c9
+ bl_0_9 br_0_9 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c9
+ bl_0_9 br_0_9 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c10
+ bl_0_10 br_0_10 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c10
+ bl_0_10 br_0_10 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c10
+ bl_0_10 br_0_10 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c10
+ bl_0_10 br_0_10 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c10
+ bl_0_10 br_0_10 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c10
+ bl_0_10 br_0_10 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c10
+ bl_0_10 br_0_10 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c10
+ bl_0_10 br_0_10 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c10
+ bl_0_10 br_0_10 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c10
+ bl_0_10 br_0_10 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c10
+ bl_0_10 br_0_10 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c10
+ bl_0_10 br_0_10 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c10
+ bl_0_10 br_0_10 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c10
+ bl_0_10 br_0_10 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c10
+ bl_0_10 br_0_10 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c10
+ bl_0_10 br_0_10 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c10
+ bl_0_10 br_0_10 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c10
+ bl_0_10 br_0_10 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c10
+ bl_0_10 br_0_10 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c10
+ bl_0_10 br_0_10 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c10
+ bl_0_10 br_0_10 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c10
+ bl_0_10 br_0_10 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c10
+ bl_0_10 br_0_10 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c10
+ bl_0_10 br_0_10 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c10
+ bl_0_10 br_0_10 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c10
+ bl_0_10 br_0_10 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c10
+ bl_0_10 br_0_10 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c10
+ bl_0_10 br_0_10 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c10
+ bl_0_10 br_0_10 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c10
+ bl_0_10 br_0_10 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c10
+ bl_0_10 br_0_10 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c10
+ bl_0_10 br_0_10 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c10
+ bl_0_10 br_0_10 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c10
+ bl_0_10 br_0_10 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c10
+ bl_0_10 br_0_10 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c10
+ bl_0_10 br_0_10 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c10
+ bl_0_10 br_0_10 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c10
+ bl_0_10 br_0_10 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c10
+ bl_0_10 br_0_10 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c10
+ bl_0_10 br_0_10 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c10
+ bl_0_10 br_0_10 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c10
+ bl_0_10 br_0_10 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c10
+ bl_0_10 br_0_10 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c10
+ bl_0_10 br_0_10 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c11
+ bl_0_11 br_0_11 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c11
+ bl_0_11 br_0_11 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c11
+ bl_0_11 br_0_11 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c11
+ bl_0_11 br_0_11 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c11
+ bl_0_11 br_0_11 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c11
+ bl_0_11 br_0_11 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c11
+ bl_0_11 br_0_11 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c11
+ bl_0_11 br_0_11 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c11
+ bl_0_11 br_0_11 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c11
+ bl_0_11 br_0_11 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c11
+ bl_0_11 br_0_11 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c11
+ bl_0_11 br_0_11 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c11
+ bl_0_11 br_0_11 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c11
+ bl_0_11 br_0_11 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c11
+ bl_0_11 br_0_11 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c11
+ bl_0_11 br_0_11 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c11
+ bl_0_11 br_0_11 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c11
+ bl_0_11 br_0_11 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c11
+ bl_0_11 br_0_11 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c11
+ bl_0_11 br_0_11 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c11
+ bl_0_11 br_0_11 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c11
+ bl_0_11 br_0_11 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c11
+ bl_0_11 br_0_11 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c11
+ bl_0_11 br_0_11 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c11
+ bl_0_11 br_0_11 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c11
+ bl_0_11 br_0_11 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c11
+ bl_0_11 br_0_11 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c11
+ bl_0_11 br_0_11 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c11
+ bl_0_11 br_0_11 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c11
+ bl_0_11 br_0_11 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c11
+ bl_0_11 br_0_11 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c11
+ bl_0_11 br_0_11 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c11
+ bl_0_11 br_0_11 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c11
+ bl_0_11 br_0_11 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c11
+ bl_0_11 br_0_11 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c11
+ bl_0_11 br_0_11 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c11
+ bl_0_11 br_0_11 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c11
+ bl_0_11 br_0_11 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c11
+ bl_0_11 br_0_11 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c11
+ bl_0_11 br_0_11 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c11
+ bl_0_11 br_0_11 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c11
+ bl_0_11 br_0_11 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c11
+ bl_0_11 br_0_11 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c11
+ bl_0_11 br_0_11 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c12
+ bl_0_12 br_0_12 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c12
+ bl_0_12 br_0_12 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c12
+ bl_0_12 br_0_12 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c12
+ bl_0_12 br_0_12 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c12
+ bl_0_12 br_0_12 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c12
+ bl_0_12 br_0_12 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c12
+ bl_0_12 br_0_12 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c12
+ bl_0_12 br_0_12 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c12
+ bl_0_12 br_0_12 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c12
+ bl_0_12 br_0_12 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c12
+ bl_0_12 br_0_12 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c12
+ bl_0_12 br_0_12 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c12
+ bl_0_12 br_0_12 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c12
+ bl_0_12 br_0_12 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c12
+ bl_0_12 br_0_12 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c12
+ bl_0_12 br_0_12 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c12
+ bl_0_12 br_0_12 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c12
+ bl_0_12 br_0_12 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c12
+ bl_0_12 br_0_12 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c12
+ bl_0_12 br_0_12 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c12
+ bl_0_12 br_0_12 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c12
+ bl_0_12 br_0_12 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c12
+ bl_0_12 br_0_12 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c12
+ bl_0_12 br_0_12 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c12
+ bl_0_12 br_0_12 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c12
+ bl_0_12 br_0_12 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c12
+ bl_0_12 br_0_12 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c12
+ bl_0_12 br_0_12 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c12
+ bl_0_12 br_0_12 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c12
+ bl_0_12 br_0_12 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c12
+ bl_0_12 br_0_12 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c12
+ bl_0_12 br_0_12 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c12
+ bl_0_12 br_0_12 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c12
+ bl_0_12 br_0_12 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c12
+ bl_0_12 br_0_12 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c12
+ bl_0_12 br_0_12 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c12
+ bl_0_12 br_0_12 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c12
+ bl_0_12 br_0_12 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c12
+ bl_0_12 br_0_12 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c12
+ bl_0_12 br_0_12 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c12
+ bl_0_12 br_0_12 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c12
+ bl_0_12 br_0_12 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c12
+ bl_0_12 br_0_12 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c12
+ bl_0_12 br_0_12 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c13
+ bl_0_13 br_0_13 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c13
+ bl_0_13 br_0_13 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c13
+ bl_0_13 br_0_13 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c13
+ bl_0_13 br_0_13 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c13
+ bl_0_13 br_0_13 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c13
+ bl_0_13 br_0_13 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c13
+ bl_0_13 br_0_13 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c13
+ bl_0_13 br_0_13 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c13
+ bl_0_13 br_0_13 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c13
+ bl_0_13 br_0_13 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c13
+ bl_0_13 br_0_13 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c13
+ bl_0_13 br_0_13 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c13
+ bl_0_13 br_0_13 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c13
+ bl_0_13 br_0_13 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c13
+ bl_0_13 br_0_13 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c13
+ bl_0_13 br_0_13 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c13
+ bl_0_13 br_0_13 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c13
+ bl_0_13 br_0_13 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c13
+ bl_0_13 br_0_13 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c13
+ bl_0_13 br_0_13 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c13
+ bl_0_13 br_0_13 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c13
+ bl_0_13 br_0_13 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c13
+ bl_0_13 br_0_13 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c13
+ bl_0_13 br_0_13 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c13
+ bl_0_13 br_0_13 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c13
+ bl_0_13 br_0_13 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c13
+ bl_0_13 br_0_13 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c13
+ bl_0_13 br_0_13 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c13
+ bl_0_13 br_0_13 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c13
+ bl_0_13 br_0_13 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c13
+ bl_0_13 br_0_13 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c13
+ bl_0_13 br_0_13 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c13
+ bl_0_13 br_0_13 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c13
+ bl_0_13 br_0_13 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c13
+ bl_0_13 br_0_13 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c13
+ bl_0_13 br_0_13 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c13
+ bl_0_13 br_0_13 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c13
+ bl_0_13 br_0_13 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c13
+ bl_0_13 br_0_13 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c13
+ bl_0_13 br_0_13 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c13
+ bl_0_13 br_0_13 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c13
+ bl_0_13 br_0_13 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c13
+ bl_0_13 br_0_13 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c13
+ bl_0_13 br_0_13 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c14
+ bl_0_14 br_0_14 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c14
+ bl_0_14 br_0_14 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c14
+ bl_0_14 br_0_14 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c14
+ bl_0_14 br_0_14 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c14
+ bl_0_14 br_0_14 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c14
+ bl_0_14 br_0_14 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c14
+ bl_0_14 br_0_14 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c14
+ bl_0_14 br_0_14 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c14
+ bl_0_14 br_0_14 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c14
+ bl_0_14 br_0_14 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c14
+ bl_0_14 br_0_14 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c14
+ bl_0_14 br_0_14 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c14
+ bl_0_14 br_0_14 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c14
+ bl_0_14 br_0_14 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c14
+ bl_0_14 br_0_14 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c14
+ bl_0_14 br_0_14 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c14
+ bl_0_14 br_0_14 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c14
+ bl_0_14 br_0_14 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c14
+ bl_0_14 br_0_14 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c14
+ bl_0_14 br_0_14 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c14
+ bl_0_14 br_0_14 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c14
+ bl_0_14 br_0_14 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c14
+ bl_0_14 br_0_14 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c14
+ bl_0_14 br_0_14 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c14
+ bl_0_14 br_0_14 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c14
+ bl_0_14 br_0_14 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c14
+ bl_0_14 br_0_14 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c14
+ bl_0_14 br_0_14 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c14
+ bl_0_14 br_0_14 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c14
+ bl_0_14 br_0_14 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c14
+ bl_0_14 br_0_14 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c14
+ bl_0_14 br_0_14 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c14
+ bl_0_14 br_0_14 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c14
+ bl_0_14 br_0_14 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c14
+ bl_0_14 br_0_14 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c14
+ bl_0_14 br_0_14 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c14
+ bl_0_14 br_0_14 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c14
+ bl_0_14 br_0_14 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c14
+ bl_0_14 br_0_14 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c14
+ bl_0_14 br_0_14 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c14
+ bl_0_14 br_0_14 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c14
+ bl_0_14 br_0_14 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c14
+ bl_0_14 br_0_14 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c14
+ bl_0_14 br_0_14 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c15
+ bl_0_15 br_0_15 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c15
+ bl_0_15 br_0_15 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c15
+ bl_0_15 br_0_15 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c15
+ bl_0_15 br_0_15 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c15
+ bl_0_15 br_0_15 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c15
+ bl_0_15 br_0_15 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c15
+ bl_0_15 br_0_15 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c15
+ bl_0_15 br_0_15 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c15
+ bl_0_15 br_0_15 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c15
+ bl_0_15 br_0_15 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c15
+ bl_0_15 br_0_15 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c15
+ bl_0_15 br_0_15 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c15
+ bl_0_15 br_0_15 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c15
+ bl_0_15 br_0_15 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c15
+ bl_0_15 br_0_15 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c15
+ bl_0_15 br_0_15 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c15
+ bl_0_15 br_0_15 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c15
+ bl_0_15 br_0_15 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c15
+ bl_0_15 br_0_15 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c15
+ bl_0_15 br_0_15 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c15
+ bl_0_15 br_0_15 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c15
+ bl_0_15 br_0_15 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c15
+ bl_0_15 br_0_15 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c15
+ bl_0_15 br_0_15 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c15
+ bl_0_15 br_0_15 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c15
+ bl_0_15 br_0_15 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c15
+ bl_0_15 br_0_15 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c15
+ bl_0_15 br_0_15 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c15
+ bl_0_15 br_0_15 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c15
+ bl_0_15 br_0_15 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c15
+ bl_0_15 br_0_15 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c15
+ bl_0_15 br_0_15 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c15
+ bl_0_15 br_0_15 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c15
+ bl_0_15 br_0_15 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c15
+ bl_0_15 br_0_15 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c15
+ bl_0_15 br_0_15 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c15
+ bl_0_15 br_0_15 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c15
+ bl_0_15 br_0_15 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c15
+ bl_0_15 br_0_15 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c15
+ bl_0_15 br_0_15 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c15
+ bl_0_15 br_0_15 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c15
+ bl_0_15 br_0_15 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c15
+ bl_0_15 br_0_15 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c15
+ bl_0_15 br_0_15 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c16
+ bl_0_16 br_0_16 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c16
+ bl_0_16 br_0_16 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c16
+ bl_0_16 br_0_16 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c16
+ bl_0_16 br_0_16 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c16
+ bl_0_16 br_0_16 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c16
+ bl_0_16 br_0_16 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c16
+ bl_0_16 br_0_16 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c16
+ bl_0_16 br_0_16 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c16
+ bl_0_16 br_0_16 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c16
+ bl_0_16 br_0_16 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c16
+ bl_0_16 br_0_16 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c16
+ bl_0_16 br_0_16 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c16
+ bl_0_16 br_0_16 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c16
+ bl_0_16 br_0_16 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c16
+ bl_0_16 br_0_16 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c16
+ bl_0_16 br_0_16 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c16
+ bl_0_16 br_0_16 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c16
+ bl_0_16 br_0_16 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c16
+ bl_0_16 br_0_16 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c16
+ bl_0_16 br_0_16 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c16
+ bl_0_16 br_0_16 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c16
+ bl_0_16 br_0_16 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c16
+ bl_0_16 br_0_16 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c16
+ bl_0_16 br_0_16 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c16
+ bl_0_16 br_0_16 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c16
+ bl_0_16 br_0_16 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c16
+ bl_0_16 br_0_16 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c16
+ bl_0_16 br_0_16 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c16
+ bl_0_16 br_0_16 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c16
+ bl_0_16 br_0_16 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c16
+ bl_0_16 br_0_16 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c16
+ bl_0_16 br_0_16 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c16
+ bl_0_16 br_0_16 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c16
+ bl_0_16 br_0_16 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c16
+ bl_0_16 br_0_16 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c16
+ bl_0_16 br_0_16 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c16
+ bl_0_16 br_0_16 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c16
+ bl_0_16 br_0_16 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c16
+ bl_0_16 br_0_16 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c16
+ bl_0_16 br_0_16 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c16
+ bl_0_16 br_0_16 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c16
+ bl_0_16 br_0_16 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c16
+ bl_0_16 br_0_16 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c16
+ bl_0_16 br_0_16 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c17
+ bl_0_17 br_0_17 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c17
+ bl_0_17 br_0_17 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c17
+ bl_0_17 br_0_17 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c17
+ bl_0_17 br_0_17 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c17
+ bl_0_17 br_0_17 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c17
+ bl_0_17 br_0_17 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c17
+ bl_0_17 br_0_17 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c17
+ bl_0_17 br_0_17 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c17
+ bl_0_17 br_0_17 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c17
+ bl_0_17 br_0_17 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c17
+ bl_0_17 br_0_17 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c17
+ bl_0_17 br_0_17 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c17
+ bl_0_17 br_0_17 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c17
+ bl_0_17 br_0_17 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c17
+ bl_0_17 br_0_17 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c17
+ bl_0_17 br_0_17 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c17
+ bl_0_17 br_0_17 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c17
+ bl_0_17 br_0_17 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c17
+ bl_0_17 br_0_17 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c17
+ bl_0_17 br_0_17 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c17
+ bl_0_17 br_0_17 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c17
+ bl_0_17 br_0_17 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c17
+ bl_0_17 br_0_17 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c17
+ bl_0_17 br_0_17 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c17
+ bl_0_17 br_0_17 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c17
+ bl_0_17 br_0_17 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c17
+ bl_0_17 br_0_17 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c17
+ bl_0_17 br_0_17 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c17
+ bl_0_17 br_0_17 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c17
+ bl_0_17 br_0_17 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c17
+ bl_0_17 br_0_17 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c17
+ bl_0_17 br_0_17 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c17
+ bl_0_17 br_0_17 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c17
+ bl_0_17 br_0_17 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c17
+ bl_0_17 br_0_17 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c17
+ bl_0_17 br_0_17 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c17
+ bl_0_17 br_0_17 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c17
+ bl_0_17 br_0_17 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c17
+ bl_0_17 br_0_17 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c17
+ bl_0_17 br_0_17 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c17
+ bl_0_17 br_0_17 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c17
+ bl_0_17 br_0_17 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c17
+ bl_0_17 br_0_17 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c17
+ bl_0_17 br_0_17 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c18
+ bl_0_18 br_0_18 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c18
+ bl_0_18 br_0_18 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c18
+ bl_0_18 br_0_18 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c18
+ bl_0_18 br_0_18 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c18
+ bl_0_18 br_0_18 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c18
+ bl_0_18 br_0_18 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c18
+ bl_0_18 br_0_18 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c18
+ bl_0_18 br_0_18 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c18
+ bl_0_18 br_0_18 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c18
+ bl_0_18 br_0_18 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c18
+ bl_0_18 br_0_18 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c18
+ bl_0_18 br_0_18 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c18
+ bl_0_18 br_0_18 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c18
+ bl_0_18 br_0_18 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c18
+ bl_0_18 br_0_18 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c18
+ bl_0_18 br_0_18 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c18
+ bl_0_18 br_0_18 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c18
+ bl_0_18 br_0_18 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c18
+ bl_0_18 br_0_18 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c18
+ bl_0_18 br_0_18 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c18
+ bl_0_18 br_0_18 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c18
+ bl_0_18 br_0_18 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c18
+ bl_0_18 br_0_18 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c18
+ bl_0_18 br_0_18 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c18
+ bl_0_18 br_0_18 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c18
+ bl_0_18 br_0_18 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c18
+ bl_0_18 br_0_18 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c18
+ bl_0_18 br_0_18 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c18
+ bl_0_18 br_0_18 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c18
+ bl_0_18 br_0_18 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c18
+ bl_0_18 br_0_18 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c18
+ bl_0_18 br_0_18 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c18
+ bl_0_18 br_0_18 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c18
+ bl_0_18 br_0_18 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c18
+ bl_0_18 br_0_18 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c18
+ bl_0_18 br_0_18 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c18
+ bl_0_18 br_0_18 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c18
+ bl_0_18 br_0_18 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c18
+ bl_0_18 br_0_18 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c18
+ bl_0_18 br_0_18 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c18
+ bl_0_18 br_0_18 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c18
+ bl_0_18 br_0_18 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c18
+ bl_0_18 br_0_18 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c18
+ bl_0_18 br_0_18 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c19
+ bl_0_19 br_0_19 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c19
+ bl_0_19 br_0_19 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c19
+ bl_0_19 br_0_19 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c19
+ bl_0_19 br_0_19 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c19
+ bl_0_19 br_0_19 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c19
+ bl_0_19 br_0_19 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c19
+ bl_0_19 br_0_19 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c19
+ bl_0_19 br_0_19 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c19
+ bl_0_19 br_0_19 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c19
+ bl_0_19 br_0_19 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c19
+ bl_0_19 br_0_19 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c19
+ bl_0_19 br_0_19 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c19
+ bl_0_19 br_0_19 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c19
+ bl_0_19 br_0_19 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c19
+ bl_0_19 br_0_19 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c19
+ bl_0_19 br_0_19 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c19
+ bl_0_19 br_0_19 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c19
+ bl_0_19 br_0_19 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c19
+ bl_0_19 br_0_19 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c19
+ bl_0_19 br_0_19 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c19
+ bl_0_19 br_0_19 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c19
+ bl_0_19 br_0_19 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c19
+ bl_0_19 br_0_19 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c19
+ bl_0_19 br_0_19 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c19
+ bl_0_19 br_0_19 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c19
+ bl_0_19 br_0_19 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c19
+ bl_0_19 br_0_19 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c19
+ bl_0_19 br_0_19 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c19
+ bl_0_19 br_0_19 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c19
+ bl_0_19 br_0_19 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c19
+ bl_0_19 br_0_19 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c19
+ bl_0_19 br_0_19 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c19
+ bl_0_19 br_0_19 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c19
+ bl_0_19 br_0_19 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c19
+ bl_0_19 br_0_19 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c19
+ bl_0_19 br_0_19 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c19
+ bl_0_19 br_0_19 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c19
+ bl_0_19 br_0_19 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c19
+ bl_0_19 br_0_19 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c19
+ bl_0_19 br_0_19 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c19
+ bl_0_19 br_0_19 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c19
+ bl_0_19 br_0_19 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c19
+ bl_0_19 br_0_19 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c19
+ bl_0_19 br_0_19 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c20
+ bl_0_20 br_0_20 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c20
+ bl_0_20 br_0_20 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c20
+ bl_0_20 br_0_20 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c20
+ bl_0_20 br_0_20 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c20
+ bl_0_20 br_0_20 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c20
+ bl_0_20 br_0_20 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c20
+ bl_0_20 br_0_20 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c20
+ bl_0_20 br_0_20 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c20
+ bl_0_20 br_0_20 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c20
+ bl_0_20 br_0_20 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c20
+ bl_0_20 br_0_20 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c20
+ bl_0_20 br_0_20 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c20
+ bl_0_20 br_0_20 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c20
+ bl_0_20 br_0_20 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c20
+ bl_0_20 br_0_20 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c20
+ bl_0_20 br_0_20 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c20
+ bl_0_20 br_0_20 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c20
+ bl_0_20 br_0_20 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c20
+ bl_0_20 br_0_20 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c20
+ bl_0_20 br_0_20 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c20
+ bl_0_20 br_0_20 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c20
+ bl_0_20 br_0_20 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c20
+ bl_0_20 br_0_20 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c20
+ bl_0_20 br_0_20 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c20
+ bl_0_20 br_0_20 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c20
+ bl_0_20 br_0_20 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c20
+ bl_0_20 br_0_20 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c20
+ bl_0_20 br_0_20 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c20
+ bl_0_20 br_0_20 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c20
+ bl_0_20 br_0_20 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c20
+ bl_0_20 br_0_20 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c20
+ bl_0_20 br_0_20 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c20
+ bl_0_20 br_0_20 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c20
+ bl_0_20 br_0_20 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c20
+ bl_0_20 br_0_20 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c20
+ bl_0_20 br_0_20 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c20
+ bl_0_20 br_0_20 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c20
+ bl_0_20 br_0_20 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c20
+ bl_0_20 br_0_20 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c20
+ bl_0_20 br_0_20 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c20
+ bl_0_20 br_0_20 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c20
+ bl_0_20 br_0_20 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c20
+ bl_0_20 br_0_20 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c20
+ bl_0_20 br_0_20 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c21
+ bl_0_21 br_0_21 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c21
+ bl_0_21 br_0_21 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c21
+ bl_0_21 br_0_21 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c21
+ bl_0_21 br_0_21 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c21
+ bl_0_21 br_0_21 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c21
+ bl_0_21 br_0_21 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c21
+ bl_0_21 br_0_21 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c21
+ bl_0_21 br_0_21 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c21
+ bl_0_21 br_0_21 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c21
+ bl_0_21 br_0_21 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c21
+ bl_0_21 br_0_21 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c21
+ bl_0_21 br_0_21 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c21
+ bl_0_21 br_0_21 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c21
+ bl_0_21 br_0_21 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c21
+ bl_0_21 br_0_21 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c21
+ bl_0_21 br_0_21 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c21
+ bl_0_21 br_0_21 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c21
+ bl_0_21 br_0_21 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c21
+ bl_0_21 br_0_21 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c21
+ bl_0_21 br_0_21 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c21
+ bl_0_21 br_0_21 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c21
+ bl_0_21 br_0_21 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c21
+ bl_0_21 br_0_21 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c21
+ bl_0_21 br_0_21 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c21
+ bl_0_21 br_0_21 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c21
+ bl_0_21 br_0_21 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c21
+ bl_0_21 br_0_21 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c21
+ bl_0_21 br_0_21 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c21
+ bl_0_21 br_0_21 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c21
+ bl_0_21 br_0_21 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c21
+ bl_0_21 br_0_21 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c21
+ bl_0_21 br_0_21 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c21
+ bl_0_21 br_0_21 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c21
+ bl_0_21 br_0_21 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c21
+ bl_0_21 br_0_21 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c21
+ bl_0_21 br_0_21 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c21
+ bl_0_21 br_0_21 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c21
+ bl_0_21 br_0_21 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c21
+ bl_0_21 br_0_21 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c21
+ bl_0_21 br_0_21 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c21
+ bl_0_21 br_0_21 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c21
+ bl_0_21 br_0_21 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c21
+ bl_0_21 br_0_21 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c21
+ bl_0_21 br_0_21 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c22
+ bl_0_22 br_0_22 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c22
+ bl_0_22 br_0_22 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c22
+ bl_0_22 br_0_22 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c22
+ bl_0_22 br_0_22 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c22
+ bl_0_22 br_0_22 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c22
+ bl_0_22 br_0_22 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c22
+ bl_0_22 br_0_22 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c22
+ bl_0_22 br_0_22 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c22
+ bl_0_22 br_0_22 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c22
+ bl_0_22 br_0_22 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c22
+ bl_0_22 br_0_22 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c22
+ bl_0_22 br_0_22 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c22
+ bl_0_22 br_0_22 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c22
+ bl_0_22 br_0_22 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c22
+ bl_0_22 br_0_22 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c22
+ bl_0_22 br_0_22 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c22
+ bl_0_22 br_0_22 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c22
+ bl_0_22 br_0_22 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c22
+ bl_0_22 br_0_22 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c22
+ bl_0_22 br_0_22 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c22
+ bl_0_22 br_0_22 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c22
+ bl_0_22 br_0_22 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c22
+ bl_0_22 br_0_22 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c22
+ bl_0_22 br_0_22 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c22
+ bl_0_22 br_0_22 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c22
+ bl_0_22 br_0_22 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c22
+ bl_0_22 br_0_22 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c22
+ bl_0_22 br_0_22 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c22
+ bl_0_22 br_0_22 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c22
+ bl_0_22 br_0_22 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c22
+ bl_0_22 br_0_22 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c22
+ bl_0_22 br_0_22 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c22
+ bl_0_22 br_0_22 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c22
+ bl_0_22 br_0_22 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c22
+ bl_0_22 br_0_22 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c22
+ bl_0_22 br_0_22 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c22
+ bl_0_22 br_0_22 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c22
+ bl_0_22 br_0_22 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c22
+ bl_0_22 br_0_22 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c22
+ bl_0_22 br_0_22 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c22
+ bl_0_22 br_0_22 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c22
+ bl_0_22 br_0_22 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c22
+ bl_0_22 br_0_22 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c22
+ bl_0_22 br_0_22 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c23
+ bl_0_23 br_0_23 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c23
+ bl_0_23 br_0_23 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c23
+ bl_0_23 br_0_23 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c23
+ bl_0_23 br_0_23 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c23
+ bl_0_23 br_0_23 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c23
+ bl_0_23 br_0_23 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c23
+ bl_0_23 br_0_23 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c23
+ bl_0_23 br_0_23 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c23
+ bl_0_23 br_0_23 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c23
+ bl_0_23 br_0_23 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c23
+ bl_0_23 br_0_23 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c23
+ bl_0_23 br_0_23 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c23
+ bl_0_23 br_0_23 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c23
+ bl_0_23 br_0_23 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c23
+ bl_0_23 br_0_23 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c23
+ bl_0_23 br_0_23 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c23
+ bl_0_23 br_0_23 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c23
+ bl_0_23 br_0_23 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c23
+ bl_0_23 br_0_23 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c23
+ bl_0_23 br_0_23 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c23
+ bl_0_23 br_0_23 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c23
+ bl_0_23 br_0_23 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c23
+ bl_0_23 br_0_23 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c23
+ bl_0_23 br_0_23 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c23
+ bl_0_23 br_0_23 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c23
+ bl_0_23 br_0_23 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c23
+ bl_0_23 br_0_23 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c23
+ bl_0_23 br_0_23 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c23
+ bl_0_23 br_0_23 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c23
+ bl_0_23 br_0_23 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c23
+ bl_0_23 br_0_23 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c23
+ bl_0_23 br_0_23 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c23
+ bl_0_23 br_0_23 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c23
+ bl_0_23 br_0_23 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c23
+ bl_0_23 br_0_23 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c23
+ bl_0_23 br_0_23 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c23
+ bl_0_23 br_0_23 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c23
+ bl_0_23 br_0_23 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c23
+ bl_0_23 br_0_23 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c23
+ bl_0_23 br_0_23 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c23
+ bl_0_23 br_0_23 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c23
+ bl_0_23 br_0_23 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c23
+ bl_0_23 br_0_23 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c23
+ bl_0_23 br_0_23 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c24
+ bl_0_24 br_0_24 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c24
+ bl_0_24 br_0_24 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c24
+ bl_0_24 br_0_24 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c24
+ bl_0_24 br_0_24 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c24
+ bl_0_24 br_0_24 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c24
+ bl_0_24 br_0_24 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c24
+ bl_0_24 br_0_24 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c24
+ bl_0_24 br_0_24 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c24
+ bl_0_24 br_0_24 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c24
+ bl_0_24 br_0_24 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c24
+ bl_0_24 br_0_24 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c24
+ bl_0_24 br_0_24 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c24
+ bl_0_24 br_0_24 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c24
+ bl_0_24 br_0_24 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c24
+ bl_0_24 br_0_24 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c24
+ bl_0_24 br_0_24 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c24
+ bl_0_24 br_0_24 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c24
+ bl_0_24 br_0_24 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c24
+ bl_0_24 br_0_24 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c24
+ bl_0_24 br_0_24 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c24
+ bl_0_24 br_0_24 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c24
+ bl_0_24 br_0_24 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c24
+ bl_0_24 br_0_24 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c24
+ bl_0_24 br_0_24 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c24
+ bl_0_24 br_0_24 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c24
+ bl_0_24 br_0_24 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c24
+ bl_0_24 br_0_24 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c24
+ bl_0_24 br_0_24 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c24
+ bl_0_24 br_0_24 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c24
+ bl_0_24 br_0_24 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c24
+ bl_0_24 br_0_24 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c24
+ bl_0_24 br_0_24 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c24
+ bl_0_24 br_0_24 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c24
+ bl_0_24 br_0_24 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c24
+ bl_0_24 br_0_24 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c24
+ bl_0_24 br_0_24 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c24
+ bl_0_24 br_0_24 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c24
+ bl_0_24 br_0_24 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c24
+ bl_0_24 br_0_24 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c24
+ bl_0_24 br_0_24 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c24
+ bl_0_24 br_0_24 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c24
+ bl_0_24 br_0_24 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c24
+ bl_0_24 br_0_24 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c24
+ bl_0_24 br_0_24 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c25
+ bl_0_25 br_0_25 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c25
+ bl_0_25 br_0_25 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c25
+ bl_0_25 br_0_25 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c25
+ bl_0_25 br_0_25 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c25
+ bl_0_25 br_0_25 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c25
+ bl_0_25 br_0_25 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c25
+ bl_0_25 br_0_25 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c25
+ bl_0_25 br_0_25 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c25
+ bl_0_25 br_0_25 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c25
+ bl_0_25 br_0_25 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c25
+ bl_0_25 br_0_25 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c25
+ bl_0_25 br_0_25 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c25
+ bl_0_25 br_0_25 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c25
+ bl_0_25 br_0_25 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c25
+ bl_0_25 br_0_25 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c25
+ bl_0_25 br_0_25 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c25
+ bl_0_25 br_0_25 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c25
+ bl_0_25 br_0_25 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c25
+ bl_0_25 br_0_25 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c25
+ bl_0_25 br_0_25 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c25
+ bl_0_25 br_0_25 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c25
+ bl_0_25 br_0_25 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c25
+ bl_0_25 br_0_25 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c25
+ bl_0_25 br_0_25 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c25
+ bl_0_25 br_0_25 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c25
+ bl_0_25 br_0_25 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c25
+ bl_0_25 br_0_25 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c25
+ bl_0_25 br_0_25 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c25
+ bl_0_25 br_0_25 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c25
+ bl_0_25 br_0_25 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c25
+ bl_0_25 br_0_25 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c25
+ bl_0_25 br_0_25 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c25
+ bl_0_25 br_0_25 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c25
+ bl_0_25 br_0_25 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c25
+ bl_0_25 br_0_25 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c25
+ bl_0_25 br_0_25 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c25
+ bl_0_25 br_0_25 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c25
+ bl_0_25 br_0_25 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c25
+ bl_0_25 br_0_25 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c25
+ bl_0_25 br_0_25 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c25
+ bl_0_25 br_0_25 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c25
+ bl_0_25 br_0_25 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c25
+ bl_0_25 br_0_25 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c25
+ bl_0_25 br_0_25 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c26
+ bl_0_26 br_0_26 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c26
+ bl_0_26 br_0_26 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c26
+ bl_0_26 br_0_26 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c26
+ bl_0_26 br_0_26 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c26
+ bl_0_26 br_0_26 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c26
+ bl_0_26 br_0_26 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c26
+ bl_0_26 br_0_26 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c26
+ bl_0_26 br_0_26 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c26
+ bl_0_26 br_0_26 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c26
+ bl_0_26 br_0_26 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c26
+ bl_0_26 br_0_26 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c26
+ bl_0_26 br_0_26 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c26
+ bl_0_26 br_0_26 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c26
+ bl_0_26 br_0_26 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c26
+ bl_0_26 br_0_26 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c26
+ bl_0_26 br_0_26 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c26
+ bl_0_26 br_0_26 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c26
+ bl_0_26 br_0_26 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c26
+ bl_0_26 br_0_26 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c26
+ bl_0_26 br_0_26 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c26
+ bl_0_26 br_0_26 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c26
+ bl_0_26 br_0_26 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c26
+ bl_0_26 br_0_26 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c26
+ bl_0_26 br_0_26 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c26
+ bl_0_26 br_0_26 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c26
+ bl_0_26 br_0_26 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c26
+ bl_0_26 br_0_26 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c26
+ bl_0_26 br_0_26 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c26
+ bl_0_26 br_0_26 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c26
+ bl_0_26 br_0_26 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c26
+ bl_0_26 br_0_26 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c26
+ bl_0_26 br_0_26 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c26
+ bl_0_26 br_0_26 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c26
+ bl_0_26 br_0_26 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c26
+ bl_0_26 br_0_26 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c26
+ bl_0_26 br_0_26 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c26
+ bl_0_26 br_0_26 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c26
+ bl_0_26 br_0_26 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c26
+ bl_0_26 br_0_26 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c26
+ bl_0_26 br_0_26 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c26
+ bl_0_26 br_0_26 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c26
+ bl_0_26 br_0_26 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c26
+ bl_0_26 br_0_26 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c26
+ bl_0_26 br_0_26 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c27
+ bl_0_27 br_0_27 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c27
+ bl_0_27 br_0_27 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c27
+ bl_0_27 br_0_27 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c27
+ bl_0_27 br_0_27 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c27
+ bl_0_27 br_0_27 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c27
+ bl_0_27 br_0_27 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c27
+ bl_0_27 br_0_27 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c27
+ bl_0_27 br_0_27 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c27
+ bl_0_27 br_0_27 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c27
+ bl_0_27 br_0_27 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c27
+ bl_0_27 br_0_27 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c27
+ bl_0_27 br_0_27 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c27
+ bl_0_27 br_0_27 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c27
+ bl_0_27 br_0_27 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c27
+ bl_0_27 br_0_27 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c27
+ bl_0_27 br_0_27 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c27
+ bl_0_27 br_0_27 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c27
+ bl_0_27 br_0_27 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c27
+ bl_0_27 br_0_27 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c27
+ bl_0_27 br_0_27 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c27
+ bl_0_27 br_0_27 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c27
+ bl_0_27 br_0_27 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c27
+ bl_0_27 br_0_27 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c27
+ bl_0_27 br_0_27 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c27
+ bl_0_27 br_0_27 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c27
+ bl_0_27 br_0_27 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c27
+ bl_0_27 br_0_27 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c27
+ bl_0_27 br_0_27 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c27
+ bl_0_27 br_0_27 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c27
+ bl_0_27 br_0_27 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c27
+ bl_0_27 br_0_27 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c27
+ bl_0_27 br_0_27 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c27
+ bl_0_27 br_0_27 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c27
+ bl_0_27 br_0_27 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c27
+ bl_0_27 br_0_27 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c27
+ bl_0_27 br_0_27 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c27
+ bl_0_27 br_0_27 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c27
+ bl_0_27 br_0_27 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c27
+ bl_0_27 br_0_27 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c27
+ bl_0_27 br_0_27 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c27
+ bl_0_27 br_0_27 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c27
+ bl_0_27 br_0_27 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c27
+ bl_0_27 br_0_27 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c27
+ bl_0_27 br_0_27 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c28
+ bl_0_28 br_0_28 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c28
+ bl_0_28 br_0_28 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c28
+ bl_0_28 br_0_28 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c28
+ bl_0_28 br_0_28 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c28
+ bl_0_28 br_0_28 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c28
+ bl_0_28 br_0_28 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c28
+ bl_0_28 br_0_28 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c28
+ bl_0_28 br_0_28 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c28
+ bl_0_28 br_0_28 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c28
+ bl_0_28 br_0_28 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c28
+ bl_0_28 br_0_28 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c28
+ bl_0_28 br_0_28 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c28
+ bl_0_28 br_0_28 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c28
+ bl_0_28 br_0_28 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c28
+ bl_0_28 br_0_28 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c28
+ bl_0_28 br_0_28 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c28
+ bl_0_28 br_0_28 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c28
+ bl_0_28 br_0_28 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c28
+ bl_0_28 br_0_28 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c28
+ bl_0_28 br_0_28 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c28
+ bl_0_28 br_0_28 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c28
+ bl_0_28 br_0_28 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c28
+ bl_0_28 br_0_28 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c28
+ bl_0_28 br_0_28 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c28
+ bl_0_28 br_0_28 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c28
+ bl_0_28 br_0_28 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c28
+ bl_0_28 br_0_28 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c28
+ bl_0_28 br_0_28 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c28
+ bl_0_28 br_0_28 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c28
+ bl_0_28 br_0_28 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c28
+ bl_0_28 br_0_28 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c28
+ bl_0_28 br_0_28 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c28
+ bl_0_28 br_0_28 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c28
+ bl_0_28 br_0_28 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c28
+ bl_0_28 br_0_28 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c28
+ bl_0_28 br_0_28 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c28
+ bl_0_28 br_0_28 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c28
+ bl_0_28 br_0_28 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c28
+ bl_0_28 br_0_28 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c28
+ bl_0_28 br_0_28 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c28
+ bl_0_28 br_0_28 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c28
+ bl_0_28 br_0_28 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c28
+ bl_0_28 br_0_28 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c28
+ bl_0_28 br_0_28 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c29
+ bl_0_29 br_0_29 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c29
+ bl_0_29 br_0_29 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c29
+ bl_0_29 br_0_29 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c29
+ bl_0_29 br_0_29 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c29
+ bl_0_29 br_0_29 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c29
+ bl_0_29 br_0_29 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c29
+ bl_0_29 br_0_29 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c29
+ bl_0_29 br_0_29 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c29
+ bl_0_29 br_0_29 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c29
+ bl_0_29 br_0_29 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c29
+ bl_0_29 br_0_29 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c29
+ bl_0_29 br_0_29 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c29
+ bl_0_29 br_0_29 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c29
+ bl_0_29 br_0_29 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c29
+ bl_0_29 br_0_29 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c29
+ bl_0_29 br_0_29 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c29
+ bl_0_29 br_0_29 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c29
+ bl_0_29 br_0_29 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c29
+ bl_0_29 br_0_29 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c29
+ bl_0_29 br_0_29 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c29
+ bl_0_29 br_0_29 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c29
+ bl_0_29 br_0_29 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c29
+ bl_0_29 br_0_29 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c29
+ bl_0_29 br_0_29 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c29
+ bl_0_29 br_0_29 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c29
+ bl_0_29 br_0_29 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c29
+ bl_0_29 br_0_29 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c29
+ bl_0_29 br_0_29 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c29
+ bl_0_29 br_0_29 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c29
+ bl_0_29 br_0_29 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c29
+ bl_0_29 br_0_29 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c29
+ bl_0_29 br_0_29 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c29
+ bl_0_29 br_0_29 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c29
+ bl_0_29 br_0_29 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c29
+ bl_0_29 br_0_29 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c29
+ bl_0_29 br_0_29 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c29
+ bl_0_29 br_0_29 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c29
+ bl_0_29 br_0_29 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c29
+ bl_0_29 br_0_29 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c29
+ bl_0_29 br_0_29 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c29
+ bl_0_29 br_0_29 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c29
+ bl_0_29 br_0_29 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c29
+ bl_0_29 br_0_29 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c29
+ bl_0_29 br_0_29 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c30
+ bl_0_30 br_0_30 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c30
+ bl_0_30 br_0_30 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c30
+ bl_0_30 br_0_30 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c30
+ bl_0_30 br_0_30 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c30
+ bl_0_30 br_0_30 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c30
+ bl_0_30 br_0_30 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c30
+ bl_0_30 br_0_30 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c30
+ bl_0_30 br_0_30 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c30
+ bl_0_30 br_0_30 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c30
+ bl_0_30 br_0_30 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c30
+ bl_0_30 br_0_30 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c30
+ bl_0_30 br_0_30 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c30
+ bl_0_30 br_0_30 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c30
+ bl_0_30 br_0_30 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c30
+ bl_0_30 br_0_30 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c30
+ bl_0_30 br_0_30 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c30
+ bl_0_30 br_0_30 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c30
+ bl_0_30 br_0_30 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c30
+ bl_0_30 br_0_30 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c30
+ bl_0_30 br_0_30 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c30
+ bl_0_30 br_0_30 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c30
+ bl_0_30 br_0_30 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c30
+ bl_0_30 br_0_30 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c30
+ bl_0_30 br_0_30 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c30
+ bl_0_30 br_0_30 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c30
+ bl_0_30 br_0_30 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c30
+ bl_0_30 br_0_30 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c30
+ bl_0_30 br_0_30 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c30
+ bl_0_30 br_0_30 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c30
+ bl_0_30 br_0_30 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c30
+ bl_0_30 br_0_30 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c30
+ bl_0_30 br_0_30 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c30
+ bl_0_30 br_0_30 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c30
+ bl_0_30 br_0_30 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c30
+ bl_0_30 br_0_30 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c30
+ bl_0_30 br_0_30 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c30
+ bl_0_30 br_0_30 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c30
+ bl_0_30 br_0_30 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c30
+ bl_0_30 br_0_30 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c30
+ bl_0_30 br_0_30 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c30
+ bl_0_30 br_0_30 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c30
+ bl_0_30 br_0_30 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c30
+ bl_0_30 br_0_30 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c30
+ bl_0_30 br_0_30 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c31
+ bl_0_31 br_0_31 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c31
+ bl_0_31 br_0_31 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c31
+ bl_0_31 br_0_31 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c31
+ bl_0_31 br_0_31 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c31
+ bl_0_31 br_0_31 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c31
+ bl_0_31 br_0_31 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c31
+ bl_0_31 br_0_31 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c31
+ bl_0_31 br_0_31 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c31
+ bl_0_31 br_0_31 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c31
+ bl_0_31 br_0_31 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c31
+ bl_0_31 br_0_31 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c31
+ bl_0_31 br_0_31 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c31
+ bl_0_31 br_0_31 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c31
+ bl_0_31 br_0_31 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c31
+ bl_0_31 br_0_31 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c31
+ bl_0_31 br_0_31 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c31
+ bl_0_31 br_0_31 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c31
+ bl_0_31 br_0_31 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c31
+ bl_0_31 br_0_31 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c31
+ bl_0_31 br_0_31 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c31
+ bl_0_31 br_0_31 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c31
+ bl_0_31 br_0_31 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c31
+ bl_0_31 br_0_31 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c31
+ bl_0_31 br_0_31 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c31
+ bl_0_31 br_0_31 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c31
+ bl_0_31 br_0_31 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c31
+ bl_0_31 br_0_31 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c31
+ bl_0_31 br_0_31 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c31
+ bl_0_31 br_0_31 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c31
+ bl_0_31 br_0_31 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c31
+ bl_0_31 br_0_31 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c31
+ bl_0_31 br_0_31 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c31
+ bl_0_31 br_0_31 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c31
+ bl_0_31 br_0_31 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c31
+ bl_0_31 br_0_31 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c31
+ bl_0_31 br_0_31 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c31
+ bl_0_31 br_0_31 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c31
+ bl_0_31 br_0_31 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c31
+ bl_0_31 br_0_31 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c31
+ bl_0_31 br_0_31 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c31
+ bl_0_31 br_0_31 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c31
+ bl_0_31 br_0_31 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c31
+ bl_0_31 br_0_31 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c31
+ bl_0_31 br_0_31 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c32
+ bl_0_32 br_0_32 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c32
+ bl_0_32 br_0_32 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c32
+ bl_0_32 br_0_32 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c32
+ bl_0_32 br_0_32 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c32
+ bl_0_32 br_0_32 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c32
+ bl_0_32 br_0_32 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c32
+ bl_0_32 br_0_32 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c32
+ bl_0_32 br_0_32 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c32
+ bl_0_32 br_0_32 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c32
+ bl_0_32 br_0_32 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c32
+ bl_0_32 br_0_32 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c32
+ bl_0_32 br_0_32 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c32
+ bl_0_32 br_0_32 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c32
+ bl_0_32 br_0_32 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c32
+ bl_0_32 br_0_32 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c32
+ bl_0_32 br_0_32 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c32
+ bl_0_32 br_0_32 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c32
+ bl_0_32 br_0_32 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c32
+ bl_0_32 br_0_32 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c32
+ bl_0_32 br_0_32 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c32
+ bl_0_32 br_0_32 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c32
+ bl_0_32 br_0_32 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c32
+ bl_0_32 br_0_32 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c32
+ bl_0_32 br_0_32 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c32
+ bl_0_32 br_0_32 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c32
+ bl_0_32 br_0_32 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c32
+ bl_0_32 br_0_32 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c32
+ bl_0_32 br_0_32 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c32
+ bl_0_32 br_0_32 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c32
+ bl_0_32 br_0_32 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c32
+ bl_0_32 br_0_32 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c32
+ bl_0_32 br_0_32 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c32
+ bl_0_32 br_0_32 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c32
+ bl_0_32 br_0_32 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c32
+ bl_0_32 br_0_32 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c32
+ bl_0_32 br_0_32 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c32
+ bl_0_32 br_0_32 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c32
+ bl_0_32 br_0_32 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c32
+ bl_0_32 br_0_32 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c32
+ bl_0_32 br_0_32 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c32
+ bl_0_32 br_0_32 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c32
+ bl_0_32 br_0_32 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c32
+ bl_0_32 br_0_32 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c32
+ bl_0_32 br_0_32 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c33
+ bl_0_33 br_0_33 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c33
+ bl_0_33 br_0_33 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c33
+ bl_0_33 br_0_33 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c33
+ bl_0_33 br_0_33 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c33
+ bl_0_33 br_0_33 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c33
+ bl_0_33 br_0_33 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c33
+ bl_0_33 br_0_33 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c33
+ bl_0_33 br_0_33 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c33
+ bl_0_33 br_0_33 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c33
+ bl_0_33 br_0_33 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c33
+ bl_0_33 br_0_33 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c33
+ bl_0_33 br_0_33 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c33
+ bl_0_33 br_0_33 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c33
+ bl_0_33 br_0_33 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c33
+ bl_0_33 br_0_33 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c33
+ bl_0_33 br_0_33 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c33
+ bl_0_33 br_0_33 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c33
+ bl_0_33 br_0_33 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c33
+ bl_0_33 br_0_33 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c33
+ bl_0_33 br_0_33 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c33
+ bl_0_33 br_0_33 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c33
+ bl_0_33 br_0_33 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c33
+ bl_0_33 br_0_33 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c33
+ bl_0_33 br_0_33 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c33
+ bl_0_33 br_0_33 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c33
+ bl_0_33 br_0_33 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c33
+ bl_0_33 br_0_33 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c33
+ bl_0_33 br_0_33 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c33
+ bl_0_33 br_0_33 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c33
+ bl_0_33 br_0_33 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c33
+ bl_0_33 br_0_33 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c33
+ bl_0_33 br_0_33 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c33
+ bl_0_33 br_0_33 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c33
+ bl_0_33 br_0_33 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c33
+ bl_0_33 br_0_33 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c33
+ bl_0_33 br_0_33 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c33
+ bl_0_33 br_0_33 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c33
+ bl_0_33 br_0_33 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c33
+ bl_0_33 br_0_33 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c33
+ bl_0_33 br_0_33 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c33
+ bl_0_33 br_0_33 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c33
+ bl_0_33 br_0_33 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c33
+ bl_0_33 br_0_33 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c33
+ bl_0_33 br_0_33 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c34
+ bl_0_34 br_0_34 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c34
+ bl_0_34 br_0_34 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c34
+ bl_0_34 br_0_34 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c34
+ bl_0_34 br_0_34 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c34
+ bl_0_34 br_0_34 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c34
+ bl_0_34 br_0_34 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c34
+ bl_0_34 br_0_34 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c34
+ bl_0_34 br_0_34 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c34
+ bl_0_34 br_0_34 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c34
+ bl_0_34 br_0_34 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c34
+ bl_0_34 br_0_34 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c34
+ bl_0_34 br_0_34 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c34
+ bl_0_34 br_0_34 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c34
+ bl_0_34 br_0_34 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c34
+ bl_0_34 br_0_34 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c34
+ bl_0_34 br_0_34 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c34
+ bl_0_34 br_0_34 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c34
+ bl_0_34 br_0_34 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c34
+ bl_0_34 br_0_34 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c34
+ bl_0_34 br_0_34 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c34
+ bl_0_34 br_0_34 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c34
+ bl_0_34 br_0_34 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c34
+ bl_0_34 br_0_34 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c34
+ bl_0_34 br_0_34 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c34
+ bl_0_34 br_0_34 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c34
+ bl_0_34 br_0_34 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c34
+ bl_0_34 br_0_34 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c34
+ bl_0_34 br_0_34 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c34
+ bl_0_34 br_0_34 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c34
+ bl_0_34 br_0_34 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c34
+ bl_0_34 br_0_34 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c34
+ bl_0_34 br_0_34 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c34
+ bl_0_34 br_0_34 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c34
+ bl_0_34 br_0_34 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c34
+ bl_0_34 br_0_34 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c34
+ bl_0_34 br_0_34 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c34
+ bl_0_34 br_0_34 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c34
+ bl_0_34 br_0_34 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c34
+ bl_0_34 br_0_34 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c34
+ bl_0_34 br_0_34 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c34
+ bl_0_34 br_0_34 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c34
+ bl_0_34 br_0_34 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c34
+ bl_0_34 br_0_34 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c34
+ bl_0_34 br_0_34 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c35
+ bl_0_35 br_0_35 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c35
+ bl_0_35 br_0_35 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c35
+ bl_0_35 br_0_35 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c35
+ bl_0_35 br_0_35 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c35
+ bl_0_35 br_0_35 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c35
+ bl_0_35 br_0_35 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c35
+ bl_0_35 br_0_35 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c35
+ bl_0_35 br_0_35 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c35
+ bl_0_35 br_0_35 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c35
+ bl_0_35 br_0_35 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c35
+ bl_0_35 br_0_35 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c35
+ bl_0_35 br_0_35 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c35
+ bl_0_35 br_0_35 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c35
+ bl_0_35 br_0_35 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c35
+ bl_0_35 br_0_35 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c35
+ bl_0_35 br_0_35 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c35
+ bl_0_35 br_0_35 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c35
+ bl_0_35 br_0_35 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c35
+ bl_0_35 br_0_35 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c35
+ bl_0_35 br_0_35 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c35
+ bl_0_35 br_0_35 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c35
+ bl_0_35 br_0_35 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c35
+ bl_0_35 br_0_35 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c35
+ bl_0_35 br_0_35 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c35
+ bl_0_35 br_0_35 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c35
+ bl_0_35 br_0_35 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c35
+ bl_0_35 br_0_35 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c35
+ bl_0_35 br_0_35 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c35
+ bl_0_35 br_0_35 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c35
+ bl_0_35 br_0_35 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c35
+ bl_0_35 br_0_35 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c35
+ bl_0_35 br_0_35 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c35
+ bl_0_35 br_0_35 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c35
+ bl_0_35 br_0_35 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c35
+ bl_0_35 br_0_35 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c35
+ bl_0_35 br_0_35 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c35
+ bl_0_35 br_0_35 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c35
+ bl_0_35 br_0_35 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c35
+ bl_0_35 br_0_35 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c35
+ bl_0_35 br_0_35 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c35
+ bl_0_35 br_0_35 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c35
+ bl_0_35 br_0_35 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c35
+ bl_0_35 br_0_35 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c35
+ bl_0_35 br_0_35 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c36
+ bl_0_36 br_0_36 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c36
+ bl_0_36 br_0_36 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c36
+ bl_0_36 br_0_36 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c36
+ bl_0_36 br_0_36 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c36
+ bl_0_36 br_0_36 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c36
+ bl_0_36 br_0_36 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c36
+ bl_0_36 br_0_36 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c36
+ bl_0_36 br_0_36 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c36
+ bl_0_36 br_0_36 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c36
+ bl_0_36 br_0_36 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c36
+ bl_0_36 br_0_36 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c36
+ bl_0_36 br_0_36 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c36
+ bl_0_36 br_0_36 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c36
+ bl_0_36 br_0_36 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c36
+ bl_0_36 br_0_36 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c36
+ bl_0_36 br_0_36 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c36
+ bl_0_36 br_0_36 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c36
+ bl_0_36 br_0_36 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c36
+ bl_0_36 br_0_36 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c36
+ bl_0_36 br_0_36 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c36
+ bl_0_36 br_0_36 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c36
+ bl_0_36 br_0_36 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c36
+ bl_0_36 br_0_36 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c36
+ bl_0_36 br_0_36 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c36
+ bl_0_36 br_0_36 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c36
+ bl_0_36 br_0_36 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c36
+ bl_0_36 br_0_36 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c36
+ bl_0_36 br_0_36 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c36
+ bl_0_36 br_0_36 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c36
+ bl_0_36 br_0_36 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c36
+ bl_0_36 br_0_36 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c36
+ bl_0_36 br_0_36 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c36
+ bl_0_36 br_0_36 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c36
+ bl_0_36 br_0_36 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c36
+ bl_0_36 br_0_36 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c36
+ bl_0_36 br_0_36 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c36
+ bl_0_36 br_0_36 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c36
+ bl_0_36 br_0_36 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c36
+ bl_0_36 br_0_36 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c36
+ bl_0_36 br_0_36 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c36
+ bl_0_36 br_0_36 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c36
+ bl_0_36 br_0_36 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c36
+ bl_0_36 br_0_36 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c36
+ bl_0_36 br_0_36 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c37
+ bl_0_37 br_0_37 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c37
+ bl_0_37 br_0_37 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c37
+ bl_0_37 br_0_37 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c37
+ bl_0_37 br_0_37 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c37
+ bl_0_37 br_0_37 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c37
+ bl_0_37 br_0_37 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c37
+ bl_0_37 br_0_37 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c37
+ bl_0_37 br_0_37 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c37
+ bl_0_37 br_0_37 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c37
+ bl_0_37 br_0_37 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c37
+ bl_0_37 br_0_37 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c37
+ bl_0_37 br_0_37 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c37
+ bl_0_37 br_0_37 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c37
+ bl_0_37 br_0_37 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c37
+ bl_0_37 br_0_37 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c37
+ bl_0_37 br_0_37 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c37
+ bl_0_37 br_0_37 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c37
+ bl_0_37 br_0_37 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c37
+ bl_0_37 br_0_37 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c37
+ bl_0_37 br_0_37 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c37
+ bl_0_37 br_0_37 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c37
+ bl_0_37 br_0_37 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c37
+ bl_0_37 br_0_37 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c37
+ bl_0_37 br_0_37 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c37
+ bl_0_37 br_0_37 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c37
+ bl_0_37 br_0_37 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c37
+ bl_0_37 br_0_37 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c37
+ bl_0_37 br_0_37 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c37
+ bl_0_37 br_0_37 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c37
+ bl_0_37 br_0_37 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c37
+ bl_0_37 br_0_37 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c37
+ bl_0_37 br_0_37 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c37
+ bl_0_37 br_0_37 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c37
+ bl_0_37 br_0_37 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c37
+ bl_0_37 br_0_37 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c37
+ bl_0_37 br_0_37 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c37
+ bl_0_37 br_0_37 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c37
+ bl_0_37 br_0_37 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c37
+ bl_0_37 br_0_37 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c37
+ bl_0_37 br_0_37 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c37
+ bl_0_37 br_0_37 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c37
+ bl_0_37 br_0_37 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c37
+ bl_0_37 br_0_37 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c37
+ bl_0_37 br_0_37 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c38
+ bl_0_38 br_0_38 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c38
+ bl_0_38 br_0_38 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c38
+ bl_0_38 br_0_38 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c38
+ bl_0_38 br_0_38 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c38
+ bl_0_38 br_0_38 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c38
+ bl_0_38 br_0_38 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c38
+ bl_0_38 br_0_38 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c38
+ bl_0_38 br_0_38 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c38
+ bl_0_38 br_0_38 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c38
+ bl_0_38 br_0_38 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c38
+ bl_0_38 br_0_38 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c38
+ bl_0_38 br_0_38 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c38
+ bl_0_38 br_0_38 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c38
+ bl_0_38 br_0_38 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c38
+ bl_0_38 br_0_38 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c38
+ bl_0_38 br_0_38 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c38
+ bl_0_38 br_0_38 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c38
+ bl_0_38 br_0_38 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c38
+ bl_0_38 br_0_38 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c38
+ bl_0_38 br_0_38 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c38
+ bl_0_38 br_0_38 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c38
+ bl_0_38 br_0_38 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c38
+ bl_0_38 br_0_38 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c38
+ bl_0_38 br_0_38 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c38
+ bl_0_38 br_0_38 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c38
+ bl_0_38 br_0_38 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c38
+ bl_0_38 br_0_38 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c38
+ bl_0_38 br_0_38 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c38
+ bl_0_38 br_0_38 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c38
+ bl_0_38 br_0_38 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c38
+ bl_0_38 br_0_38 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c38
+ bl_0_38 br_0_38 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c38
+ bl_0_38 br_0_38 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c38
+ bl_0_38 br_0_38 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c38
+ bl_0_38 br_0_38 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c38
+ bl_0_38 br_0_38 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c38
+ bl_0_38 br_0_38 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c38
+ bl_0_38 br_0_38 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c38
+ bl_0_38 br_0_38 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c38
+ bl_0_38 br_0_38 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c38
+ bl_0_38 br_0_38 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c38
+ bl_0_38 br_0_38 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c38
+ bl_0_38 br_0_38 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c38
+ bl_0_38 br_0_38 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c39
+ bl_0_39 br_0_39 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c39
+ bl_0_39 br_0_39 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c39
+ bl_0_39 br_0_39 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c39
+ bl_0_39 br_0_39 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c39
+ bl_0_39 br_0_39 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c39
+ bl_0_39 br_0_39 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c39
+ bl_0_39 br_0_39 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c39
+ bl_0_39 br_0_39 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c39
+ bl_0_39 br_0_39 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c39
+ bl_0_39 br_0_39 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c39
+ bl_0_39 br_0_39 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c39
+ bl_0_39 br_0_39 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c39
+ bl_0_39 br_0_39 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c39
+ bl_0_39 br_0_39 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c39
+ bl_0_39 br_0_39 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c39
+ bl_0_39 br_0_39 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c39
+ bl_0_39 br_0_39 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c39
+ bl_0_39 br_0_39 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c39
+ bl_0_39 br_0_39 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c39
+ bl_0_39 br_0_39 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c39
+ bl_0_39 br_0_39 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c39
+ bl_0_39 br_0_39 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c39
+ bl_0_39 br_0_39 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c39
+ bl_0_39 br_0_39 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c39
+ bl_0_39 br_0_39 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c39
+ bl_0_39 br_0_39 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c39
+ bl_0_39 br_0_39 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c39
+ bl_0_39 br_0_39 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c39
+ bl_0_39 br_0_39 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c39
+ bl_0_39 br_0_39 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c39
+ bl_0_39 br_0_39 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c39
+ bl_0_39 br_0_39 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c39
+ bl_0_39 br_0_39 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c39
+ bl_0_39 br_0_39 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c39
+ bl_0_39 br_0_39 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c39
+ bl_0_39 br_0_39 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c39
+ bl_0_39 br_0_39 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c39
+ bl_0_39 br_0_39 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c39
+ bl_0_39 br_0_39 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c39
+ bl_0_39 br_0_39 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c39
+ bl_0_39 br_0_39 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c39
+ bl_0_39 br_0_39 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c39
+ bl_0_39 br_0_39 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c39
+ bl_0_39 br_0_39 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c40
+ bl_0_40 br_0_40 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c40
+ bl_0_40 br_0_40 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c40
+ bl_0_40 br_0_40 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c40
+ bl_0_40 br_0_40 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c40
+ bl_0_40 br_0_40 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c40
+ bl_0_40 br_0_40 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c40
+ bl_0_40 br_0_40 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c40
+ bl_0_40 br_0_40 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c40
+ bl_0_40 br_0_40 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c40
+ bl_0_40 br_0_40 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c40
+ bl_0_40 br_0_40 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c40
+ bl_0_40 br_0_40 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c40
+ bl_0_40 br_0_40 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c40
+ bl_0_40 br_0_40 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c40
+ bl_0_40 br_0_40 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c40
+ bl_0_40 br_0_40 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c40
+ bl_0_40 br_0_40 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c40
+ bl_0_40 br_0_40 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c40
+ bl_0_40 br_0_40 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c40
+ bl_0_40 br_0_40 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c40
+ bl_0_40 br_0_40 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c40
+ bl_0_40 br_0_40 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c40
+ bl_0_40 br_0_40 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c40
+ bl_0_40 br_0_40 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c40
+ bl_0_40 br_0_40 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c40
+ bl_0_40 br_0_40 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c40
+ bl_0_40 br_0_40 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c40
+ bl_0_40 br_0_40 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c40
+ bl_0_40 br_0_40 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c40
+ bl_0_40 br_0_40 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c40
+ bl_0_40 br_0_40 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c40
+ bl_0_40 br_0_40 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c40
+ bl_0_40 br_0_40 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c40
+ bl_0_40 br_0_40 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c40
+ bl_0_40 br_0_40 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c40
+ bl_0_40 br_0_40 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c40
+ bl_0_40 br_0_40 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c40
+ bl_0_40 br_0_40 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c40
+ bl_0_40 br_0_40 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c40
+ bl_0_40 br_0_40 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c40
+ bl_0_40 br_0_40 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c40
+ bl_0_40 br_0_40 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c40
+ bl_0_40 br_0_40 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c40
+ bl_0_40 br_0_40 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c41
+ bl_0_41 br_0_41 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c41
+ bl_0_41 br_0_41 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c41
+ bl_0_41 br_0_41 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c41
+ bl_0_41 br_0_41 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c41
+ bl_0_41 br_0_41 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c41
+ bl_0_41 br_0_41 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c41
+ bl_0_41 br_0_41 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c41
+ bl_0_41 br_0_41 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c41
+ bl_0_41 br_0_41 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c41
+ bl_0_41 br_0_41 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c41
+ bl_0_41 br_0_41 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c41
+ bl_0_41 br_0_41 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c41
+ bl_0_41 br_0_41 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c41
+ bl_0_41 br_0_41 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c41
+ bl_0_41 br_0_41 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c41
+ bl_0_41 br_0_41 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c41
+ bl_0_41 br_0_41 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c41
+ bl_0_41 br_0_41 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c41
+ bl_0_41 br_0_41 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c41
+ bl_0_41 br_0_41 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c41
+ bl_0_41 br_0_41 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c41
+ bl_0_41 br_0_41 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c41
+ bl_0_41 br_0_41 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c41
+ bl_0_41 br_0_41 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c41
+ bl_0_41 br_0_41 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c41
+ bl_0_41 br_0_41 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c41
+ bl_0_41 br_0_41 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c41
+ bl_0_41 br_0_41 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c41
+ bl_0_41 br_0_41 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c41
+ bl_0_41 br_0_41 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c41
+ bl_0_41 br_0_41 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c41
+ bl_0_41 br_0_41 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c41
+ bl_0_41 br_0_41 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c41
+ bl_0_41 br_0_41 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c41
+ bl_0_41 br_0_41 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c41
+ bl_0_41 br_0_41 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c41
+ bl_0_41 br_0_41 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c41
+ bl_0_41 br_0_41 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c41
+ bl_0_41 br_0_41 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c41
+ bl_0_41 br_0_41 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c41
+ bl_0_41 br_0_41 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c41
+ bl_0_41 br_0_41 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c41
+ bl_0_41 br_0_41 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c41
+ bl_0_41 br_0_41 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c42
+ bl_0_42 br_0_42 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c42
+ bl_0_42 br_0_42 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c42
+ bl_0_42 br_0_42 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c42
+ bl_0_42 br_0_42 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c42
+ bl_0_42 br_0_42 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c42
+ bl_0_42 br_0_42 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c42
+ bl_0_42 br_0_42 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c42
+ bl_0_42 br_0_42 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c42
+ bl_0_42 br_0_42 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c42
+ bl_0_42 br_0_42 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c42
+ bl_0_42 br_0_42 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c42
+ bl_0_42 br_0_42 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c42
+ bl_0_42 br_0_42 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c42
+ bl_0_42 br_0_42 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c42
+ bl_0_42 br_0_42 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c42
+ bl_0_42 br_0_42 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c42
+ bl_0_42 br_0_42 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c42
+ bl_0_42 br_0_42 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c42
+ bl_0_42 br_0_42 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c42
+ bl_0_42 br_0_42 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c42
+ bl_0_42 br_0_42 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c42
+ bl_0_42 br_0_42 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c42
+ bl_0_42 br_0_42 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c42
+ bl_0_42 br_0_42 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c42
+ bl_0_42 br_0_42 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c42
+ bl_0_42 br_0_42 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c42
+ bl_0_42 br_0_42 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c42
+ bl_0_42 br_0_42 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c42
+ bl_0_42 br_0_42 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c42
+ bl_0_42 br_0_42 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c42
+ bl_0_42 br_0_42 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c42
+ bl_0_42 br_0_42 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c42
+ bl_0_42 br_0_42 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c42
+ bl_0_42 br_0_42 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c42
+ bl_0_42 br_0_42 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c42
+ bl_0_42 br_0_42 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c42
+ bl_0_42 br_0_42 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c42
+ bl_0_42 br_0_42 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c42
+ bl_0_42 br_0_42 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c42
+ bl_0_42 br_0_42 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c42
+ bl_0_42 br_0_42 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c42
+ bl_0_42 br_0_42 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c42
+ bl_0_42 br_0_42 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c42
+ bl_0_42 br_0_42 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c43
+ bl_0_43 br_0_43 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c43
+ bl_0_43 br_0_43 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c43
+ bl_0_43 br_0_43 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c43
+ bl_0_43 br_0_43 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c43
+ bl_0_43 br_0_43 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c43
+ bl_0_43 br_0_43 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c43
+ bl_0_43 br_0_43 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c43
+ bl_0_43 br_0_43 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c43
+ bl_0_43 br_0_43 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c43
+ bl_0_43 br_0_43 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c43
+ bl_0_43 br_0_43 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c43
+ bl_0_43 br_0_43 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c43
+ bl_0_43 br_0_43 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c43
+ bl_0_43 br_0_43 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c43
+ bl_0_43 br_0_43 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c43
+ bl_0_43 br_0_43 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c43
+ bl_0_43 br_0_43 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c43
+ bl_0_43 br_0_43 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c43
+ bl_0_43 br_0_43 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c43
+ bl_0_43 br_0_43 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c43
+ bl_0_43 br_0_43 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c43
+ bl_0_43 br_0_43 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c43
+ bl_0_43 br_0_43 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c43
+ bl_0_43 br_0_43 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c43
+ bl_0_43 br_0_43 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c43
+ bl_0_43 br_0_43 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c43
+ bl_0_43 br_0_43 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c43
+ bl_0_43 br_0_43 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c43
+ bl_0_43 br_0_43 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c43
+ bl_0_43 br_0_43 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c43
+ bl_0_43 br_0_43 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c43
+ bl_0_43 br_0_43 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c43
+ bl_0_43 br_0_43 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c43
+ bl_0_43 br_0_43 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c43
+ bl_0_43 br_0_43 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c43
+ bl_0_43 br_0_43 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c43
+ bl_0_43 br_0_43 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c43
+ bl_0_43 br_0_43 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c43
+ bl_0_43 br_0_43 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c43
+ bl_0_43 br_0_43 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c43
+ bl_0_43 br_0_43 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c43
+ bl_0_43 br_0_43 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c43
+ bl_0_43 br_0_43 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c43
+ bl_0_43 br_0_43 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c44
+ bl_0_44 br_0_44 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c44
+ bl_0_44 br_0_44 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c44
+ bl_0_44 br_0_44 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c44
+ bl_0_44 br_0_44 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c44
+ bl_0_44 br_0_44 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c44
+ bl_0_44 br_0_44 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c44
+ bl_0_44 br_0_44 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c44
+ bl_0_44 br_0_44 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c44
+ bl_0_44 br_0_44 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c44
+ bl_0_44 br_0_44 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c44
+ bl_0_44 br_0_44 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c44
+ bl_0_44 br_0_44 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c44
+ bl_0_44 br_0_44 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c44
+ bl_0_44 br_0_44 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c44
+ bl_0_44 br_0_44 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c44
+ bl_0_44 br_0_44 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c44
+ bl_0_44 br_0_44 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c44
+ bl_0_44 br_0_44 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c44
+ bl_0_44 br_0_44 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c44
+ bl_0_44 br_0_44 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c44
+ bl_0_44 br_0_44 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c44
+ bl_0_44 br_0_44 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c44
+ bl_0_44 br_0_44 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c44
+ bl_0_44 br_0_44 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c44
+ bl_0_44 br_0_44 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c44
+ bl_0_44 br_0_44 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c44
+ bl_0_44 br_0_44 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c44
+ bl_0_44 br_0_44 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c44
+ bl_0_44 br_0_44 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c44
+ bl_0_44 br_0_44 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c44
+ bl_0_44 br_0_44 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c44
+ bl_0_44 br_0_44 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c44
+ bl_0_44 br_0_44 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c44
+ bl_0_44 br_0_44 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c44
+ bl_0_44 br_0_44 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c44
+ bl_0_44 br_0_44 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c44
+ bl_0_44 br_0_44 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c44
+ bl_0_44 br_0_44 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c44
+ bl_0_44 br_0_44 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c44
+ bl_0_44 br_0_44 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c44
+ bl_0_44 br_0_44 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c44
+ bl_0_44 br_0_44 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c44
+ bl_0_44 br_0_44 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c44
+ bl_0_44 br_0_44 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c45
+ bl_0_45 br_0_45 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c45
+ bl_0_45 br_0_45 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c45
+ bl_0_45 br_0_45 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c45
+ bl_0_45 br_0_45 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c45
+ bl_0_45 br_0_45 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c45
+ bl_0_45 br_0_45 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c45
+ bl_0_45 br_0_45 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c45
+ bl_0_45 br_0_45 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c45
+ bl_0_45 br_0_45 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c45
+ bl_0_45 br_0_45 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c45
+ bl_0_45 br_0_45 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c45
+ bl_0_45 br_0_45 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c45
+ bl_0_45 br_0_45 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c45
+ bl_0_45 br_0_45 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c45
+ bl_0_45 br_0_45 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c45
+ bl_0_45 br_0_45 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c45
+ bl_0_45 br_0_45 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c45
+ bl_0_45 br_0_45 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c45
+ bl_0_45 br_0_45 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c45
+ bl_0_45 br_0_45 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c45
+ bl_0_45 br_0_45 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c45
+ bl_0_45 br_0_45 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c45
+ bl_0_45 br_0_45 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c45
+ bl_0_45 br_0_45 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c45
+ bl_0_45 br_0_45 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c45
+ bl_0_45 br_0_45 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c45
+ bl_0_45 br_0_45 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c45
+ bl_0_45 br_0_45 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c45
+ bl_0_45 br_0_45 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c45
+ bl_0_45 br_0_45 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c45
+ bl_0_45 br_0_45 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c45
+ bl_0_45 br_0_45 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c45
+ bl_0_45 br_0_45 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c45
+ bl_0_45 br_0_45 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c45
+ bl_0_45 br_0_45 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c45
+ bl_0_45 br_0_45 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c45
+ bl_0_45 br_0_45 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c45
+ bl_0_45 br_0_45 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c45
+ bl_0_45 br_0_45 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c45
+ bl_0_45 br_0_45 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c45
+ bl_0_45 br_0_45 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c45
+ bl_0_45 br_0_45 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c45
+ bl_0_45 br_0_45 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c45
+ bl_0_45 br_0_45 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c46
+ bl_0_46 br_0_46 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c46
+ bl_0_46 br_0_46 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c46
+ bl_0_46 br_0_46 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c46
+ bl_0_46 br_0_46 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c46
+ bl_0_46 br_0_46 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c46
+ bl_0_46 br_0_46 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c46
+ bl_0_46 br_0_46 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c46
+ bl_0_46 br_0_46 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c46
+ bl_0_46 br_0_46 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c46
+ bl_0_46 br_0_46 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c46
+ bl_0_46 br_0_46 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c46
+ bl_0_46 br_0_46 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c46
+ bl_0_46 br_0_46 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c46
+ bl_0_46 br_0_46 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c46
+ bl_0_46 br_0_46 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c46
+ bl_0_46 br_0_46 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c46
+ bl_0_46 br_0_46 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c46
+ bl_0_46 br_0_46 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c46
+ bl_0_46 br_0_46 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c46
+ bl_0_46 br_0_46 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c46
+ bl_0_46 br_0_46 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c46
+ bl_0_46 br_0_46 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c46
+ bl_0_46 br_0_46 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c46
+ bl_0_46 br_0_46 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c46
+ bl_0_46 br_0_46 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c46
+ bl_0_46 br_0_46 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c46
+ bl_0_46 br_0_46 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c46
+ bl_0_46 br_0_46 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c46
+ bl_0_46 br_0_46 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c46
+ bl_0_46 br_0_46 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c46
+ bl_0_46 br_0_46 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c46
+ bl_0_46 br_0_46 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c46
+ bl_0_46 br_0_46 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c46
+ bl_0_46 br_0_46 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c46
+ bl_0_46 br_0_46 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c46
+ bl_0_46 br_0_46 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c46
+ bl_0_46 br_0_46 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c46
+ bl_0_46 br_0_46 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c46
+ bl_0_46 br_0_46 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c46
+ bl_0_46 br_0_46 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c46
+ bl_0_46 br_0_46 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c46
+ bl_0_46 br_0_46 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c46
+ bl_0_46 br_0_46 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c46
+ bl_0_46 br_0_46 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c47
+ bl_0_47 br_0_47 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c47
+ bl_0_47 br_0_47 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c47
+ bl_0_47 br_0_47 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c47
+ bl_0_47 br_0_47 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c47
+ bl_0_47 br_0_47 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c47
+ bl_0_47 br_0_47 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c47
+ bl_0_47 br_0_47 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c47
+ bl_0_47 br_0_47 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c47
+ bl_0_47 br_0_47 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c47
+ bl_0_47 br_0_47 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c47
+ bl_0_47 br_0_47 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c47
+ bl_0_47 br_0_47 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c47
+ bl_0_47 br_0_47 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c47
+ bl_0_47 br_0_47 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c47
+ bl_0_47 br_0_47 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c47
+ bl_0_47 br_0_47 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c47
+ bl_0_47 br_0_47 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c47
+ bl_0_47 br_0_47 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c47
+ bl_0_47 br_0_47 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c47
+ bl_0_47 br_0_47 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c47
+ bl_0_47 br_0_47 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c47
+ bl_0_47 br_0_47 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c47
+ bl_0_47 br_0_47 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c47
+ bl_0_47 br_0_47 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c47
+ bl_0_47 br_0_47 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c47
+ bl_0_47 br_0_47 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c47
+ bl_0_47 br_0_47 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c47
+ bl_0_47 br_0_47 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c47
+ bl_0_47 br_0_47 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c47
+ bl_0_47 br_0_47 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c47
+ bl_0_47 br_0_47 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c47
+ bl_0_47 br_0_47 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c47
+ bl_0_47 br_0_47 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c47
+ bl_0_47 br_0_47 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c47
+ bl_0_47 br_0_47 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c47
+ bl_0_47 br_0_47 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c47
+ bl_0_47 br_0_47 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c47
+ bl_0_47 br_0_47 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c47
+ bl_0_47 br_0_47 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c47
+ bl_0_47 br_0_47 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c47
+ bl_0_47 br_0_47 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c47
+ bl_0_47 br_0_47 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c47
+ bl_0_47 br_0_47 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c47
+ bl_0_47 br_0_47 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c48
+ bl_0_48 br_0_48 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c48
+ bl_0_48 br_0_48 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c48
+ bl_0_48 br_0_48 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c48
+ bl_0_48 br_0_48 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c48
+ bl_0_48 br_0_48 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c48
+ bl_0_48 br_0_48 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c48
+ bl_0_48 br_0_48 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c48
+ bl_0_48 br_0_48 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c48
+ bl_0_48 br_0_48 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c48
+ bl_0_48 br_0_48 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c48
+ bl_0_48 br_0_48 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c48
+ bl_0_48 br_0_48 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c48
+ bl_0_48 br_0_48 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c48
+ bl_0_48 br_0_48 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c48
+ bl_0_48 br_0_48 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c48
+ bl_0_48 br_0_48 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c48
+ bl_0_48 br_0_48 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c48
+ bl_0_48 br_0_48 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c48
+ bl_0_48 br_0_48 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c48
+ bl_0_48 br_0_48 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c48
+ bl_0_48 br_0_48 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c48
+ bl_0_48 br_0_48 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c48
+ bl_0_48 br_0_48 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c48
+ bl_0_48 br_0_48 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c48
+ bl_0_48 br_0_48 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c48
+ bl_0_48 br_0_48 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c48
+ bl_0_48 br_0_48 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c48
+ bl_0_48 br_0_48 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c48
+ bl_0_48 br_0_48 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c48
+ bl_0_48 br_0_48 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c48
+ bl_0_48 br_0_48 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c48
+ bl_0_48 br_0_48 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c48
+ bl_0_48 br_0_48 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c48
+ bl_0_48 br_0_48 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c48
+ bl_0_48 br_0_48 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c48
+ bl_0_48 br_0_48 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c48
+ bl_0_48 br_0_48 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c48
+ bl_0_48 br_0_48 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c48
+ bl_0_48 br_0_48 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c48
+ bl_0_48 br_0_48 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c48
+ bl_0_48 br_0_48 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c48
+ bl_0_48 br_0_48 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c48
+ bl_0_48 br_0_48 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c48
+ bl_0_48 br_0_48 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c49
+ bl_0_49 br_0_49 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c49
+ bl_0_49 br_0_49 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c49
+ bl_0_49 br_0_49 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c49
+ bl_0_49 br_0_49 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c49
+ bl_0_49 br_0_49 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c49
+ bl_0_49 br_0_49 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c49
+ bl_0_49 br_0_49 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c49
+ bl_0_49 br_0_49 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c49
+ bl_0_49 br_0_49 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c49
+ bl_0_49 br_0_49 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c49
+ bl_0_49 br_0_49 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c49
+ bl_0_49 br_0_49 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c49
+ bl_0_49 br_0_49 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c49
+ bl_0_49 br_0_49 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c49
+ bl_0_49 br_0_49 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c49
+ bl_0_49 br_0_49 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c49
+ bl_0_49 br_0_49 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c49
+ bl_0_49 br_0_49 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c49
+ bl_0_49 br_0_49 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c49
+ bl_0_49 br_0_49 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c49
+ bl_0_49 br_0_49 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c49
+ bl_0_49 br_0_49 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c49
+ bl_0_49 br_0_49 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c49
+ bl_0_49 br_0_49 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c49
+ bl_0_49 br_0_49 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c49
+ bl_0_49 br_0_49 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c49
+ bl_0_49 br_0_49 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c49
+ bl_0_49 br_0_49 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c49
+ bl_0_49 br_0_49 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c49
+ bl_0_49 br_0_49 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c49
+ bl_0_49 br_0_49 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c49
+ bl_0_49 br_0_49 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c49
+ bl_0_49 br_0_49 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c49
+ bl_0_49 br_0_49 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c49
+ bl_0_49 br_0_49 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c49
+ bl_0_49 br_0_49 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c49
+ bl_0_49 br_0_49 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c49
+ bl_0_49 br_0_49 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c49
+ bl_0_49 br_0_49 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c49
+ bl_0_49 br_0_49 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c49
+ bl_0_49 br_0_49 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c49
+ bl_0_49 br_0_49 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c49
+ bl_0_49 br_0_49 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c49
+ bl_0_49 br_0_49 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c50
+ bl_0_50 br_0_50 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c50
+ bl_0_50 br_0_50 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c50
+ bl_0_50 br_0_50 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c50
+ bl_0_50 br_0_50 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c50
+ bl_0_50 br_0_50 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c50
+ bl_0_50 br_0_50 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c50
+ bl_0_50 br_0_50 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c50
+ bl_0_50 br_0_50 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c50
+ bl_0_50 br_0_50 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c50
+ bl_0_50 br_0_50 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c50
+ bl_0_50 br_0_50 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c50
+ bl_0_50 br_0_50 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c50
+ bl_0_50 br_0_50 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c50
+ bl_0_50 br_0_50 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c50
+ bl_0_50 br_0_50 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c50
+ bl_0_50 br_0_50 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c50
+ bl_0_50 br_0_50 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c50
+ bl_0_50 br_0_50 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c50
+ bl_0_50 br_0_50 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c50
+ bl_0_50 br_0_50 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c50
+ bl_0_50 br_0_50 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c50
+ bl_0_50 br_0_50 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c50
+ bl_0_50 br_0_50 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c50
+ bl_0_50 br_0_50 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c50
+ bl_0_50 br_0_50 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c50
+ bl_0_50 br_0_50 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c50
+ bl_0_50 br_0_50 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c50
+ bl_0_50 br_0_50 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c50
+ bl_0_50 br_0_50 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c50
+ bl_0_50 br_0_50 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c50
+ bl_0_50 br_0_50 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c50
+ bl_0_50 br_0_50 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c50
+ bl_0_50 br_0_50 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c50
+ bl_0_50 br_0_50 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c50
+ bl_0_50 br_0_50 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c50
+ bl_0_50 br_0_50 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c50
+ bl_0_50 br_0_50 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c50
+ bl_0_50 br_0_50 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c50
+ bl_0_50 br_0_50 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c50
+ bl_0_50 br_0_50 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c50
+ bl_0_50 br_0_50 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c50
+ bl_0_50 br_0_50 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c50
+ bl_0_50 br_0_50 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c50
+ bl_0_50 br_0_50 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c51
+ bl_0_51 br_0_51 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c51
+ bl_0_51 br_0_51 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c51
+ bl_0_51 br_0_51 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c51
+ bl_0_51 br_0_51 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c51
+ bl_0_51 br_0_51 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c51
+ bl_0_51 br_0_51 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c51
+ bl_0_51 br_0_51 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c51
+ bl_0_51 br_0_51 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c51
+ bl_0_51 br_0_51 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c51
+ bl_0_51 br_0_51 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c51
+ bl_0_51 br_0_51 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c51
+ bl_0_51 br_0_51 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c51
+ bl_0_51 br_0_51 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c51
+ bl_0_51 br_0_51 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c51
+ bl_0_51 br_0_51 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c51
+ bl_0_51 br_0_51 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c51
+ bl_0_51 br_0_51 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c51
+ bl_0_51 br_0_51 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c51
+ bl_0_51 br_0_51 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c51
+ bl_0_51 br_0_51 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c51
+ bl_0_51 br_0_51 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c51
+ bl_0_51 br_0_51 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c51
+ bl_0_51 br_0_51 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c51
+ bl_0_51 br_0_51 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c51
+ bl_0_51 br_0_51 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c51
+ bl_0_51 br_0_51 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c51
+ bl_0_51 br_0_51 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c51
+ bl_0_51 br_0_51 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c51
+ bl_0_51 br_0_51 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c51
+ bl_0_51 br_0_51 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c51
+ bl_0_51 br_0_51 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c51
+ bl_0_51 br_0_51 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c51
+ bl_0_51 br_0_51 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c51
+ bl_0_51 br_0_51 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c51
+ bl_0_51 br_0_51 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c51
+ bl_0_51 br_0_51 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c51
+ bl_0_51 br_0_51 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c51
+ bl_0_51 br_0_51 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c51
+ bl_0_51 br_0_51 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c51
+ bl_0_51 br_0_51 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c51
+ bl_0_51 br_0_51 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c51
+ bl_0_51 br_0_51 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c51
+ bl_0_51 br_0_51 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c51
+ bl_0_51 br_0_51 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c52
+ bl_0_52 br_0_52 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c52
+ bl_0_52 br_0_52 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c52
+ bl_0_52 br_0_52 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c52
+ bl_0_52 br_0_52 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c52
+ bl_0_52 br_0_52 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c52
+ bl_0_52 br_0_52 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c52
+ bl_0_52 br_0_52 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c52
+ bl_0_52 br_0_52 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c52
+ bl_0_52 br_0_52 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c52
+ bl_0_52 br_0_52 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c52
+ bl_0_52 br_0_52 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c52
+ bl_0_52 br_0_52 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c52
+ bl_0_52 br_0_52 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c52
+ bl_0_52 br_0_52 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c52
+ bl_0_52 br_0_52 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c52
+ bl_0_52 br_0_52 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c52
+ bl_0_52 br_0_52 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c52
+ bl_0_52 br_0_52 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c52
+ bl_0_52 br_0_52 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c52
+ bl_0_52 br_0_52 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c52
+ bl_0_52 br_0_52 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c52
+ bl_0_52 br_0_52 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c52
+ bl_0_52 br_0_52 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c52
+ bl_0_52 br_0_52 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c52
+ bl_0_52 br_0_52 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c52
+ bl_0_52 br_0_52 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c52
+ bl_0_52 br_0_52 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c52
+ bl_0_52 br_0_52 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c52
+ bl_0_52 br_0_52 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c52
+ bl_0_52 br_0_52 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c52
+ bl_0_52 br_0_52 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c52
+ bl_0_52 br_0_52 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c52
+ bl_0_52 br_0_52 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c52
+ bl_0_52 br_0_52 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c52
+ bl_0_52 br_0_52 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c52
+ bl_0_52 br_0_52 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c52
+ bl_0_52 br_0_52 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c52
+ bl_0_52 br_0_52 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c52
+ bl_0_52 br_0_52 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c52
+ bl_0_52 br_0_52 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c52
+ bl_0_52 br_0_52 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c52
+ bl_0_52 br_0_52 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c52
+ bl_0_52 br_0_52 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c52
+ bl_0_52 br_0_52 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c53
+ bl_0_53 br_0_53 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c53
+ bl_0_53 br_0_53 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c53
+ bl_0_53 br_0_53 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c53
+ bl_0_53 br_0_53 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c53
+ bl_0_53 br_0_53 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c53
+ bl_0_53 br_0_53 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c53
+ bl_0_53 br_0_53 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c53
+ bl_0_53 br_0_53 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c53
+ bl_0_53 br_0_53 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c53
+ bl_0_53 br_0_53 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c53
+ bl_0_53 br_0_53 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c53
+ bl_0_53 br_0_53 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c53
+ bl_0_53 br_0_53 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c53
+ bl_0_53 br_0_53 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c53
+ bl_0_53 br_0_53 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c53
+ bl_0_53 br_0_53 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c53
+ bl_0_53 br_0_53 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c53
+ bl_0_53 br_0_53 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c53
+ bl_0_53 br_0_53 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c53
+ bl_0_53 br_0_53 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c53
+ bl_0_53 br_0_53 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c53
+ bl_0_53 br_0_53 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c53
+ bl_0_53 br_0_53 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c53
+ bl_0_53 br_0_53 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c53
+ bl_0_53 br_0_53 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c53
+ bl_0_53 br_0_53 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c53
+ bl_0_53 br_0_53 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c53
+ bl_0_53 br_0_53 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c53
+ bl_0_53 br_0_53 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c53
+ bl_0_53 br_0_53 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c53
+ bl_0_53 br_0_53 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c53
+ bl_0_53 br_0_53 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c53
+ bl_0_53 br_0_53 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c53
+ bl_0_53 br_0_53 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c53
+ bl_0_53 br_0_53 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c53
+ bl_0_53 br_0_53 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c53
+ bl_0_53 br_0_53 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c53
+ bl_0_53 br_0_53 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c53
+ bl_0_53 br_0_53 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c53
+ bl_0_53 br_0_53 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c53
+ bl_0_53 br_0_53 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c53
+ bl_0_53 br_0_53 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c53
+ bl_0_53 br_0_53 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c53
+ bl_0_53 br_0_53 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c54
+ bl_0_54 br_0_54 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c54
+ bl_0_54 br_0_54 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c54
+ bl_0_54 br_0_54 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c54
+ bl_0_54 br_0_54 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c54
+ bl_0_54 br_0_54 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c54
+ bl_0_54 br_0_54 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c54
+ bl_0_54 br_0_54 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c54
+ bl_0_54 br_0_54 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c54
+ bl_0_54 br_0_54 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c54
+ bl_0_54 br_0_54 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c54
+ bl_0_54 br_0_54 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c54
+ bl_0_54 br_0_54 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c54
+ bl_0_54 br_0_54 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c54
+ bl_0_54 br_0_54 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c54
+ bl_0_54 br_0_54 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c54
+ bl_0_54 br_0_54 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c54
+ bl_0_54 br_0_54 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c54
+ bl_0_54 br_0_54 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c54
+ bl_0_54 br_0_54 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c54
+ bl_0_54 br_0_54 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c54
+ bl_0_54 br_0_54 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c54
+ bl_0_54 br_0_54 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c54
+ bl_0_54 br_0_54 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c54
+ bl_0_54 br_0_54 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c54
+ bl_0_54 br_0_54 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c54
+ bl_0_54 br_0_54 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c54
+ bl_0_54 br_0_54 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c54
+ bl_0_54 br_0_54 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c54
+ bl_0_54 br_0_54 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c54
+ bl_0_54 br_0_54 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c54
+ bl_0_54 br_0_54 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c54
+ bl_0_54 br_0_54 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c54
+ bl_0_54 br_0_54 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c54
+ bl_0_54 br_0_54 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c54
+ bl_0_54 br_0_54 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c54
+ bl_0_54 br_0_54 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c54
+ bl_0_54 br_0_54 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c54
+ bl_0_54 br_0_54 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c54
+ bl_0_54 br_0_54 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c54
+ bl_0_54 br_0_54 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c54
+ bl_0_54 br_0_54 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c54
+ bl_0_54 br_0_54 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c54
+ bl_0_54 br_0_54 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c54
+ bl_0_54 br_0_54 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c55
+ bl_0_55 br_0_55 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c55
+ bl_0_55 br_0_55 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c55
+ bl_0_55 br_0_55 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c55
+ bl_0_55 br_0_55 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c55
+ bl_0_55 br_0_55 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c55
+ bl_0_55 br_0_55 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c55
+ bl_0_55 br_0_55 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c55
+ bl_0_55 br_0_55 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c55
+ bl_0_55 br_0_55 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c55
+ bl_0_55 br_0_55 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c55
+ bl_0_55 br_0_55 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c55
+ bl_0_55 br_0_55 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c55
+ bl_0_55 br_0_55 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c55
+ bl_0_55 br_0_55 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c55
+ bl_0_55 br_0_55 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c55
+ bl_0_55 br_0_55 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c55
+ bl_0_55 br_0_55 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c55
+ bl_0_55 br_0_55 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c55
+ bl_0_55 br_0_55 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c55
+ bl_0_55 br_0_55 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c55
+ bl_0_55 br_0_55 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c55
+ bl_0_55 br_0_55 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c55
+ bl_0_55 br_0_55 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c55
+ bl_0_55 br_0_55 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c55
+ bl_0_55 br_0_55 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c55
+ bl_0_55 br_0_55 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c55
+ bl_0_55 br_0_55 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c55
+ bl_0_55 br_0_55 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c55
+ bl_0_55 br_0_55 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c55
+ bl_0_55 br_0_55 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c55
+ bl_0_55 br_0_55 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c55
+ bl_0_55 br_0_55 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c55
+ bl_0_55 br_0_55 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c55
+ bl_0_55 br_0_55 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c55
+ bl_0_55 br_0_55 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c55
+ bl_0_55 br_0_55 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c55
+ bl_0_55 br_0_55 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c55
+ bl_0_55 br_0_55 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c55
+ bl_0_55 br_0_55 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c55
+ bl_0_55 br_0_55 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c55
+ bl_0_55 br_0_55 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c55
+ bl_0_55 br_0_55 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c55
+ bl_0_55 br_0_55 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c55
+ bl_0_55 br_0_55 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c56
+ bl_0_56 br_0_56 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c56
+ bl_0_56 br_0_56 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c56
+ bl_0_56 br_0_56 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c56
+ bl_0_56 br_0_56 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c56
+ bl_0_56 br_0_56 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c56
+ bl_0_56 br_0_56 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c56
+ bl_0_56 br_0_56 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c56
+ bl_0_56 br_0_56 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c56
+ bl_0_56 br_0_56 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c56
+ bl_0_56 br_0_56 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c56
+ bl_0_56 br_0_56 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c56
+ bl_0_56 br_0_56 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c56
+ bl_0_56 br_0_56 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c56
+ bl_0_56 br_0_56 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c56
+ bl_0_56 br_0_56 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c56
+ bl_0_56 br_0_56 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c56
+ bl_0_56 br_0_56 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c56
+ bl_0_56 br_0_56 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c56
+ bl_0_56 br_0_56 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c56
+ bl_0_56 br_0_56 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c56
+ bl_0_56 br_0_56 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c56
+ bl_0_56 br_0_56 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c56
+ bl_0_56 br_0_56 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c56
+ bl_0_56 br_0_56 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c56
+ bl_0_56 br_0_56 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c56
+ bl_0_56 br_0_56 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c56
+ bl_0_56 br_0_56 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c56
+ bl_0_56 br_0_56 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c56
+ bl_0_56 br_0_56 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c56
+ bl_0_56 br_0_56 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c56
+ bl_0_56 br_0_56 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c56
+ bl_0_56 br_0_56 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c56
+ bl_0_56 br_0_56 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c56
+ bl_0_56 br_0_56 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c56
+ bl_0_56 br_0_56 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c56
+ bl_0_56 br_0_56 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c56
+ bl_0_56 br_0_56 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c56
+ bl_0_56 br_0_56 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c56
+ bl_0_56 br_0_56 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c56
+ bl_0_56 br_0_56 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c56
+ bl_0_56 br_0_56 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c56
+ bl_0_56 br_0_56 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c56
+ bl_0_56 br_0_56 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c56
+ bl_0_56 br_0_56 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c57
+ bl_0_57 br_0_57 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c57
+ bl_0_57 br_0_57 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c57
+ bl_0_57 br_0_57 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c57
+ bl_0_57 br_0_57 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c57
+ bl_0_57 br_0_57 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c57
+ bl_0_57 br_0_57 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c57
+ bl_0_57 br_0_57 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c57
+ bl_0_57 br_0_57 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c57
+ bl_0_57 br_0_57 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c57
+ bl_0_57 br_0_57 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c57
+ bl_0_57 br_0_57 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c57
+ bl_0_57 br_0_57 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c57
+ bl_0_57 br_0_57 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c57
+ bl_0_57 br_0_57 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c57
+ bl_0_57 br_0_57 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c57
+ bl_0_57 br_0_57 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c57
+ bl_0_57 br_0_57 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c57
+ bl_0_57 br_0_57 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c57
+ bl_0_57 br_0_57 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c57
+ bl_0_57 br_0_57 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c57
+ bl_0_57 br_0_57 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c57
+ bl_0_57 br_0_57 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c57
+ bl_0_57 br_0_57 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c57
+ bl_0_57 br_0_57 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c57
+ bl_0_57 br_0_57 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c57
+ bl_0_57 br_0_57 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c57
+ bl_0_57 br_0_57 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c57
+ bl_0_57 br_0_57 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c57
+ bl_0_57 br_0_57 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c57
+ bl_0_57 br_0_57 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c57
+ bl_0_57 br_0_57 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c57
+ bl_0_57 br_0_57 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c57
+ bl_0_57 br_0_57 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c57
+ bl_0_57 br_0_57 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c57
+ bl_0_57 br_0_57 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c57
+ bl_0_57 br_0_57 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c57
+ bl_0_57 br_0_57 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c57
+ bl_0_57 br_0_57 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c57
+ bl_0_57 br_0_57 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c57
+ bl_0_57 br_0_57 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c57
+ bl_0_57 br_0_57 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c57
+ bl_0_57 br_0_57 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c57
+ bl_0_57 br_0_57 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c57
+ bl_0_57 br_0_57 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c58
+ bl_0_58 br_0_58 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c58
+ bl_0_58 br_0_58 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c58
+ bl_0_58 br_0_58 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c58
+ bl_0_58 br_0_58 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c58
+ bl_0_58 br_0_58 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c58
+ bl_0_58 br_0_58 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c58
+ bl_0_58 br_0_58 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c58
+ bl_0_58 br_0_58 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c58
+ bl_0_58 br_0_58 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c58
+ bl_0_58 br_0_58 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c58
+ bl_0_58 br_0_58 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c58
+ bl_0_58 br_0_58 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c58
+ bl_0_58 br_0_58 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c58
+ bl_0_58 br_0_58 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c58
+ bl_0_58 br_0_58 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c58
+ bl_0_58 br_0_58 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c58
+ bl_0_58 br_0_58 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c58
+ bl_0_58 br_0_58 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c58
+ bl_0_58 br_0_58 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c58
+ bl_0_58 br_0_58 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c58
+ bl_0_58 br_0_58 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c58
+ bl_0_58 br_0_58 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c58
+ bl_0_58 br_0_58 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c58
+ bl_0_58 br_0_58 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c58
+ bl_0_58 br_0_58 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c58
+ bl_0_58 br_0_58 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c58
+ bl_0_58 br_0_58 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c58
+ bl_0_58 br_0_58 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c58
+ bl_0_58 br_0_58 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c58
+ bl_0_58 br_0_58 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c58
+ bl_0_58 br_0_58 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c58
+ bl_0_58 br_0_58 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c58
+ bl_0_58 br_0_58 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c58
+ bl_0_58 br_0_58 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c58
+ bl_0_58 br_0_58 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c58
+ bl_0_58 br_0_58 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c58
+ bl_0_58 br_0_58 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c58
+ bl_0_58 br_0_58 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c58
+ bl_0_58 br_0_58 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c58
+ bl_0_58 br_0_58 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c58
+ bl_0_58 br_0_58 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c58
+ bl_0_58 br_0_58 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c58
+ bl_0_58 br_0_58 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c58
+ bl_0_58 br_0_58 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c59
+ bl_0_59 br_0_59 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c59
+ bl_0_59 br_0_59 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c59
+ bl_0_59 br_0_59 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c59
+ bl_0_59 br_0_59 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c59
+ bl_0_59 br_0_59 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c59
+ bl_0_59 br_0_59 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c59
+ bl_0_59 br_0_59 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c59
+ bl_0_59 br_0_59 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c59
+ bl_0_59 br_0_59 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c59
+ bl_0_59 br_0_59 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c59
+ bl_0_59 br_0_59 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c59
+ bl_0_59 br_0_59 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c59
+ bl_0_59 br_0_59 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c59
+ bl_0_59 br_0_59 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c59
+ bl_0_59 br_0_59 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c59
+ bl_0_59 br_0_59 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c59
+ bl_0_59 br_0_59 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c59
+ bl_0_59 br_0_59 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c59
+ bl_0_59 br_0_59 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c59
+ bl_0_59 br_0_59 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c59
+ bl_0_59 br_0_59 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c59
+ bl_0_59 br_0_59 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c59
+ bl_0_59 br_0_59 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c59
+ bl_0_59 br_0_59 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c59
+ bl_0_59 br_0_59 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c59
+ bl_0_59 br_0_59 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c59
+ bl_0_59 br_0_59 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c59
+ bl_0_59 br_0_59 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c59
+ bl_0_59 br_0_59 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c59
+ bl_0_59 br_0_59 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c59
+ bl_0_59 br_0_59 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c59
+ bl_0_59 br_0_59 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c59
+ bl_0_59 br_0_59 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c59
+ bl_0_59 br_0_59 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c59
+ bl_0_59 br_0_59 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c59
+ bl_0_59 br_0_59 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c59
+ bl_0_59 br_0_59 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c59
+ bl_0_59 br_0_59 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c59
+ bl_0_59 br_0_59 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c59
+ bl_0_59 br_0_59 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c59
+ bl_0_59 br_0_59 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c59
+ bl_0_59 br_0_59 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c59
+ bl_0_59 br_0_59 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c59
+ bl_0_59 br_0_59 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c60
+ bl_0_60 br_0_60 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c60
+ bl_0_60 br_0_60 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c60
+ bl_0_60 br_0_60 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c60
+ bl_0_60 br_0_60 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c60
+ bl_0_60 br_0_60 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c60
+ bl_0_60 br_0_60 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c60
+ bl_0_60 br_0_60 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c60
+ bl_0_60 br_0_60 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c60
+ bl_0_60 br_0_60 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c60
+ bl_0_60 br_0_60 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c60
+ bl_0_60 br_0_60 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c60
+ bl_0_60 br_0_60 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c60
+ bl_0_60 br_0_60 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c60
+ bl_0_60 br_0_60 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c60
+ bl_0_60 br_0_60 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c60
+ bl_0_60 br_0_60 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c60
+ bl_0_60 br_0_60 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c60
+ bl_0_60 br_0_60 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c60
+ bl_0_60 br_0_60 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c60
+ bl_0_60 br_0_60 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c60
+ bl_0_60 br_0_60 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c60
+ bl_0_60 br_0_60 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c60
+ bl_0_60 br_0_60 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c60
+ bl_0_60 br_0_60 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c60
+ bl_0_60 br_0_60 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c60
+ bl_0_60 br_0_60 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c60
+ bl_0_60 br_0_60 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c60
+ bl_0_60 br_0_60 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c60
+ bl_0_60 br_0_60 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c60
+ bl_0_60 br_0_60 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c60
+ bl_0_60 br_0_60 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c60
+ bl_0_60 br_0_60 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c60
+ bl_0_60 br_0_60 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c60
+ bl_0_60 br_0_60 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c60
+ bl_0_60 br_0_60 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c60
+ bl_0_60 br_0_60 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c60
+ bl_0_60 br_0_60 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c60
+ bl_0_60 br_0_60 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c60
+ bl_0_60 br_0_60 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c60
+ bl_0_60 br_0_60 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c60
+ bl_0_60 br_0_60 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c60
+ bl_0_60 br_0_60 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c60
+ bl_0_60 br_0_60 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c60
+ bl_0_60 br_0_60 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c61
+ bl_0_61 br_0_61 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c61
+ bl_0_61 br_0_61 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c61
+ bl_0_61 br_0_61 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c61
+ bl_0_61 br_0_61 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c61
+ bl_0_61 br_0_61 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c61
+ bl_0_61 br_0_61 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c61
+ bl_0_61 br_0_61 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c61
+ bl_0_61 br_0_61 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c61
+ bl_0_61 br_0_61 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c61
+ bl_0_61 br_0_61 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c61
+ bl_0_61 br_0_61 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c61
+ bl_0_61 br_0_61 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c61
+ bl_0_61 br_0_61 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c61
+ bl_0_61 br_0_61 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c61
+ bl_0_61 br_0_61 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c61
+ bl_0_61 br_0_61 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c61
+ bl_0_61 br_0_61 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c61
+ bl_0_61 br_0_61 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c61
+ bl_0_61 br_0_61 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c61
+ bl_0_61 br_0_61 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c61
+ bl_0_61 br_0_61 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c61
+ bl_0_61 br_0_61 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c61
+ bl_0_61 br_0_61 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c61
+ bl_0_61 br_0_61 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c61
+ bl_0_61 br_0_61 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c61
+ bl_0_61 br_0_61 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c61
+ bl_0_61 br_0_61 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c61
+ bl_0_61 br_0_61 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c61
+ bl_0_61 br_0_61 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c61
+ bl_0_61 br_0_61 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c61
+ bl_0_61 br_0_61 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c61
+ bl_0_61 br_0_61 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c61
+ bl_0_61 br_0_61 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c61
+ bl_0_61 br_0_61 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c61
+ bl_0_61 br_0_61 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c61
+ bl_0_61 br_0_61 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c61
+ bl_0_61 br_0_61 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c61
+ bl_0_61 br_0_61 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c61
+ bl_0_61 br_0_61 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c61
+ bl_0_61 br_0_61 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c61
+ bl_0_61 br_0_61 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c61
+ bl_0_61 br_0_61 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c61
+ bl_0_61 br_0_61 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c61
+ bl_0_61 br_0_61 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c62
+ bl_0_62 br_0_62 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c62
+ bl_0_62 br_0_62 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c62
+ bl_0_62 br_0_62 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c62
+ bl_0_62 br_0_62 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c62
+ bl_0_62 br_0_62 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c62
+ bl_0_62 br_0_62 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c62
+ bl_0_62 br_0_62 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c62
+ bl_0_62 br_0_62 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c62
+ bl_0_62 br_0_62 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c62
+ bl_0_62 br_0_62 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c62
+ bl_0_62 br_0_62 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c62
+ bl_0_62 br_0_62 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c62
+ bl_0_62 br_0_62 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c62
+ bl_0_62 br_0_62 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c62
+ bl_0_62 br_0_62 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c62
+ bl_0_62 br_0_62 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c62
+ bl_0_62 br_0_62 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c62
+ bl_0_62 br_0_62 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c62
+ bl_0_62 br_0_62 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c62
+ bl_0_62 br_0_62 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c62
+ bl_0_62 br_0_62 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c62
+ bl_0_62 br_0_62 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c62
+ bl_0_62 br_0_62 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c62
+ bl_0_62 br_0_62 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c62
+ bl_0_62 br_0_62 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c62
+ bl_0_62 br_0_62 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c62
+ bl_0_62 br_0_62 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c62
+ bl_0_62 br_0_62 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c62
+ bl_0_62 br_0_62 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c62
+ bl_0_62 br_0_62 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c62
+ bl_0_62 br_0_62 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c62
+ bl_0_62 br_0_62 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c62
+ bl_0_62 br_0_62 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c62
+ bl_0_62 br_0_62 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c62
+ bl_0_62 br_0_62 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c62
+ bl_0_62 br_0_62 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c62
+ bl_0_62 br_0_62 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c62
+ bl_0_62 br_0_62 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c62
+ bl_0_62 br_0_62 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c62
+ bl_0_62 br_0_62 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c62
+ bl_0_62 br_0_62 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c62
+ bl_0_62 br_0_62 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c62
+ bl_0_62 br_0_62 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c62
+ bl_0_62 br_0_62 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c63
+ bl_0_63 br_0_63 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c63
+ bl_0_63 br_0_63 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c63
+ bl_0_63 br_0_63 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c63
+ bl_0_63 br_0_63 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c63
+ bl_0_63 br_0_63 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c63
+ bl_0_63 br_0_63 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c63
+ bl_0_63 br_0_63 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c63
+ bl_0_63 br_0_63 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c63
+ bl_0_63 br_0_63 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c63
+ bl_0_63 br_0_63 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c63
+ bl_0_63 br_0_63 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c63
+ bl_0_63 br_0_63 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c63
+ bl_0_63 br_0_63 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c63
+ bl_0_63 br_0_63 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c63
+ bl_0_63 br_0_63 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c63
+ bl_0_63 br_0_63 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c63
+ bl_0_63 br_0_63 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c63
+ bl_0_63 br_0_63 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c63
+ bl_0_63 br_0_63 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c63
+ bl_0_63 br_0_63 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c63
+ bl_0_63 br_0_63 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c63
+ bl_0_63 br_0_63 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c63
+ bl_0_63 br_0_63 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c63
+ bl_0_63 br_0_63 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c63
+ bl_0_63 br_0_63 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c63
+ bl_0_63 br_0_63 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c63
+ bl_0_63 br_0_63 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c63
+ bl_0_63 br_0_63 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c63
+ bl_0_63 br_0_63 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c63
+ bl_0_63 br_0_63 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c63
+ bl_0_63 br_0_63 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c63
+ bl_0_63 br_0_63 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c63
+ bl_0_63 br_0_63 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c63
+ bl_0_63 br_0_63 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c63
+ bl_0_63 br_0_63 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c63
+ bl_0_63 br_0_63 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c63
+ bl_0_63 br_0_63 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c63
+ bl_0_63 br_0_63 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c63
+ bl_0_63 br_0_63 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c63
+ bl_0_63 br_0_63 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c63
+ bl_0_63 br_0_63 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c63
+ bl_0_63 br_0_63 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c63
+ bl_0_63 br_0_63 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c63
+ bl_0_63 br_0_63 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c64
+ bl_0_64 br_0_64 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c64
+ bl_0_64 br_0_64 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c64
+ bl_0_64 br_0_64 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c64
+ bl_0_64 br_0_64 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c64
+ bl_0_64 br_0_64 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c64
+ bl_0_64 br_0_64 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c64
+ bl_0_64 br_0_64 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c64
+ bl_0_64 br_0_64 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c64
+ bl_0_64 br_0_64 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c64
+ bl_0_64 br_0_64 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c64
+ bl_0_64 br_0_64 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c64
+ bl_0_64 br_0_64 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c64
+ bl_0_64 br_0_64 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c64
+ bl_0_64 br_0_64 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c64
+ bl_0_64 br_0_64 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c64
+ bl_0_64 br_0_64 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c64
+ bl_0_64 br_0_64 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c64
+ bl_0_64 br_0_64 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c64
+ bl_0_64 br_0_64 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c64
+ bl_0_64 br_0_64 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c64
+ bl_0_64 br_0_64 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c64
+ bl_0_64 br_0_64 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c64
+ bl_0_64 br_0_64 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c64
+ bl_0_64 br_0_64 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c64
+ bl_0_64 br_0_64 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c64
+ bl_0_64 br_0_64 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c64
+ bl_0_64 br_0_64 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c64
+ bl_0_64 br_0_64 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c64
+ bl_0_64 br_0_64 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c64
+ bl_0_64 br_0_64 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c64
+ bl_0_64 br_0_64 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c64
+ bl_0_64 br_0_64 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c64
+ bl_0_64 br_0_64 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c64
+ bl_0_64 br_0_64 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c64
+ bl_0_64 br_0_64 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c64
+ bl_0_64 br_0_64 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c64
+ bl_0_64 br_0_64 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c64
+ bl_0_64 br_0_64 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c64
+ bl_0_64 br_0_64 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c64
+ bl_0_64 br_0_64 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c64
+ bl_0_64 br_0_64 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c64
+ bl_0_64 br_0_64 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c64
+ bl_0_64 br_0_64 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c64
+ bl_0_64 br_0_64 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c65
+ bl_0_65 br_0_65 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c65
+ bl_0_65 br_0_65 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c65
+ bl_0_65 br_0_65 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c65
+ bl_0_65 br_0_65 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c65
+ bl_0_65 br_0_65 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c65
+ bl_0_65 br_0_65 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c65
+ bl_0_65 br_0_65 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c65
+ bl_0_65 br_0_65 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c65
+ bl_0_65 br_0_65 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c65
+ bl_0_65 br_0_65 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c65
+ bl_0_65 br_0_65 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c65
+ bl_0_65 br_0_65 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c65
+ bl_0_65 br_0_65 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c65
+ bl_0_65 br_0_65 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c65
+ bl_0_65 br_0_65 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c65
+ bl_0_65 br_0_65 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c65
+ bl_0_65 br_0_65 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c65
+ bl_0_65 br_0_65 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c65
+ bl_0_65 br_0_65 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c65
+ bl_0_65 br_0_65 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c65
+ bl_0_65 br_0_65 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c65
+ bl_0_65 br_0_65 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c65
+ bl_0_65 br_0_65 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c65
+ bl_0_65 br_0_65 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c65
+ bl_0_65 br_0_65 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c65
+ bl_0_65 br_0_65 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c65
+ bl_0_65 br_0_65 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c65
+ bl_0_65 br_0_65 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c65
+ bl_0_65 br_0_65 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c65
+ bl_0_65 br_0_65 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c65
+ bl_0_65 br_0_65 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c65
+ bl_0_65 br_0_65 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c65
+ bl_0_65 br_0_65 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c65
+ bl_0_65 br_0_65 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c65
+ bl_0_65 br_0_65 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c65
+ bl_0_65 br_0_65 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c65
+ bl_0_65 br_0_65 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c65
+ bl_0_65 br_0_65 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c65
+ bl_0_65 br_0_65 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c65
+ bl_0_65 br_0_65 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c65
+ bl_0_65 br_0_65 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c65
+ bl_0_65 br_0_65 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c65
+ bl_0_65 br_0_65 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c65
+ bl_0_65 br_0_65 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c66
+ bl_0_66 br_0_66 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c66
+ bl_0_66 br_0_66 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c66
+ bl_0_66 br_0_66 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c66
+ bl_0_66 br_0_66 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c66
+ bl_0_66 br_0_66 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c66
+ bl_0_66 br_0_66 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c66
+ bl_0_66 br_0_66 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c66
+ bl_0_66 br_0_66 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c66
+ bl_0_66 br_0_66 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c66
+ bl_0_66 br_0_66 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c66
+ bl_0_66 br_0_66 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c66
+ bl_0_66 br_0_66 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c66
+ bl_0_66 br_0_66 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c66
+ bl_0_66 br_0_66 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c66
+ bl_0_66 br_0_66 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c66
+ bl_0_66 br_0_66 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c66
+ bl_0_66 br_0_66 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c66
+ bl_0_66 br_0_66 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c66
+ bl_0_66 br_0_66 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c66
+ bl_0_66 br_0_66 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c66
+ bl_0_66 br_0_66 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c66
+ bl_0_66 br_0_66 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c66
+ bl_0_66 br_0_66 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c66
+ bl_0_66 br_0_66 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c66
+ bl_0_66 br_0_66 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c66
+ bl_0_66 br_0_66 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c66
+ bl_0_66 br_0_66 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c66
+ bl_0_66 br_0_66 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c66
+ bl_0_66 br_0_66 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c66
+ bl_0_66 br_0_66 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c66
+ bl_0_66 br_0_66 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c66
+ bl_0_66 br_0_66 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c66
+ bl_0_66 br_0_66 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c66
+ bl_0_66 br_0_66 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c66
+ bl_0_66 br_0_66 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c66
+ bl_0_66 br_0_66 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c66
+ bl_0_66 br_0_66 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c66
+ bl_0_66 br_0_66 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c66
+ bl_0_66 br_0_66 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c66
+ bl_0_66 br_0_66 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c66
+ bl_0_66 br_0_66 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c66
+ bl_0_66 br_0_66 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c66
+ bl_0_66 br_0_66 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c66
+ bl_0_66 br_0_66 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c67
+ bl_0_67 br_0_67 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c67
+ bl_0_67 br_0_67 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c67
+ bl_0_67 br_0_67 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c67
+ bl_0_67 br_0_67 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c67
+ bl_0_67 br_0_67 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c67
+ bl_0_67 br_0_67 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c67
+ bl_0_67 br_0_67 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c67
+ bl_0_67 br_0_67 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c67
+ bl_0_67 br_0_67 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c67
+ bl_0_67 br_0_67 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c67
+ bl_0_67 br_0_67 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c67
+ bl_0_67 br_0_67 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c67
+ bl_0_67 br_0_67 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c67
+ bl_0_67 br_0_67 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c67
+ bl_0_67 br_0_67 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c67
+ bl_0_67 br_0_67 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c67
+ bl_0_67 br_0_67 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c67
+ bl_0_67 br_0_67 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c67
+ bl_0_67 br_0_67 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c67
+ bl_0_67 br_0_67 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c67
+ bl_0_67 br_0_67 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c67
+ bl_0_67 br_0_67 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c67
+ bl_0_67 br_0_67 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c67
+ bl_0_67 br_0_67 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c67
+ bl_0_67 br_0_67 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c67
+ bl_0_67 br_0_67 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c67
+ bl_0_67 br_0_67 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c67
+ bl_0_67 br_0_67 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c67
+ bl_0_67 br_0_67 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c67
+ bl_0_67 br_0_67 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c67
+ bl_0_67 br_0_67 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c67
+ bl_0_67 br_0_67 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c67
+ bl_0_67 br_0_67 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c67
+ bl_0_67 br_0_67 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c67
+ bl_0_67 br_0_67 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c67
+ bl_0_67 br_0_67 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c67
+ bl_0_67 br_0_67 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c67
+ bl_0_67 br_0_67 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c67
+ bl_0_67 br_0_67 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c67
+ bl_0_67 br_0_67 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c67
+ bl_0_67 br_0_67 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c67
+ bl_0_67 br_0_67 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c67
+ bl_0_67 br_0_67 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c67
+ bl_0_67 br_0_67 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c68
+ bl_0_68 br_0_68 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c68
+ bl_0_68 br_0_68 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c68
+ bl_0_68 br_0_68 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c68
+ bl_0_68 br_0_68 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c68
+ bl_0_68 br_0_68 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c68
+ bl_0_68 br_0_68 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c68
+ bl_0_68 br_0_68 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c68
+ bl_0_68 br_0_68 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c68
+ bl_0_68 br_0_68 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c68
+ bl_0_68 br_0_68 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c68
+ bl_0_68 br_0_68 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c68
+ bl_0_68 br_0_68 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c68
+ bl_0_68 br_0_68 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c68
+ bl_0_68 br_0_68 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c68
+ bl_0_68 br_0_68 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c68
+ bl_0_68 br_0_68 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c68
+ bl_0_68 br_0_68 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c68
+ bl_0_68 br_0_68 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c68
+ bl_0_68 br_0_68 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c68
+ bl_0_68 br_0_68 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c68
+ bl_0_68 br_0_68 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c68
+ bl_0_68 br_0_68 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c68
+ bl_0_68 br_0_68 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c68
+ bl_0_68 br_0_68 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c68
+ bl_0_68 br_0_68 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c68
+ bl_0_68 br_0_68 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c68
+ bl_0_68 br_0_68 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c68
+ bl_0_68 br_0_68 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c68
+ bl_0_68 br_0_68 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c68
+ bl_0_68 br_0_68 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c68
+ bl_0_68 br_0_68 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c68
+ bl_0_68 br_0_68 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c68
+ bl_0_68 br_0_68 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c68
+ bl_0_68 br_0_68 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c68
+ bl_0_68 br_0_68 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c68
+ bl_0_68 br_0_68 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c68
+ bl_0_68 br_0_68 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c68
+ bl_0_68 br_0_68 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c68
+ bl_0_68 br_0_68 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c68
+ bl_0_68 br_0_68 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c68
+ bl_0_68 br_0_68 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c68
+ bl_0_68 br_0_68 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c68
+ bl_0_68 br_0_68 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c68
+ bl_0_68 br_0_68 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c69
+ bl_0_69 br_0_69 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c69
+ bl_0_69 br_0_69 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c69
+ bl_0_69 br_0_69 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c69
+ bl_0_69 br_0_69 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c69
+ bl_0_69 br_0_69 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c69
+ bl_0_69 br_0_69 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c69
+ bl_0_69 br_0_69 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c69
+ bl_0_69 br_0_69 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c69
+ bl_0_69 br_0_69 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c69
+ bl_0_69 br_0_69 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c69
+ bl_0_69 br_0_69 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c69
+ bl_0_69 br_0_69 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c69
+ bl_0_69 br_0_69 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c69
+ bl_0_69 br_0_69 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c69
+ bl_0_69 br_0_69 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c69
+ bl_0_69 br_0_69 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c69
+ bl_0_69 br_0_69 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c69
+ bl_0_69 br_0_69 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c69
+ bl_0_69 br_0_69 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c69
+ bl_0_69 br_0_69 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c69
+ bl_0_69 br_0_69 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c69
+ bl_0_69 br_0_69 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c69
+ bl_0_69 br_0_69 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c69
+ bl_0_69 br_0_69 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c69
+ bl_0_69 br_0_69 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c69
+ bl_0_69 br_0_69 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c69
+ bl_0_69 br_0_69 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c69
+ bl_0_69 br_0_69 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c69
+ bl_0_69 br_0_69 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c69
+ bl_0_69 br_0_69 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c69
+ bl_0_69 br_0_69 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c69
+ bl_0_69 br_0_69 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c69
+ bl_0_69 br_0_69 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c69
+ bl_0_69 br_0_69 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c69
+ bl_0_69 br_0_69 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c69
+ bl_0_69 br_0_69 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c69
+ bl_0_69 br_0_69 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c69
+ bl_0_69 br_0_69 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c69
+ bl_0_69 br_0_69 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c69
+ bl_0_69 br_0_69 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c69
+ bl_0_69 br_0_69 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c69
+ bl_0_69 br_0_69 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c69
+ bl_0_69 br_0_69 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c69
+ bl_0_69 br_0_69 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c70
+ bl_0_70 br_0_70 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c70
+ bl_0_70 br_0_70 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c70
+ bl_0_70 br_0_70 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c70
+ bl_0_70 br_0_70 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c70
+ bl_0_70 br_0_70 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c70
+ bl_0_70 br_0_70 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c70
+ bl_0_70 br_0_70 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c70
+ bl_0_70 br_0_70 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c70
+ bl_0_70 br_0_70 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c70
+ bl_0_70 br_0_70 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c70
+ bl_0_70 br_0_70 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c70
+ bl_0_70 br_0_70 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c70
+ bl_0_70 br_0_70 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c70
+ bl_0_70 br_0_70 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c70
+ bl_0_70 br_0_70 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c70
+ bl_0_70 br_0_70 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c70
+ bl_0_70 br_0_70 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c70
+ bl_0_70 br_0_70 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c70
+ bl_0_70 br_0_70 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c70
+ bl_0_70 br_0_70 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c70
+ bl_0_70 br_0_70 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c70
+ bl_0_70 br_0_70 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c70
+ bl_0_70 br_0_70 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c70
+ bl_0_70 br_0_70 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c70
+ bl_0_70 br_0_70 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c70
+ bl_0_70 br_0_70 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c70
+ bl_0_70 br_0_70 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c70
+ bl_0_70 br_0_70 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c70
+ bl_0_70 br_0_70 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c70
+ bl_0_70 br_0_70 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c70
+ bl_0_70 br_0_70 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c70
+ bl_0_70 br_0_70 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c70
+ bl_0_70 br_0_70 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c70
+ bl_0_70 br_0_70 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c70
+ bl_0_70 br_0_70 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c70
+ bl_0_70 br_0_70 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c70
+ bl_0_70 br_0_70 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c70
+ bl_0_70 br_0_70 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c70
+ bl_0_70 br_0_70 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c70
+ bl_0_70 br_0_70 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c70
+ bl_0_70 br_0_70 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c70
+ bl_0_70 br_0_70 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c70
+ bl_0_70 br_0_70 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c70
+ bl_0_70 br_0_70 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c71
+ bl_0_71 br_0_71 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c71
+ bl_0_71 br_0_71 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c71
+ bl_0_71 br_0_71 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c71
+ bl_0_71 br_0_71 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c71
+ bl_0_71 br_0_71 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c71
+ bl_0_71 br_0_71 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c71
+ bl_0_71 br_0_71 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c71
+ bl_0_71 br_0_71 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c71
+ bl_0_71 br_0_71 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c71
+ bl_0_71 br_0_71 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c71
+ bl_0_71 br_0_71 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c71
+ bl_0_71 br_0_71 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c71
+ bl_0_71 br_0_71 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c71
+ bl_0_71 br_0_71 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c71
+ bl_0_71 br_0_71 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c71
+ bl_0_71 br_0_71 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c71
+ bl_0_71 br_0_71 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c71
+ bl_0_71 br_0_71 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c71
+ bl_0_71 br_0_71 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c71
+ bl_0_71 br_0_71 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c71
+ bl_0_71 br_0_71 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c71
+ bl_0_71 br_0_71 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c71
+ bl_0_71 br_0_71 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c71
+ bl_0_71 br_0_71 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c71
+ bl_0_71 br_0_71 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c71
+ bl_0_71 br_0_71 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c71
+ bl_0_71 br_0_71 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c71
+ bl_0_71 br_0_71 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c71
+ bl_0_71 br_0_71 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c71
+ bl_0_71 br_0_71 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c71
+ bl_0_71 br_0_71 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c71
+ bl_0_71 br_0_71 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c71
+ bl_0_71 br_0_71 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c71
+ bl_0_71 br_0_71 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c71
+ bl_0_71 br_0_71 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c71
+ bl_0_71 br_0_71 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c71
+ bl_0_71 br_0_71 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c71
+ bl_0_71 br_0_71 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c71
+ bl_0_71 br_0_71 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c71
+ bl_0_71 br_0_71 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c71
+ bl_0_71 br_0_71 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c71
+ bl_0_71 br_0_71 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c71
+ bl_0_71 br_0_71 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c71
+ bl_0_71 br_0_71 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c72
+ bl_0_72 br_0_72 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c72
+ bl_0_72 br_0_72 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c72
+ bl_0_72 br_0_72 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c72
+ bl_0_72 br_0_72 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c72
+ bl_0_72 br_0_72 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c72
+ bl_0_72 br_0_72 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c72
+ bl_0_72 br_0_72 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c72
+ bl_0_72 br_0_72 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c72
+ bl_0_72 br_0_72 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c72
+ bl_0_72 br_0_72 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c72
+ bl_0_72 br_0_72 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c72
+ bl_0_72 br_0_72 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c72
+ bl_0_72 br_0_72 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c72
+ bl_0_72 br_0_72 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c72
+ bl_0_72 br_0_72 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c72
+ bl_0_72 br_0_72 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c72
+ bl_0_72 br_0_72 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c72
+ bl_0_72 br_0_72 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c72
+ bl_0_72 br_0_72 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c72
+ bl_0_72 br_0_72 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c72
+ bl_0_72 br_0_72 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c72
+ bl_0_72 br_0_72 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c72
+ bl_0_72 br_0_72 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c72
+ bl_0_72 br_0_72 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c72
+ bl_0_72 br_0_72 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c72
+ bl_0_72 br_0_72 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c72
+ bl_0_72 br_0_72 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c72
+ bl_0_72 br_0_72 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c72
+ bl_0_72 br_0_72 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c72
+ bl_0_72 br_0_72 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c72
+ bl_0_72 br_0_72 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c72
+ bl_0_72 br_0_72 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c72
+ bl_0_72 br_0_72 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c72
+ bl_0_72 br_0_72 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c72
+ bl_0_72 br_0_72 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c72
+ bl_0_72 br_0_72 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c72
+ bl_0_72 br_0_72 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c72
+ bl_0_72 br_0_72 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c72
+ bl_0_72 br_0_72 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c72
+ bl_0_72 br_0_72 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c72
+ bl_0_72 br_0_72 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c72
+ bl_0_72 br_0_72 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c72
+ bl_0_72 br_0_72 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c72
+ bl_0_72 br_0_72 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c73
+ bl_0_73 br_0_73 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c73
+ bl_0_73 br_0_73 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c73
+ bl_0_73 br_0_73 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c73
+ bl_0_73 br_0_73 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c73
+ bl_0_73 br_0_73 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c73
+ bl_0_73 br_0_73 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c73
+ bl_0_73 br_0_73 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c73
+ bl_0_73 br_0_73 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c73
+ bl_0_73 br_0_73 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c73
+ bl_0_73 br_0_73 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c73
+ bl_0_73 br_0_73 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c73
+ bl_0_73 br_0_73 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c73
+ bl_0_73 br_0_73 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c73
+ bl_0_73 br_0_73 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c73
+ bl_0_73 br_0_73 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c73
+ bl_0_73 br_0_73 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c73
+ bl_0_73 br_0_73 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c73
+ bl_0_73 br_0_73 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c73
+ bl_0_73 br_0_73 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c73
+ bl_0_73 br_0_73 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c73
+ bl_0_73 br_0_73 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c73
+ bl_0_73 br_0_73 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c73
+ bl_0_73 br_0_73 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c73
+ bl_0_73 br_0_73 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c73
+ bl_0_73 br_0_73 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c73
+ bl_0_73 br_0_73 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c73
+ bl_0_73 br_0_73 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c73
+ bl_0_73 br_0_73 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c73
+ bl_0_73 br_0_73 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c73
+ bl_0_73 br_0_73 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c73
+ bl_0_73 br_0_73 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c73
+ bl_0_73 br_0_73 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c73
+ bl_0_73 br_0_73 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c73
+ bl_0_73 br_0_73 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c73
+ bl_0_73 br_0_73 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c73
+ bl_0_73 br_0_73 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c73
+ bl_0_73 br_0_73 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c73
+ bl_0_73 br_0_73 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c73
+ bl_0_73 br_0_73 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c73
+ bl_0_73 br_0_73 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c73
+ bl_0_73 br_0_73 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c73
+ bl_0_73 br_0_73 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c73
+ bl_0_73 br_0_73 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c73
+ bl_0_73 br_0_73 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c74
+ bl_0_74 br_0_74 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c74
+ bl_0_74 br_0_74 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c74
+ bl_0_74 br_0_74 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c74
+ bl_0_74 br_0_74 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c74
+ bl_0_74 br_0_74 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c74
+ bl_0_74 br_0_74 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c74
+ bl_0_74 br_0_74 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c74
+ bl_0_74 br_0_74 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c74
+ bl_0_74 br_0_74 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c74
+ bl_0_74 br_0_74 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c74
+ bl_0_74 br_0_74 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c74
+ bl_0_74 br_0_74 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c74
+ bl_0_74 br_0_74 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c74
+ bl_0_74 br_0_74 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c74
+ bl_0_74 br_0_74 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c74
+ bl_0_74 br_0_74 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c74
+ bl_0_74 br_0_74 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c74
+ bl_0_74 br_0_74 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c74
+ bl_0_74 br_0_74 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c74
+ bl_0_74 br_0_74 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c74
+ bl_0_74 br_0_74 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c74
+ bl_0_74 br_0_74 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c74
+ bl_0_74 br_0_74 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c74
+ bl_0_74 br_0_74 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c74
+ bl_0_74 br_0_74 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c74
+ bl_0_74 br_0_74 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c74
+ bl_0_74 br_0_74 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c74
+ bl_0_74 br_0_74 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c74
+ bl_0_74 br_0_74 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c74
+ bl_0_74 br_0_74 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c74
+ bl_0_74 br_0_74 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c74
+ bl_0_74 br_0_74 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c74
+ bl_0_74 br_0_74 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c74
+ bl_0_74 br_0_74 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c74
+ bl_0_74 br_0_74 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c74
+ bl_0_74 br_0_74 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c74
+ bl_0_74 br_0_74 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c74
+ bl_0_74 br_0_74 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c74
+ bl_0_74 br_0_74 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c74
+ bl_0_74 br_0_74 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c74
+ bl_0_74 br_0_74 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c74
+ bl_0_74 br_0_74 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c74
+ bl_0_74 br_0_74 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c74
+ bl_0_74 br_0_74 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c75
+ bl_0_75 br_0_75 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c75
+ bl_0_75 br_0_75 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c75
+ bl_0_75 br_0_75 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c75
+ bl_0_75 br_0_75 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c75
+ bl_0_75 br_0_75 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c75
+ bl_0_75 br_0_75 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c75
+ bl_0_75 br_0_75 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c75
+ bl_0_75 br_0_75 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c75
+ bl_0_75 br_0_75 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c75
+ bl_0_75 br_0_75 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c75
+ bl_0_75 br_0_75 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c75
+ bl_0_75 br_0_75 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c75
+ bl_0_75 br_0_75 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c75
+ bl_0_75 br_0_75 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c75
+ bl_0_75 br_0_75 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c75
+ bl_0_75 br_0_75 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c75
+ bl_0_75 br_0_75 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c75
+ bl_0_75 br_0_75 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c75
+ bl_0_75 br_0_75 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c75
+ bl_0_75 br_0_75 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c75
+ bl_0_75 br_0_75 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c75
+ bl_0_75 br_0_75 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c75
+ bl_0_75 br_0_75 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c75
+ bl_0_75 br_0_75 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c75
+ bl_0_75 br_0_75 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c75
+ bl_0_75 br_0_75 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c75
+ bl_0_75 br_0_75 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c75
+ bl_0_75 br_0_75 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c75
+ bl_0_75 br_0_75 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c75
+ bl_0_75 br_0_75 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c75
+ bl_0_75 br_0_75 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c75
+ bl_0_75 br_0_75 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c75
+ bl_0_75 br_0_75 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c75
+ bl_0_75 br_0_75 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c75
+ bl_0_75 br_0_75 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c75
+ bl_0_75 br_0_75 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c75
+ bl_0_75 br_0_75 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c75
+ bl_0_75 br_0_75 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c75
+ bl_0_75 br_0_75 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c75
+ bl_0_75 br_0_75 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c75
+ bl_0_75 br_0_75 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c75
+ bl_0_75 br_0_75 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c75
+ bl_0_75 br_0_75 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c75
+ bl_0_75 br_0_75 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c76
+ bl_0_76 br_0_76 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c76
+ bl_0_76 br_0_76 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c76
+ bl_0_76 br_0_76 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c76
+ bl_0_76 br_0_76 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c76
+ bl_0_76 br_0_76 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c76
+ bl_0_76 br_0_76 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c76
+ bl_0_76 br_0_76 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c76
+ bl_0_76 br_0_76 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c76
+ bl_0_76 br_0_76 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c76
+ bl_0_76 br_0_76 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c76
+ bl_0_76 br_0_76 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c76
+ bl_0_76 br_0_76 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c76
+ bl_0_76 br_0_76 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c76
+ bl_0_76 br_0_76 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c76
+ bl_0_76 br_0_76 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c76
+ bl_0_76 br_0_76 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c76
+ bl_0_76 br_0_76 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c76
+ bl_0_76 br_0_76 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c76
+ bl_0_76 br_0_76 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c76
+ bl_0_76 br_0_76 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c76
+ bl_0_76 br_0_76 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c76
+ bl_0_76 br_0_76 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c76
+ bl_0_76 br_0_76 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c76
+ bl_0_76 br_0_76 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c76
+ bl_0_76 br_0_76 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c76
+ bl_0_76 br_0_76 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c76
+ bl_0_76 br_0_76 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c76
+ bl_0_76 br_0_76 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c76
+ bl_0_76 br_0_76 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c76
+ bl_0_76 br_0_76 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c76
+ bl_0_76 br_0_76 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c76
+ bl_0_76 br_0_76 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c76
+ bl_0_76 br_0_76 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c76
+ bl_0_76 br_0_76 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c76
+ bl_0_76 br_0_76 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c76
+ bl_0_76 br_0_76 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c76
+ bl_0_76 br_0_76 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c76
+ bl_0_76 br_0_76 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c76
+ bl_0_76 br_0_76 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c76
+ bl_0_76 br_0_76 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c76
+ bl_0_76 br_0_76 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c76
+ bl_0_76 br_0_76 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c76
+ bl_0_76 br_0_76 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c76
+ bl_0_76 br_0_76 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c77
+ bl_0_77 br_0_77 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c77
+ bl_0_77 br_0_77 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c77
+ bl_0_77 br_0_77 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c77
+ bl_0_77 br_0_77 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c77
+ bl_0_77 br_0_77 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c77
+ bl_0_77 br_0_77 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c77
+ bl_0_77 br_0_77 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c77
+ bl_0_77 br_0_77 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c77
+ bl_0_77 br_0_77 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c77
+ bl_0_77 br_0_77 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c77
+ bl_0_77 br_0_77 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c77
+ bl_0_77 br_0_77 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c77
+ bl_0_77 br_0_77 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c77
+ bl_0_77 br_0_77 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c77
+ bl_0_77 br_0_77 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c77
+ bl_0_77 br_0_77 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c77
+ bl_0_77 br_0_77 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c77
+ bl_0_77 br_0_77 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c77
+ bl_0_77 br_0_77 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c77
+ bl_0_77 br_0_77 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c77
+ bl_0_77 br_0_77 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c77
+ bl_0_77 br_0_77 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c77
+ bl_0_77 br_0_77 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c77
+ bl_0_77 br_0_77 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c77
+ bl_0_77 br_0_77 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c77
+ bl_0_77 br_0_77 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c77
+ bl_0_77 br_0_77 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c77
+ bl_0_77 br_0_77 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c77
+ bl_0_77 br_0_77 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c77
+ bl_0_77 br_0_77 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c77
+ bl_0_77 br_0_77 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c77
+ bl_0_77 br_0_77 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c77
+ bl_0_77 br_0_77 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c77
+ bl_0_77 br_0_77 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c77
+ bl_0_77 br_0_77 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c77
+ bl_0_77 br_0_77 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c77
+ bl_0_77 br_0_77 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c77
+ bl_0_77 br_0_77 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c77
+ bl_0_77 br_0_77 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c77
+ bl_0_77 br_0_77 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c77
+ bl_0_77 br_0_77 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c77
+ bl_0_77 br_0_77 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c77
+ bl_0_77 br_0_77 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c77
+ bl_0_77 br_0_77 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c78
+ bl_0_78 br_0_78 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c78
+ bl_0_78 br_0_78 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c78
+ bl_0_78 br_0_78 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c78
+ bl_0_78 br_0_78 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c78
+ bl_0_78 br_0_78 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c78
+ bl_0_78 br_0_78 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c78
+ bl_0_78 br_0_78 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c78
+ bl_0_78 br_0_78 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c78
+ bl_0_78 br_0_78 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c78
+ bl_0_78 br_0_78 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c78
+ bl_0_78 br_0_78 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c78
+ bl_0_78 br_0_78 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c78
+ bl_0_78 br_0_78 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c78
+ bl_0_78 br_0_78 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c78
+ bl_0_78 br_0_78 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c78
+ bl_0_78 br_0_78 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c78
+ bl_0_78 br_0_78 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c78
+ bl_0_78 br_0_78 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c78
+ bl_0_78 br_0_78 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c78
+ bl_0_78 br_0_78 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c78
+ bl_0_78 br_0_78 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c78
+ bl_0_78 br_0_78 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c78
+ bl_0_78 br_0_78 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c78
+ bl_0_78 br_0_78 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c78
+ bl_0_78 br_0_78 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c78
+ bl_0_78 br_0_78 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c78
+ bl_0_78 br_0_78 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c78
+ bl_0_78 br_0_78 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c78
+ bl_0_78 br_0_78 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c78
+ bl_0_78 br_0_78 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c78
+ bl_0_78 br_0_78 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c78
+ bl_0_78 br_0_78 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c78
+ bl_0_78 br_0_78 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c78
+ bl_0_78 br_0_78 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c78
+ bl_0_78 br_0_78 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c78
+ bl_0_78 br_0_78 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c78
+ bl_0_78 br_0_78 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c78
+ bl_0_78 br_0_78 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c78
+ bl_0_78 br_0_78 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c78
+ bl_0_78 br_0_78 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c78
+ bl_0_78 br_0_78 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c78
+ bl_0_78 br_0_78 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c78
+ bl_0_78 br_0_78 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c78
+ bl_0_78 br_0_78 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c79
+ bl_0_79 br_0_79 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c79
+ bl_0_79 br_0_79 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c79
+ bl_0_79 br_0_79 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c79
+ bl_0_79 br_0_79 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c79
+ bl_0_79 br_0_79 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c79
+ bl_0_79 br_0_79 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c79
+ bl_0_79 br_0_79 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c79
+ bl_0_79 br_0_79 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c79
+ bl_0_79 br_0_79 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c79
+ bl_0_79 br_0_79 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c79
+ bl_0_79 br_0_79 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c79
+ bl_0_79 br_0_79 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c79
+ bl_0_79 br_0_79 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c79
+ bl_0_79 br_0_79 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c79
+ bl_0_79 br_0_79 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c79
+ bl_0_79 br_0_79 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c79
+ bl_0_79 br_0_79 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c79
+ bl_0_79 br_0_79 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c79
+ bl_0_79 br_0_79 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c79
+ bl_0_79 br_0_79 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c79
+ bl_0_79 br_0_79 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c79
+ bl_0_79 br_0_79 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c79
+ bl_0_79 br_0_79 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c79
+ bl_0_79 br_0_79 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c79
+ bl_0_79 br_0_79 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c79
+ bl_0_79 br_0_79 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c79
+ bl_0_79 br_0_79 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c79
+ bl_0_79 br_0_79 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c79
+ bl_0_79 br_0_79 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c79
+ bl_0_79 br_0_79 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c79
+ bl_0_79 br_0_79 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c79
+ bl_0_79 br_0_79 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c79
+ bl_0_79 br_0_79 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c79
+ bl_0_79 br_0_79 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c79
+ bl_0_79 br_0_79 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c79
+ bl_0_79 br_0_79 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c79
+ bl_0_79 br_0_79 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c79
+ bl_0_79 br_0_79 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c79
+ bl_0_79 br_0_79 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c79
+ bl_0_79 br_0_79 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c79
+ bl_0_79 br_0_79 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c79
+ bl_0_79 br_0_79 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c79
+ bl_0_79 br_0_79 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c79
+ bl_0_79 br_0_79 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c80
+ bl_0_80 br_0_80 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c80
+ bl_0_80 br_0_80 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c80
+ bl_0_80 br_0_80 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c80
+ bl_0_80 br_0_80 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c80
+ bl_0_80 br_0_80 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c80
+ bl_0_80 br_0_80 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c80
+ bl_0_80 br_0_80 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c80
+ bl_0_80 br_0_80 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c80
+ bl_0_80 br_0_80 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c80
+ bl_0_80 br_0_80 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c80
+ bl_0_80 br_0_80 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c80
+ bl_0_80 br_0_80 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c80
+ bl_0_80 br_0_80 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c80
+ bl_0_80 br_0_80 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c80
+ bl_0_80 br_0_80 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c80
+ bl_0_80 br_0_80 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c80
+ bl_0_80 br_0_80 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c80
+ bl_0_80 br_0_80 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c80
+ bl_0_80 br_0_80 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c80
+ bl_0_80 br_0_80 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c80
+ bl_0_80 br_0_80 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c80
+ bl_0_80 br_0_80 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c80
+ bl_0_80 br_0_80 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c80
+ bl_0_80 br_0_80 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c80
+ bl_0_80 br_0_80 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c80
+ bl_0_80 br_0_80 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c80
+ bl_0_80 br_0_80 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c80
+ bl_0_80 br_0_80 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c80
+ bl_0_80 br_0_80 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c80
+ bl_0_80 br_0_80 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c80
+ bl_0_80 br_0_80 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c80
+ bl_0_80 br_0_80 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c80
+ bl_0_80 br_0_80 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c80
+ bl_0_80 br_0_80 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c80
+ bl_0_80 br_0_80 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c80
+ bl_0_80 br_0_80 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c80
+ bl_0_80 br_0_80 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c80
+ bl_0_80 br_0_80 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c80
+ bl_0_80 br_0_80 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c80
+ bl_0_80 br_0_80 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c80
+ bl_0_80 br_0_80 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c80
+ bl_0_80 br_0_80 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c80
+ bl_0_80 br_0_80 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c80
+ bl_0_80 br_0_80 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c81
+ bl_0_81 br_0_81 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c81
+ bl_0_81 br_0_81 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c81
+ bl_0_81 br_0_81 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c81
+ bl_0_81 br_0_81 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c81
+ bl_0_81 br_0_81 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c81
+ bl_0_81 br_0_81 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c81
+ bl_0_81 br_0_81 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c81
+ bl_0_81 br_0_81 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c81
+ bl_0_81 br_0_81 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c81
+ bl_0_81 br_0_81 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c81
+ bl_0_81 br_0_81 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c81
+ bl_0_81 br_0_81 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c81
+ bl_0_81 br_0_81 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c81
+ bl_0_81 br_0_81 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c81
+ bl_0_81 br_0_81 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c81
+ bl_0_81 br_0_81 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c81
+ bl_0_81 br_0_81 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c81
+ bl_0_81 br_0_81 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c81
+ bl_0_81 br_0_81 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c81
+ bl_0_81 br_0_81 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c81
+ bl_0_81 br_0_81 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c81
+ bl_0_81 br_0_81 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c81
+ bl_0_81 br_0_81 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c81
+ bl_0_81 br_0_81 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c81
+ bl_0_81 br_0_81 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c81
+ bl_0_81 br_0_81 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c81
+ bl_0_81 br_0_81 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c81
+ bl_0_81 br_0_81 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c81
+ bl_0_81 br_0_81 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c81
+ bl_0_81 br_0_81 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c81
+ bl_0_81 br_0_81 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c81
+ bl_0_81 br_0_81 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c81
+ bl_0_81 br_0_81 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c81
+ bl_0_81 br_0_81 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c81
+ bl_0_81 br_0_81 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c81
+ bl_0_81 br_0_81 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c81
+ bl_0_81 br_0_81 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c81
+ bl_0_81 br_0_81 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c81
+ bl_0_81 br_0_81 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c81
+ bl_0_81 br_0_81 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c81
+ bl_0_81 br_0_81 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c81
+ bl_0_81 br_0_81 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c81
+ bl_0_81 br_0_81 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c81
+ bl_0_81 br_0_81 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c82
+ bl_0_82 br_0_82 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c82
+ bl_0_82 br_0_82 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c82
+ bl_0_82 br_0_82 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c82
+ bl_0_82 br_0_82 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c82
+ bl_0_82 br_0_82 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c82
+ bl_0_82 br_0_82 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c82
+ bl_0_82 br_0_82 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c82
+ bl_0_82 br_0_82 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c82
+ bl_0_82 br_0_82 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c82
+ bl_0_82 br_0_82 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c82
+ bl_0_82 br_0_82 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c82
+ bl_0_82 br_0_82 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c82
+ bl_0_82 br_0_82 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c82
+ bl_0_82 br_0_82 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c82
+ bl_0_82 br_0_82 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c82
+ bl_0_82 br_0_82 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c82
+ bl_0_82 br_0_82 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c82
+ bl_0_82 br_0_82 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c82
+ bl_0_82 br_0_82 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c82
+ bl_0_82 br_0_82 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c82
+ bl_0_82 br_0_82 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c82
+ bl_0_82 br_0_82 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c82
+ bl_0_82 br_0_82 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c82
+ bl_0_82 br_0_82 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c82
+ bl_0_82 br_0_82 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c82
+ bl_0_82 br_0_82 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c82
+ bl_0_82 br_0_82 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c82
+ bl_0_82 br_0_82 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c82
+ bl_0_82 br_0_82 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c82
+ bl_0_82 br_0_82 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c82
+ bl_0_82 br_0_82 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c82
+ bl_0_82 br_0_82 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c82
+ bl_0_82 br_0_82 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c82
+ bl_0_82 br_0_82 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c82
+ bl_0_82 br_0_82 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c82
+ bl_0_82 br_0_82 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c82
+ bl_0_82 br_0_82 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c82
+ bl_0_82 br_0_82 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c82
+ bl_0_82 br_0_82 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c82
+ bl_0_82 br_0_82 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c82
+ bl_0_82 br_0_82 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c82
+ bl_0_82 br_0_82 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c82
+ bl_0_82 br_0_82 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c82
+ bl_0_82 br_0_82 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c83
+ bl_0_83 br_0_83 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c83
+ bl_0_83 br_0_83 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c83
+ bl_0_83 br_0_83 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c83
+ bl_0_83 br_0_83 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c83
+ bl_0_83 br_0_83 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c83
+ bl_0_83 br_0_83 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c83
+ bl_0_83 br_0_83 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c83
+ bl_0_83 br_0_83 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c83
+ bl_0_83 br_0_83 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c83
+ bl_0_83 br_0_83 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c83
+ bl_0_83 br_0_83 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c83
+ bl_0_83 br_0_83 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c83
+ bl_0_83 br_0_83 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c83
+ bl_0_83 br_0_83 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c83
+ bl_0_83 br_0_83 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c83
+ bl_0_83 br_0_83 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c83
+ bl_0_83 br_0_83 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c83
+ bl_0_83 br_0_83 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c83
+ bl_0_83 br_0_83 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c83
+ bl_0_83 br_0_83 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c83
+ bl_0_83 br_0_83 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c83
+ bl_0_83 br_0_83 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c83
+ bl_0_83 br_0_83 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c83
+ bl_0_83 br_0_83 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c83
+ bl_0_83 br_0_83 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c83
+ bl_0_83 br_0_83 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c83
+ bl_0_83 br_0_83 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c83
+ bl_0_83 br_0_83 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c83
+ bl_0_83 br_0_83 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c83
+ bl_0_83 br_0_83 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c83
+ bl_0_83 br_0_83 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c83
+ bl_0_83 br_0_83 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c83
+ bl_0_83 br_0_83 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c83
+ bl_0_83 br_0_83 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c83
+ bl_0_83 br_0_83 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c83
+ bl_0_83 br_0_83 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c83
+ bl_0_83 br_0_83 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c83
+ bl_0_83 br_0_83 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c83
+ bl_0_83 br_0_83 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c83
+ bl_0_83 br_0_83 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c83
+ bl_0_83 br_0_83 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c83
+ bl_0_83 br_0_83 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c83
+ bl_0_83 br_0_83 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c83
+ bl_0_83 br_0_83 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c84
+ bl_0_84 br_0_84 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c84
+ bl_0_84 br_0_84 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c84
+ bl_0_84 br_0_84 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c84
+ bl_0_84 br_0_84 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c84
+ bl_0_84 br_0_84 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c84
+ bl_0_84 br_0_84 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c84
+ bl_0_84 br_0_84 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c84
+ bl_0_84 br_0_84 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c84
+ bl_0_84 br_0_84 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c84
+ bl_0_84 br_0_84 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c84
+ bl_0_84 br_0_84 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c84
+ bl_0_84 br_0_84 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c84
+ bl_0_84 br_0_84 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c84
+ bl_0_84 br_0_84 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c84
+ bl_0_84 br_0_84 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c84
+ bl_0_84 br_0_84 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c84
+ bl_0_84 br_0_84 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c84
+ bl_0_84 br_0_84 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c84
+ bl_0_84 br_0_84 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c84
+ bl_0_84 br_0_84 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c84
+ bl_0_84 br_0_84 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c84
+ bl_0_84 br_0_84 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c84
+ bl_0_84 br_0_84 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c84
+ bl_0_84 br_0_84 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c84
+ bl_0_84 br_0_84 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c84
+ bl_0_84 br_0_84 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c84
+ bl_0_84 br_0_84 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c84
+ bl_0_84 br_0_84 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c84
+ bl_0_84 br_0_84 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c84
+ bl_0_84 br_0_84 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c84
+ bl_0_84 br_0_84 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c84
+ bl_0_84 br_0_84 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c84
+ bl_0_84 br_0_84 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c84
+ bl_0_84 br_0_84 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c84
+ bl_0_84 br_0_84 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c84
+ bl_0_84 br_0_84 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c84
+ bl_0_84 br_0_84 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c84
+ bl_0_84 br_0_84 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c84
+ bl_0_84 br_0_84 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c84
+ bl_0_84 br_0_84 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c84
+ bl_0_84 br_0_84 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c84
+ bl_0_84 br_0_84 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c84
+ bl_0_84 br_0_84 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c84
+ bl_0_84 br_0_84 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c85
+ bl_0_85 br_0_85 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c85
+ bl_0_85 br_0_85 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c85
+ bl_0_85 br_0_85 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c85
+ bl_0_85 br_0_85 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c85
+ bl_0_85 br_0_85 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c85
+ bl_0_85 br_0_85 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c85
+ bl_0_85 br_0_85 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c85
+ bl_0_85 br_0_85 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c85
+ bl_0_85 br_0_85 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c85
+ bl_0_85 br_0_85 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c85
+ bl_0_85 br_0_85 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c85
+ bl_0_85 br_0_85 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c85
+ bl_0_85 br_0_85 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c85
+ bl_0_85 br_0_85 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c85
+ bl_0_85 br_0_85 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c85
+ bl_0_85 br_0_85 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c85
+ bl_0_85 br_0_85 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c85
+ bl_0_85 br_0_85 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c85
+ bl_0_85 br_0_85 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c85
+ bl_0_85 br_0_85 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c85
+ bl_0_85 br_0_85 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c85
+ bl_0_85 br_0_85 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c85
+ bl_0_85 br_0_85 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c85
+ bl_0_85 br_0_85 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c85
+ bl_0_85 br_0_85 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c85
+ bl_0_85 br_0_85 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c85
+ bl_0_85 br_0_85 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c85
+ bl_0_85 br_0_85 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c85
+ bl_0_85 br_0_85 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c85
+ bl_0_85 br_0_85 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c85
+ bl_0_85 br_0_85 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c85
+ bl_0_85 br_0_85 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c85
+ bl_0_85 br_0_85 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c85
+ bl_0_85 br_0_85 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c85
+ bl_0_85 br_0_85 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c85
+ bl_0_85 br_0_85 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c85
+ bl_0_85 br_0_85 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c85
+ bl_0_85 br_0_85 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c85
+ bl_0_85 br_0_85 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c85
+ bl_0_85 br_0_85 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c85
+ bl_0_85 br_0_85 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c85
+ bl_0_85 br_0_85 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c85
+ bl_0_85 br_0_85 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c85
+ bl_0_85 br_0_85 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c86
+ bl_0_86 br_0_86 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c86
+ bl_0_86 br_0_86 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c86
+ bl_0_86 br_0_86 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c86
+ bl_0_86 br_0_86 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c86
+ bl_0_86 br_0_86 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c86
+ bl_0_86 br_0_86 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c86
+ bl_0_86 br_0_86 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c86
+ bl_0_86 br_0_86 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c86
+ bl_0_86 br_0_86 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c86
+ bl_0_86 br_0_86 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c86
+ bl_0_86 br_0_86 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c86
+ bl_0_86 br_0_86 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c86
+ bl_0_86 br_0_86 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c86
+ bl_0_86 br_0_86 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c86
+ bl_0_86 br_0_86 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c86
+ bl_0_86 br_0_86 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c86
+ bl_0_86 br_0_86 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c86
+ bl_0_86 br_0_86 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c86
+ bl_0_86 br_0_86 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c86
+ bl_0_86 br_0_86 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c86
+ bl_0_86 br_0_86 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c86
+ bl_0_86 br_0_86 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c86
+ bl_0_86 br_0_86 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c86
+ bl_0_86 br_0_86 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c86
+ bl_0_86 br_0_86 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c86
+ bl_0_86 br_0_86 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c86
+ bl_0_86 br_0_86 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c86
+ bl_0_86 br_0_86 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c86
+ bl_0_86 br_0_86 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c86
+ bl_0_86 br_0_86 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c86
+ bl_0_86 br_0_86 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c86
+ bl_0_86 br_0_86 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c86
+ bl_0_86 br_0_86 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c86
+ bl_0_86 br_0_86 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c86
+ bl_0_86 br_0_86 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c86
+ bl_0_86 br_0_86 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c86
+ bl_0_86 br_0_86 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c86
+ bl_0_86 br_0_86 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c86
+ bl_0_86 br_0_86 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c86
+ bl_0_86 br_0_86 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c86
+ bl_0_86 br_0_86 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c86
+ bl_0_86 br_0_86 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c86
+ bl_0_86 br_0_86 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c86
+ bl_0_86 br_0_86 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c87
+ bl_0_87 br_0_87 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c87
+ bl_0_87 br_0_87 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c87
+ bl_0_87 br_0_87 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c87
+ bl_0_87 br_0_87 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c87
+ bl_0_87 br_0_87 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c87
+ bl_0_87 br_0_87 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c87
+ bl_0_87 br_0_87 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c87
+ bl_0_87 br_0_87 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c87
+ bl_0_87 br_0_87 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c87
+ bl_0_87 br_0_87 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c87
+ bl_0_87 br_0_87 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c87
+ bl_0_87 br_0_87 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c87
+ bl_0_87 br_0_87 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c87
+ bl_0_87 br_0_87 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c87
+ bl_0_87 br_0_87 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c87
+ bl_0_87 br_0_87 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c87
+ bl_0_87 br_0_87 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c87
+ bl_0_87 br_0_87 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c87
+ bl_0_87 br_0_87 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c87
+ bl_0_87 br_0_87 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c87
+ bl_0_87 br_0_87 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c87
+ bl_0_87 br_0_87 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c87
+ bl_0_87 br_0_87 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c87
+ bl_0_87 br_0_87 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c87
+ bl_0_87 br_0_87 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c87
+ bl_0_87 br_0_87 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c87
+ bl_0_87 br_0_87 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c87
+ bl_0_87 br_0_87 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c87
+ bl_0_87 br_0_87 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c87
+ bl_0_87 br_0_87 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c87
+ bl_0_87 br_0_87 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c87
+ bl_0_87 br_0_87 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c87
+ bl_0_87 br_0_87 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c87
+ bl_0_87 br_0_87 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c87
+ bl_0_87 br_0_87 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c87
+ bl_0_87 br_0_87 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c87
+ bl_0_87 br_0_87 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c87
+ bl_0_87 br_0_87 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c87
+ bl_0_87 br_0_87 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c87
+ bl_0_87 br_0_87 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c87
+ bl_0_87 br_0_87 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c87
+ bl_0_87 br_0_87 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c87
+ bl_0_87 br_0_87 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c87
+ bl_0_87 br_0_87 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c88
+ bl_0_88 br_0_88 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c88
+ bl_0_88 br_0_88 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c88
+ bl_0_88 br_0_88 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c88
+ bl_0_88 br_0_88 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c88
+ bl_0_88 br_0_88 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c88
+ bl_0_88 br_0_88 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c88
+ bl_0_88 br_0_88 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c88
+ bl_0_88 br_0_88 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c88
+ bl_0_88 br_0_88 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c88
+ bl_0_88 br_0_88 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c88
+ bl_0_88 br_0_88 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c88
+ bl_0_88 br_0_88 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c88
+ bl_0_88 br_0_88 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c88
+ bl_0_88 br_0_88 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c88
+ bl_0_88 br_0_88 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c88
+ bl_0_88 br_0_88 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c88
+ bl_0_88 br_0_88 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c88
+ bl_0_88 br_0_88 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c88
+ bl_0_88 br_0_88 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c88
+ bl_0_88 br_0_88 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c88
+ bl_0_88 br_0_88 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c88
+ bl_0_88 br_0_88 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c88
+ bl_0_88 br_0_88 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c88
+ bl_0_88 br_0_88 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c88
+ bl_0_88 br_0_88 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c88
+ bl_0_88 br_0_88 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c88
+ bl_0_88 br_0_88 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c88
+ bl_0_88 br_0_88 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c88
+ bl_0_88 br_0_88 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c88
+ bl_0_88 br_0_88 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c88
+ bl_0_88 br_0_88 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c88
+ bl_0_88 br_0_88 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c88
+ bl_0_88 br_0_88 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c88
+ bl_0_88 br_0_88 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c88
+ bl_0_88 br_0_88 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c88
+ bl_0_88 br_0_88 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c88
+ bl_0_88 br_0_88 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c88
+ bl_0_88 br_0_88 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c88
+ bl_0_88 br_0_88 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c88
+ bl_0_88 br_0_88 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c88
+ bl_0_88 br_0_88 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c88
+ bl_0_88 br_0_88 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c88
+ bl_0_88 br_0_88 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c88
+ bl_0_88 br_0_88 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c89
+ bl_0_89 br_0_89 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c89
+ bl_0_89 br_0_89 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c89
+ bl_0_89 br_0_89 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c89
+ bl_0_89 br_0_89 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c89
+ bl_0_89 br_0_89 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c89
+ bl_0_89 br_0_89 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c89
+ bl_0_89 br_0_89 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c89
+ bl_0_89 br_0_89 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c89
+ bl_0_89 br_0_89 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c89
+ bl_0_89 br_0_89 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c89
+ bl_0_89 br_0_89 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c89
+ bl_0_89 br_0_89 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c89
+ bl_0_89 br_0_89 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c89
+ bl_0_89 br_0_89 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c89
+ bl_0_89 br_0_89 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c89
+ bl_0_89 br_0_89 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c89
+ bl_0_89 br_0_89 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c89
+ bl_0_89 br_0_89 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c89
+ bl_0_89 br_0_89 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c89
+ bl_0_89 br_0_89 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c89
+ bl_0_89 br_0_89 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c89
+ bl_0_89 br_0_89 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c89
+ bl_0_89 br_0_89 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c89
+ bl_0_89 br_0_89 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c89
+ bl_0_89 br_0_89 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c89
+ bl_0_89 br_0_89 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c89
+ bl_0_89 br_0_89 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c89
+ bl_0_89 br_0_89 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c89
+ bl_0_89 br_0_89 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c89
+ bl_0_89 br_0_89 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c89
+ bl_0_89 br_0_89 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c89
+ bl_0_89 br_0_89 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c89
+ bl_0_89 br_0_89 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c89
+ bl_0_89 br_0_89 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c89
+ bl_0_89 br_0_89 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c89
+ bl_0_89 br_0_89 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c89
+ bl_0_89 br_0_89 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c89
+ bl_0_89 br_0_89 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c89
+ bl_0_89 br_0_89 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c89
+ bl_0_89 br_0_89 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c89
+ bl_0_89 br_0_89 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c89
+ bl_0_89 br_0_89 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c89
+ bl_0_89 br_0_89 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c89
+ bl_0_89 br_0_89 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c90
+ bl_0_90 br_0_90 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c90
+ bl_0_90 br_0_90 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c90
+ bl_0_90 br_0_90 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c90
+ bl_0_90 br_0_90 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c90
+ bl_0_90 br_0_90 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c90
+ bl_0_90 br_0_90 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c90
+ bl_0_90 br_0_90 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c90
+ bl_0_90 br_0_90 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c90
+ bl_0_90 br_0_90 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c90
+ bl_0_90 br_0_90 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c90
+ bl_0_90 br_0_90 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c90
+ bl_0_90 br_0_90 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c90
+ bl_0_90 br_0_90 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c90
+ bl_0_90 br_0_90 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c90
+ bl_0_90 br_0_90 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c90
+ bl_0_90 br_0_90 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c90
+ bl_0_90 br_0_90 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c90
+ bl_0_90 br_0_90 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c90
+ bl_0_90 br_0_90 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c90
+ bl_0_90 br_0_90 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c90
+ bl_0_90 br_0_90 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c90
+ bl_0_90 br_0_90 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c90
+ bl_0_90 br_0_90 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c90
+ bl_0_90 br_0_90 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c90
+ bl_0_90 br_0_90 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c90
+ bl_0_90 br_0_90 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c90
+ bl_0_90 br_0_90 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c90
+ bl_0_90 br_0_90 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c90
+ bl_0_90 br_0_90 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c90
+ bl_0_90 br_0_90 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c90
+ bl_0_90 br_0_90 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c90
+ bl_0_90 br_0_90 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c90
+ bl_0_90 br_0_90 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c90
+ bl_0_90 br_0_90 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c90
+ bl_0_90 br_0_90 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c90
+ bl_0_90 br_0_90 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c90
+ bl_0_90 br_0_90 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c90
+ bl_0_90 br_0_90 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c90
+ bl_0_90 br_0_90 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c90
+ bl_0_90 br_0_90 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c90
+ bl_0_90 br_0_90 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c90
+ bl_0_90 br_0_90 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c90
+ bl_0_90 br_0_90 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c90
+ bl_0_90 br_0_90 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c91
+ bl_0_91 br_0_91 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c91
+ bl_0_91 br_0_91 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c91
+ bl_0_91 br_0_91 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c91
+ bl_0_91 br_0_91 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c91
+ bl_0_91 br_0_91 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c91
+ bl_0_91 br_0_91 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c91
+ bl_0_91 br_0_91 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c91
+ bl_0_91 br_0_91 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c91
+ bl_0_91 br_0_91 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c91
+ bl_0_91 br_0_91 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c91
+ bl_0_91 br_0_91 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c91
+ bl_0_91 br_0_91 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c91
+ bl_0_91 br_0_91 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c91
+ bl_0_91 br_0_91 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c91
+ bl_0_91 br_0_91 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c91
+ bl_0_91 br_0_91 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c91
+ bl_0_91 br_0_91 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c91
+ bl_0_91 br_0_91 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c91
+ bl_0_91 br_0_91 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c91
+ bl_0_91 br_0_91 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c91
+ bl_0_91 br_0_91 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c91
+ bl_0_91 br_0_91 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c91
+ bl_0_91 br_0_91 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c91
+ bl_0_91 br_0_91 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c91
+ bl_0_91 br_0_91 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c91
+ bl_0_91 br_0_91 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c91
+ bl_0_91 br_0_91 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c91
+ bl_0_91 br_0_91 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c91
+ bl_0_91 br_0_91 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c91
+ bl_0_91 br_0_91 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c91
+ bl_0_91 br_0_91 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c91
+ bl_0_91 br_0_91 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c91
+ bl_0_91 br_0_91 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c91
+ bl_0_91 br_0_91 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c91
+ bl_0_91 br_0_91 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c91
+ bl_0_91 br_0_91 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c91
+ bl_0_91 br_0_91 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c91
+ bl_0_91 br_0_91 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c91
+ bl_0_91 br_0_91 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c91
+ bl_0_91 br_0_91 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c91
+ bl_0_91 br_0_91 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c91
+ bl_0_91 br_0_91 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c91
+ bl_0_91 br_0_91 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c91
+ bl_0_91 br_0_91 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c92
+ bl_0_92 br_0_92 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c92
+ bl_0_92 br_0_92 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c92
+ bl_0_92 br_0_92 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c92
+ bl_0_92 br_0_92 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c92
+ bl_0_92 br_0_92 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c92
+ bl_0_92 br_0_92 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c92
+ bl_0_92 br_0_92 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c92
+ bl_0_92 br_0_92 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c92
+ bl_0_92 br_0_92 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c92
+ bl_0_92 br_0_92 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c92
+ bl_0_92 br_0_92 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c92
+ bl_0_92 br_0_92 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c92
+ bl_0_92 br_0_92 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c92
+ bl_0_92 br_0_92 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c92
+ bl_0_92 br_0_92 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c92
+ bl_0_92 br_0_92 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c92
+ bl_0_92 br_0_92 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c92
+ bl_0_92 br_0_92 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c92
+ bl_0_92 br_0_92 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c92
+ bl_0_92 br_0_92 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c92
+ bl_0_92 br_0_92 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c92
+ bl_0_92 br_0_92 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c92
+ bl_0_92 br_0_92 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c92
+ bl_0_92 br_0_92 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c92
+ bl_0_92 br_0_92 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c92
+ bl_0_92 br_0_92 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c92
+ bl_0_92 br_0_92 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c92
+ bl_0_92 br_0_92 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c92
+ bl_0_92 br_0_92 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c92
+ bl_0_92 br_0_92 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c92
+ bl_0_92 br_0_92 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c92
+ bl_0_92 br_0_92 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c92
+ bl_0_92 br_0_92 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c92
+ bl_0_92 br_0_92 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c92
+ bl_0_92 br_0_92 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c92
+ bl_0_92 br_0_92 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c92
+ bl_0_92 br_0_92 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c92
+ bl_0_92 br_0_92 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c92
+ bl_0_92 br_0_92 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c92
+ bl_0_92 br_0_92 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c92
+ bl_0_92 br_0_92 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c92
+ bl_0_92 br_0_92 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c92
+ bl_0_92 br_0_92 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c92
+ bl_0_92 br_0_92 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c93
+ bl_0_93 br_0_93 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c93
+ bl_0_93 br_0_93 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c93
+ bl_0_93 br_0_93 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c93
+ bl_0_93 br_0_93 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c93
+ bl_0_93 br_0_93 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c93
+ bl_0_93 br_0_93 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c93
+ bl_0_93 br_0_93 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c93
+ bl_0_93 br_0_93 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c93
+ bl_0_93 br_0_93 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c93
+ bl_0_93 br_0_93 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c93
+ bl_0_93 br_0_93 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c93
+ bl_0_93 br_0_93 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c93
+ bl_0_93 br_0_93 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c93
+ bl_0_93 br_0_93 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c93
+ bl_0_93 br_0_93 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c93
+ bl_0_93 br_0_93 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c93
+ bl_0_93 br_0_93 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c93
+ bl_0_93 br_0_93 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c93
+ bl_0_93 br_0_93 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c93
+ bl_0_93 br_0_93 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c93
+ bl_0_93 br_0_93 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c93
+ bl_0_93 br_0_93 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c93
+ bl_0_93 br_0_93 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c93
+ bl_0_93 br_0_93 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c93
+ bl_0_93 br_0_93 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c93
+ bl_0_93 br_0_93 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c93
+ bl_0_93 br_0_93 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c93
+ bl_0_93 br_0_93 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c93
+ bl_0_93 br_0_93 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c93
+ bl_0_93 br_0_93 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c93
+ bl_0_93 br_0_93 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c93
+ bl_0_93 br_0_93 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c93
+ bl_0_93 br_0_93 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c93
+ bl_0_93 br_0_93 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c93
+ bl_0_93 br_0_93 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c93
+ bl_0_93 br_0_93 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c93
+ bl_0_93 br_0_93 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c93
+ bl_0_93 br_0_93 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c93
+ bl_0_93 br_0_93 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c93
+ bl_0_93 br_0_93 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c93
+ bl_0_93 br_0_93 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c93
+ bl_0_93 br_0_93 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c93
+ bl_0_93 br_0_93 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c93
+ bl_0_93 br_0_93 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c94
+ bl_0_94 br_0_94 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c94
+ bl_0_94 br_0_94 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c94
+ bl_0_94 br_0_94 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c94
+ bl_0_94 br_0_94 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c94
+ bl_0_94 br_0_94 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c94
+ bl_0_94 br_0_94 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c94
+ bl_0_94 br_0_94 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c94
+ bl_0_94 br_0_94 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c94
+ bl_0_94 br_0_94 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c94
+ bl_0_94 br_0_94 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c94
+ bl_0_94 br_0_94 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c94
+ bl_0_94 br_0_94 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c94
+ bl_0_94 br_0_94 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c94
+ bl_0_94 br_0_94 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c94
+ bl_0_94 br_0_94 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c94
+ bl_0_94 br_0_94 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c94
+ bl_0_94 br_0_94 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c94
+ bl_0_94 br_0_94 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c94
+ bl_0_94 br_0_94 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c94
+ bl_0_94 br_0_94 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c94
+ bl_0_94 br_0_94 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c94
+ bl_0_94 br_0_94 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c94
+ bl_0_94 br_0_94 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c94
+ bl_0_94 br_0_94 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c94
+ bl_0_94 br_0_94 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c94
+ bl_0_94 br_0_94 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c94
+ bl_0_94 br_0_94 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c94
+ bl_0_94 br_0_94 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c94
+ bl_0_94 br_0_94 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c94
+ bl_0_94 br_0_94 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c94
+ bl_0_94 br_0_94 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c94
+ bl_0_94 br_0_94 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c94
+ bl_0_94 br_0_94 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c94
+ bl_0_94 br_0_94 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c94
+ bl_0_94 br_0_94 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c94
+ bl_0_94 br_0_94 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c94
+ bl_0_94 br_0_94 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c94
+ bl_0_94 br_0_94 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c94
+ bl_0_94 br_0_94 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c94
+ bl_0_94 br_0_94 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c94
+ bl_0_94 br_0_94 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c94
+ bl_0_94 br_0_94 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c94
+ bl_0_94 br_0_94 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c94
+ bl_0_94 br_0_94 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c95
+ bl_0_95 br_0_95 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c95
+ bl_0_95 br_0_95 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c95
+ bl_0_95 br_0_95 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c95
+ bl_0_95 br_0_95 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c95
+ bl_0_95 br_0_95 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c95
+ bl_0_95 br_0_95 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c95
+ bl_0_95 br_0_95 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c95
+ bl_0_95 br_0_95 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c95
+ bl_0_95 br_0_95 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c95
+ bl_0_95 br_0_95 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c95
+ bl_0_95 br_0_95 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c95
+ bl_0_95 br_0_95 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c95
+ bl_0_95 br_0_95 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c95
+ bl_0_95 br_0_95 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c95
+ bl_0_95 br_0_95 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c95
+ bl_0_95 br_0_95 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c95
+ bl_0_95 br_0_95 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c95
+ bl_0_95 br_0_95 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c95
+ bl_0_95 br_0_95 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c95
+ bl_0_95 br_0_95 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c95
+ bl_0_95 br_0_95 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c95
+ bl_0_95 br_0_95 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c95
+ bl_0_95 br_0_95 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c95
+ bl_0_95 br_0_95 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c95
+ bl_0_95 br_0_95 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c95
+ bl_0_95 br_0_95 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c95
+ bl_0_95 br_0_95 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c95
+ bl_0_95 br_0_95 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c95
+ bl_0_95 br_0_95 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c95
+ bl_0_95 br_0_95 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c95
+ bl_0_95 br_0_95 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c95
+ bl_0_95 br_0_95 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c95
+ bl_0_95 br_0_95 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c95
+ bl_0_95 br_0_95 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c95
+ bl_0_95 br_0_95 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c95
+ bl_0_95 br_0_95 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c95
+ bl_0_95 br_0_95 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c95
+ bl_0_95 br_0_95 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c95
+ bl_0_95 br_0_95 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c95
+ bl_0_95 br_0_95 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c95
+ bl_0_95 br_0_95 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c95
+ bl_0_95 br_0_95 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c95
+ bl_0_95 br_0_95 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c95
+ bl_0_95 br_0_95 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c96
+ bl_0_96 br_0_96 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c96
+ bl_0_96 br_0_96 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c96
+ bl_0_96 br_0_96 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c96
+ bl_0_96 br_0_96 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c96
+ bl_0_96 br_0_96 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c96
+ bl_0_96 br_0_96 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c96
+ bl_0_96 br_0_96 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c96
+ bl_0_96 br_0_96 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c96
+ bl_0_96 br_0_96 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c96
+ bl_0_96 br_0_96 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c96
+ bl_0_96 br_0_96 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c96
+ bl_0_96 br_0_96 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c96
+ bl_0_96 br_0_96 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c96
+ bl_0_96 br_0_96 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c96
+ bl_0_96 br_0_96 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c96
+ bl_0_96 br_0_96 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c96
+ bl_0_96 br_0_96 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c96
+ bl_0_96 br_0_96 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c96
+ bl_0_96 br_0_96 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c96
+ bl_0_96 br_0_96 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c96
+ bl_0_96 br_0_96 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c96
+ bl_0_96 br_0_96 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c96
+ bl_0_96 br_0_96 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c96
+ bl_0_96 br_0_96 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c96
+ bl_0_96 br_0_96 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c96
+ bl_0_96 br_0_96 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c96
+ bl_0_96 br_0_96 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c96
+ bl_0_96 br_0_96 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c96
+ bl_0_96 br_0_96 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c96
+ bl_0_96 br_0_96 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c96
+ bl_0_96 br_0_96 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c96
+ bl_0_96 br_0_96 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c96
+ bl_0_96 br_0_96 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c96
+ bl_0_96 br_0_96 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c96
+ bl_0_96 br_0_96 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c96
+ bl_0_96 br_0_96 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c96
+ bl_0_96 br_0_96 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c96
+ bl_0_96 br_0_96 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c96
+ bl_0_96 br_0_96 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c96
+ bl_0_96 br_0_96 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c96
+ bl_0_96 br_0_96 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c96
+ bl_0_96 br_0_96 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c96
+ bl_0_96 br_0_96 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c96
+ bl_0_96 br_0_96 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c97
+ bl_0_97 br_0_97 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c97
+ bl_0_97 br_0_97 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c97
+ bl_0_97 br_0_97 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c97
+ bl_0_97 br_0_97 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c97
+ bl_0_97 br_0_97 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c97
+ bl_0_97 br_0_97 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c97
+ bl_0_97 br_0_97 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c97
+ bl_0_97 br_0_97 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c97
+ bl_0_97 br_0_97 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c97
+ bl_0_97 br_0_97 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c97
+ bl_0_97 br_0_97 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c97
+ bl_0_97 br_0_97 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c97
+ bl_0_97 br_0_97 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c97
+ bl_0_97 br_0_97 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c97
+ bl_0_97 br_0_97 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c97
+ bl_0_97 br_0_97 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c97
+ bl_0_97 br_0_97 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c97
+ bl_0_97 br_0_97 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c97
+ bl_0_97 br_0_97 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c97
+ bl_0_97 br_0_97 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c97
+ bl_0_97 br_0_97 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c97
+ bl_0_97 br_0_97 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c97
+ bl_0_97 br_0_97 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c97
+ bl_0_97 br_0_97 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c97
+ bl_0_97 br_0_97 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c97
+ bl_0_97 br_0_97 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c97
+ bl_0_97 br_0_97 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c97
+ bl_0_97 br_0_97 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c97
+ bl_0_97 br_0_97 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c97
+ bl_0_97 br_0_97 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c97
+ bl_0_97 br_0_97 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c97
+ bl_0_97 br_0_97 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c97
+ bl_0_97 br_0_97 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c97
+ bl_0_97 br_0_97 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c97
+ bl_0_97 br_0_97 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c97
+ bl_0_97 br_0_97 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c97
+ bl_0_97 br_0_97 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c97
+ bl_0_97 br_0_97 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c97
+ bl_0_97 br_0_97 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c97
+ bl_0_97 br_0_97 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c97
+ bl_0_97 br_0_97 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c97
+ bl_0_97 br_0_97 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c97
+ bl_0_97 br_0_97 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c97
+ bl_0_97 br_0_97 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c98
+ bl_0_98 br_0_98 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c98
+ bl_0_98 br_0_98 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c98
+ bl_0_98 br_0_98 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c98
+ bl_0_98 br_0_98 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c98
+ bl_0_98 br_0_98 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c98
+ bl_0_98 br_0_98 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c98
+ bl_0_98 br_0_98 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c98
+ bl_0_98 br_0_98 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c98
+ bl_0_98 br_0_98 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c98
+ bl_0_98 br_0_98 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c98
+ bl_0_98 br_0_98 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c98
+ bl_0_98 br_0_98 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c98
+ bl_0_98 br_0_98 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c98
+ bl_0_98 br_0_98 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c98
+ bl_0_98 br_0_98 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c98
+ bl_0_98 br_0_98 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c98
+ bl_0_98 br_0_98 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c98
+ bl_0_98 br_0_98 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c98
+ bl_0_98 br_0_98 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c98
+ bl_0_98 br_0_98 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c98
+ bl_0_98 br_0_98 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c98
+ bl_0_98 br_0_98 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c98
+ bl_0_98 br_0_98 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c98
+ bl_0_98 br_0_98 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c98
+ bl_0_98 br_0_98 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c98
+ bl_0_98 br_0_98 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c98
+ bl_0_98 br_0_98 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c98
+ bl_0_98 br_0_98 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c98
+ bl_0_98 br_0_98 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c98
+ bl_0_98 br_0_98 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c98
+ bl_0_98 br_0_98 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c98
+ bl_0_98 br_0_98 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c98
+ bl_0_98 br_0_98 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c98
+ bl_0_98 br_0_98 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c98
+ bl_0_98 br_0_98 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c98
+ bl_0_98 br_0_98 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c98
+ bl_0_98 br_0_98 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c98
+ bl_0_98 br_0_98 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c98
+ bl_0_98 br_0_98 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c98
+ bl_0_98 br_0_98 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c98
+ bl_0_98 br_0_98 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c98
+ bl_0_98 br_0_98 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c98
+ bl_0_98 br_0_98 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c98
+ bl_0_98 br_0_98 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c99
+ bl_0_99 br_0_99 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c99
+ bl_0_99 br_0_99 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c99
+ bl_0_99 br_0_99 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c99
+ bl_0_99 br_0_99 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c99
+ bl_0_99 br_0_99 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c99
+ bl_0_99 br_0_99 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c99
+ bl_0_99 br_0_99 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c99
+ bl_0_99 br_0_99 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c99
+ bl_0_99 br_0_99 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c99
+ bl_0_99 br_0_99 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c99
+ bl_0_99 br_0_99 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c99
+ bl_0_99 br_0_99 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c99
+ bl_0_99 br_0_99 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c99
+ bl_0_99 br_0_99 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c99
+ bl_0_99 br_0_99 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c99
+ bl_0_99 br_0_99 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c99
+ bl_0_99 br_0_99 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c99
+ bl_0_99 br_0_99 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c99
+ bl_0_99 br_0_99 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c99
+ bl_0_99 br_0_99 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c99
+ bl_0_99 br_0_99 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c99
+ bl_0_99 br_0_99 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c99
+ bl_0_99 br_0_99 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c99
+ bl_0_99 br_0_99 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c99
+ bl_0_99 br_0_99 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c99
+ bl_0_99 br_0_99 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c99
+ bl_0_99 br_0_99 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c99
+ bl_0_99 br_0_99 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c99
+ bl_0_99 br_0_99 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c99
+ bl_0_99 br_0_99 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c99
+ bl_0_99 br_0_99 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c99
+ bl_0_99 br_0_99 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c99
+ bl_0_99 br_0_99 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c99
+ bl_0_99 br_0_99 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c99
+ bl_0_99 br_0_99 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c99
+ bl_0_99 br_0_99 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c99
+ bl_0_99 br_0_99 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c99
+ bl_0_99 br_0_99 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c99
+ bl_0_99 br_0_99 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c99
+ bl_0_99 br_0_99 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c99
+ bl_0_99 br_0_99 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c99
+ bl_0_99 br_0_99 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c99
+ bl_0_99 br_0_99 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c99
+ bl_0_99 br_0_99 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c100
+ bl_0_100 br_0_100 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c100
+ bl_0_100 br_0_100 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c100
+ bl_0_100 br_0_100 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c100
+ bl_0_100 br_0_100 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c100
+ bl_0_100 br_0_100 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c100
+ bl_0_100 br_0_100 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c100
+ bl_0_100 br_0_100 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c100
+ bl_0_100 br_0_100 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c100
+ bl_0_100 br_0_100 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c100
+ bl_0_100 br_0_100 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c100
+ bl_0_100 br_0_100 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c100
+ bl_0_100 br_0_100 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c100
+ bl_0_100 br_0_100 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c100
+ bl_0_100 br_0_100 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c100
+ bl_0_100 br_0_100 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c100
+ bl_0_100 br_0_100 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c100
+ bl_0_100 br_0_100 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c100
+ bl_0_100 br_0_100 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c100
+ bl_0_100 br_0_100 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c100
+ bl_0_100 br_0_100 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c100
+ bl_0_100 br_0_100 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c100
+ bl_0_100 br_0_100 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c100
+ bl_0_100 br_0_100 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c100
+ bl_0_100 br_0_100 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c100
+ bl_0_100 br_0_100 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c100
+ bl_0_100 br_0_100 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c100
+ bl_0_100 br_0_100 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c100
+ bl_0_100 br_0_100 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c100
+ bl_0_100 br_0_100 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c100
+ bl_0_100 br_0_100 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c100
+ bl_0_100 br_0_100 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c100
+ bl_0_100 br_0_100 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c100
+ bl_0_100 br_0_100 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c100
+ bl_0_100 br_0_100 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c100
+ bl_0_100 br_0_100 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c100
+ bl_0_100 br_0_100 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c100
+ bl_0_100 br_0_100 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c100
+ bl_0_100 br_0_100 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c100
+ bl_0_100 br_0_100 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c100
+ bl_0_100 br_0_100 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c100
+ bl_0_100 br_0_100 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c100
+ bl_0_100 br_0_100 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c100
+ bl_0_100 br_0_100 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c100
+ bl_0_100 br_0_100 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c101
+ bl_0_101 br_0_101 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c101
+ bl_0_101 br_0_101 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c101
+ bl_0_101 br_0_101 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c101
+ bl_0_101 br_0_101 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c101
+ bl_0_101 br_0_101 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c101
+ bl_0_101 br_0_101 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c101
+ bl_0_101 br_0_101 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c101
+ bl_0_101 br_0_101 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c101
+ bl_0_101 br_0_101 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c101
+ bl_0_101 br_0_101 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c101
+ bl_0_101 br_0_101 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c101
+ bl_0_101 br_0_101 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c101
+ bl_0_101 br_0_101 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c101
+ bl_0_101 br_0_101 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c101
+ bl_0_101 br_0_101 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c101
+ bl_0_101 br_0_101 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c101
+ bl_0_101 br_0_101 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c101
+ bl_0_101 br_0_101 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c101
+ bl_0_101 br_0_101 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c101
+ bl_0_101 br_0_101 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c101
+ bl_0_101 br_0_101 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c101
+ bl_0_101 br_0_101 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c101
+ bl_0_101 br_0_101 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c101
+ bl_0_101 br_0_101 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c101
+ bl_0_101 br_0_101 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c101
+ bl_0_101 br_0_101 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c101
+ bl_0_101 br_0_101 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c101
+ bl_0_101 br_0_101 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c101
+ bl_0_101 br_0_101 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c101
+ bl_0_101 br_0_101 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c101
+ bl_0_101 br_0_101 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c101
+ bl_0_101 br_0_101 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c101
+ bl_0_101 br_0_101 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c101
+ bl_0_101 br_0_101 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c101
+ bl_0_101 br_0_101 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c101
+ bl_0_101 br_0_101 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c101
+ bl_0_101 br_0_101 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c101
+ bl_0_101 br_0_101 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c101
+ bl_0_101 br_0_101 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c101
+ bl_0_101 br_0_101 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c101
+ bl_0_101 br_0_101 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c101
+ bl_0_101 br_0_101 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c101
+ bl_0_101 br_0_101 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c101
+ bl_0_101 br_0_101 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c102
+ bl_0_102 br_0_102 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c102
+ bl_0_102 br_0_102 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c102
+ bl_0_102 br_0_102 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c102
+ bl_0_102 br_0_102 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c102
+ bl_0_102 br_0_102 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c102
+ bl_0_102 br_0_102 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c102
+ bl_0_102 br_0_102 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c102
+ bl_0_102 br_0_102 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c102
+ bl_0_102 br_0_102 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c102
+ bl_0_102 br_0_102 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c102
+ bl_0_102 br_0_102 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c102
+ bl_0_102 br_0_102 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c102
+ bl_0_102 br_0_102 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c102
+ bl_0_102 br_0_102 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c102
+ bl_0_102 br_0_102 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c102
+ bl_0_102 br_0_102 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c102
+ bl_0_102 br_0_102 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c102
+ bl_0_102 br_0_102 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c102
+ bl_0_102 br_0_102 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c102
+ bl_0_102 br_0_102 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c102
+ bl_0_102 br_0_102 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c102
+ bl_0_102 br_0_102 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c102
+ bl_0_102 br_0_102 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c102
+ bl_0_102 br_0_102 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c102
+ bl_0_102 br_0_102 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c102
+ bl_0_102 br_0_102 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c102
+ bl_0_102 br_0_102 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c102
+ bl_0_102 br_0_102 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c102
+ bl_0_102 br_0_102 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c102
+ bl_0_102 br_0_102 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c102
+ bl_0_102 br_0_102 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c102
+ bl_0_102 br_0_102 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c102
+ bl_0_102 br_0_102 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c102
+ bl_0_102 br_0_102 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c102
+ bl_0_102 br_0_102 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c102
+ bl_0_102 br_0_102 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c102
+ bl_0_102 br_0_102 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c102
+ bl_0_102 br_0_102 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c102
+ bl_0_102 br_0_102 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c102
+ bl_0_102 br_0_102 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c102
+ bl_0_102 br_0_102 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c102
+ bl_0_102 br_0_102 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c102
+ bl_0_102 br_0_102 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c102
+ bl_0_102 br_0_102 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c103
+ bl_0_103 br_0_103 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c103
+ bl_0_103 br_0_103 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c103
+ bl_0_103 br_0_103 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c103
+ bl_0_103 br_0_103 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c103
+ bl_0_103 br_0_103 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c103
+ bl_0_103 br_0_103 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c103
+ bl_0_103 br_0_103 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c103
+ bl_0_103 br_0_103 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c103
+ bl_0_103 br_0_103 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c103
+ bl_0_103 br_0_103 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c103
+ bl_0_103 br_0_103 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c103
+ bl_0_103 br_0_103 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c103
+ bl_0_103 br_0_103 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c103
+ bl_0_103 br_0_103 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c103
+ bl_0_103 br_0_103 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c103
+ bl_0_103 br_0_103 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c103
+ bl_0_103 br_0_103 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c103
+ bl_0_103 br_0_103 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c103
+ bl_0_103 br_0_103 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c103
+ bl_0_103 br_0_103 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c103
+ bl_0_103 br_0_103 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c103
+ bl_0_103 br_0_103 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c103
+ bl_0_103 br_0_103 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c103
+ bl_0_103 br_0_103 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c103
+ bl_0_103 br_0_103 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c103
+ bl_0_103 br_0_103 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c103
+ bl_0_103 br_0_103 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c103
+ bl_0_103 br_0_103 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c103
+ bl_0_103 br_0_103 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c103
+ bl_0_103 br_0_103 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c103
+ bl_0_103 br_0_103 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c103
+ bl_0_103 br_0_103 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c103
+ bl_0_103 br_0_103 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c103
+ bl_0_103 br_0_103 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c103
+ bl_0_103 br_0_103 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c103
+ bl_0_103 br_0_103 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c103
+ bl_0_103 br_0_103 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c103
+ bl_0_103 br_0_103 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c103
+ bl_0_103 br_0_103 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c103
+ bl_0_103 br_0_103 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c103
+ bl_0_103 br_0_103 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c103
+ bl_0_103 br_0_103 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c103
+ bl_0_103 br_0_103 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c103
+ bl_0_103 br_0_103 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c104
+ bl_0_104 br_0_104 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c104
+ bl_0_104 br_0_104 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c104
+ bl_0_104 br_0_104 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c104
+ bl_0_104 br_0_104 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c104
+ bl_0_104 br_0_104 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c104
+ bl_0_104 br_0_104 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c104
+ bl_0_104 br_0_104 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c104
+ bl_0_104 br_0_104 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c104
+ bl_0_104 br_0_104 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c104
+ bl_0_104 br_0_104 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c104
+ bl_0_104 br_0_104 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c104
+ bl_0_104 br_0_104 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c104
+ bl_0_104 br_0_104 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c104
+ bl_0_104 br_0_104 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c104
+ bl_0_104 br_0_104 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c104
+ bl_0_104 br_0_104 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c104
+ bl_0_104 br_0_104 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c104
+ bl_0_104 br_0_104 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c104
+ bl_0_104 br_0_104 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c104
+ bl_0_104 br_0_104 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c104
+ bl_0_104 br_0_104 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c104
+ bl_0_104 br_0_104 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c104
+ bl_0_104 br_0_104 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c104
+ bl_0_104 br_0_104 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c104
+ bl_0_104 br_0_104 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c104
+ bl_0_104 br_0_104 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c104
+ bl_0_104 br_0_104 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c104
+ bl_0_104 br_0_104 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c104
+ bl_0_104 br_0_104 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c104
+ bl_0_104 br_0_104 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c104
+ bl_0_104 br_0_104 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c104
+ bl_0_104 br_0_104 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c104
+ bl_0_104 br_0_104 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c104
+ bl_0_104 br_0_104 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c104
+ bl_0_104 br_0_104 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c104
+ bl_0_104 br_0_104 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c104
+ bl_0_104 br_0_104 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c104
+ bl_0_104 br_0_104 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c104
+ bl_0_104 br_0_104 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c104
+ bl_0_104 br_0_104 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c104
+ bl_0_104 br_0_104 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c104
+ bl_0_104 br_0_104 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c104
+ bl_0_104 br_0_104 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c104
+ bl_0_104 br_0_104 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c105
+ bl_0_105 br_0_105 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c105
+ bl_0_105 br_0_105 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c105
+ bl_0_105 br_0_105 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c105
+ bl_0_105 br_0_105 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c105
+ bl_0_105 br_0_105 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c105
+ bl_0_105 br_0_105 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c105
+ bl_0_105 br_0_105 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c105
+ bl_0_105 br_0_105 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c105
+ bl_0_105 br_0_105 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c105
+ bl_0_105 br_0_105 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c105
+ bl_0_105 br_0_105 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c105
+ bl_0_105 br_0_105 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c105
+ bl_0_105 br_0_105 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c105
+ bl_0_105 br_0_105 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c105
+ bl_0_105 br_0_105 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c105
+ bl_0_105 br_0_105 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c105
+ bl_0_105 br_0_105 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c105
+ bl_0_105 br_0_105 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c105
+ bl_0_105 br_0_105 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c105
+ bl_0_105 br_0_105 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c105
+ bl_0_105 br_0_105 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c105
+ bl_0_105 br_0_105 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c105
+ bl_0_105 br_0_105 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c105
+ bl_0_105 br_0_105 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c105
+ bl_0_105 br_0_105 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c105
+ bl_0_105 br_0_105 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c105
+ bl_0_105 br_0_105 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c105
+ bl_0_105 br_0_105 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c105
+ bl_0_105 br_0_105 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c105
+ bl_0_105 br_0_105 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c105
+ bl_0_105 br_0_105 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c105
+ bl_0_105 br_0_105 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c105
+ bl_0_105 br_0_105 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c105
+ bl_0_105 br_0_105 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c105
+ bl_0_105 br_0_105 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c105
+ bl_0_105 br_0_105 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c105
+ bl_0_105 br_0_105 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c105
+ bl_0_105 br_0_105 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c105
+ bl_0_105 br_0_105 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c105
+ bl_0_105 br_0_105 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c105
+ bl_0_105 br_0_105 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c105
+ bl_0_105 br_0_105 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c105
+ bl_0_105 br_0_105 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c105
+ bl_0_105 br_0_105 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c106
+ bl_0_106 br_0_106 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c106
+ bl_0_106 br_0_106 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c106
+ bl_0_106 br_0_106 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c106
+ bl_0_106 br_0_106 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c106
+ bl_0_106 br_0_106 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c106
+ bl_0_106 br_0_106 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c106
+ bl_0_106 br_0_106 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c106
+ bl_0_106 br_0_106 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c106
+ bl_0_106 br_0_106 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c106
+ bl_0_106 br_0_106 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c106
+ bl_0_106 br_0_106 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c106
+ bl_0_106 br_0_106 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c106
+ bl_0_106 br_0_106 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c106
+ bl_0_106 br_0_106 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c106
+ bl_0_106 br_0_106 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c106
+ bl_0_106 br_0_106 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c106
+ bl_0_106 br_0_106 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c106
+ bl_0_106 br_0_106 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c106
+ bl_0_106 br_0_106 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c106
+ bl_0_106 br_0_106 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c106
+ bl_0_106 br_0_106 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c106
+ bl_0_106 br_0_106 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c106
+ bl_0_106 br_0_106 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c106
+ bl_0_106 br_0_106 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c106
+ bl_0_106 br_0_106 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c106
+ bl_0_106 br_0_106 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c106
+ bl_0_106 br_0_106 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c106
+ bl_0_106 br_0_106 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c106
+ bl_0_106 br_0_106 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c106
+ bl_0_106 br_0_106 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c106
+ bl_0_106 br_0_106 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c106
+ bl_0_106 br_0_106 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c106
+ bl_0_106 br_0_106 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c106
+ bl_0_106 br_0_106 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c106
+ bl_0_106 br_0_106 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c106
+ bl_0_106 br_0_106 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c106
+ bl_0_106 br_0_106 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c106
+ bl_0_106 br_0_106 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c106
+ bl_0_106 br_0_106 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c106
+ bl_0_106 br_0_106 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c106
+ bl_0_106 br_0_106 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c106
+ bl_0_106 br_0_106 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c106
+ bl_0_106 br_0_106 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c106
+ bl_0_106 br_0_106 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c107
+ bl_0_107 br_0_107 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c107
+ bl_0_107 br_0_107 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c107
+ bl_0_107 br_0_107 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c107
+ bl_0_107 br_0_107 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c107
+ bl_0_107 br_0_107 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c107
+ bl_0_107 br_0_107 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c107
+ bl_0_107 br_0_107 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c107
+ bl_0_107 br_0_107 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c107
+ bl_0_107 br_0_107 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c107
+ bl_0_107 br_0_107 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c107
+ bl_0_107 br_0_107 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c107
+ bl_0_107 br_0_107 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c107
+ bl_0_107 br_0_107 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c107
+ bl_0_107 br_0_107 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c107
+ bl_0_107 br_0_107 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c107
+ bl_0_107 br_0_107 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c107
+ bl_0_107 br_0_107 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c107
+ bl_0_107 br_0_107 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c107
+ bl_0_107 br_0_107 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c107
+ bl_0_107 br_0_107 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c107
+ bl_0_107 br_0_107 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c107
+ bl_0_107 br_0_107 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c107
+ bl_0_107 br_0_107 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c107
+ bl_0_107 br_0_107 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c107
+ bl_0_107 br_0_107 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c107
+ bl_0_107 br_0_107 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c107
+ bl_0_107 br_0_107 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c107
+ bl_0_107 br_0_107 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c107
+ bl_0_107 br_0_107 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c107
+ bl_0_107 br_0_107 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c107
+ bl_0_107 br_0_107 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c107
+ bl_0_107 br_0_107 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c107
+ bl_0_107 br_0_107 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c107
+ bl_0_107 br_0_107 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c107
+ bl_0_107 br_0_107 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c107
+ bl_0_107 br_0_107 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c107
+ bl_0_107 br_0_107 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c107
+ bl_0_107 br_0_107 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c107
+ bl_0_107 br_0_107 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c107
+ bl_0_107 br_0_107 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c107
+ bl_0_107 br_0_107 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c107
+ bl_0_107 br_0_107 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c107
+ bl_0_107 br_0_107 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c107
+ bl_0_107 br_0_107 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c108
+ bl_0_108 br_0_108 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c108
+ bl_0_108 br_0_108 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c108
+ bl_0_108 br_0_108 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c108
+ bl_0_108 br_0_108 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c108
+ bl_0_108 br_0_108 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c108
+ bl_0_108 br_0_108 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c108
+ bl_0_108 br_0_108 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c108
+ bl_0_108 br_0_108 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c108
+ bl_0_108 br_0_108 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c108
+ bl_0_108 br_0_108 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c108
+ bl_0_108 br_0_108 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c108
+ bl_0_108 br_0_108 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c108
+ bl_0_108 br_0_108 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c108
+ bl_0_108 br_0_108 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c108
+ bl_0_108 br_0_108 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c108
+ bl_0_108 br_0_108 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c108
+ bl_0_108 br_0_108 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c108
+ bl_0_108 br_0_108 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c108
+ bl_0_108 br_0_108 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c108
+ bl_0_108 br_0_108 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c108
+ bl_0_108 br_0_108 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c108
+ bl_0_108 br_0_108 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c108
+ bl_0_108 br_0_108 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c108
+ bl_0_108 br_0_108 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c108
+ bl_0_108 br_0_108 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c108
+ bl_0_108 br_0_108 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c108
+ bl_0_108 br_0_108 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c108
+ bl_0_108 br_0_108 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c108
+ bl_0_108 br_0_108 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c108
+ bl_0_108 br_0_108 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c108
+ bl_0_108 br_0_108 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c108
+ bl_0_108 br_0_108 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c108
+ bl_0_108 br_0_108 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c108
+ bl_0_108 br_0_108 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c108
+ bl_0_108 br_0_108 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c108
+ bl_0_108 br_0_108 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c108
+ bl_0_108 br_0_108 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c108
+ bl_0_108 br_0_108 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c108
+ bl_0_108 br_0_108 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c108
+ bl_0_108 br_0_108 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c108
+ bl_0_108 br_0_108 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c108
+ bl_0_108 br_0_108 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c108
+ bl_0_108 br_0_108 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c108
+ bl_0_108 br_0_108 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c109
+ bl_0_109 br_0_109 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c109
+ bl_0_109 br_0_109 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c109
+ bl_0_109 br_0_109 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c109
+ bl_0_109 br_0_109 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c109
+ bl_0_109 br_0_109 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c109
+ bl_0_109 br_0_109 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c109
+ bl_0_109 br_0_109 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c109
+ bl_0_109 br_0_109 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c109
+ bl_0_109 br_0_109 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c109
+ bl_0_109 br_0_109 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c109
+ bl_0_109 br_0_109 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c109
+ bl_0_109 br_0_109 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c109
+ bl_0_109 br_0_109 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c109
+ bl_0_109 br_0_109 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c109
+ bl_0_109 br_0_109 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c109
+ bl_0_109 br_0_109 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c109
+ bl_0_109 br_0_109 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c109
+ bl_0_109 br_0_109 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c109
+ bl_0_109 br_0_109 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c109
+ bl_0_109 br_0_109 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c109
+ bl_0_109 br_0_109 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c109
+ bl_0_109 br_0_109 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c109
+ bl_0_109 br_0_109 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c109
+ bl_0_109 br_0_109 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c109
+ bl_0_109 br_0_109 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c109
+ bl_0_109 br_0_109 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c109
+ bl_0_109 br_0_109 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c109
+ bl_0_109 br_0_109 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c109
+ bl_0_109 br_0_109 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c109
+ bl_0_109 br_0_109 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c109
+ bl_0_109 br_0_109 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c109
+ bl_0_109 br_0_109 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c109
+ bl_0_109 br_0_109 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c109
+ bl_0_109 br_0_109 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c109
+ bl_0_109 br_0_109 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c109
+ bl_0_109 br_0_109 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c109
+ bl_0_109 br_0_109 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c109
+ bl_0_109 br_0_109 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c109
+ bl_0_109 br_0_109 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c109
+ bl_0_109 br_0_109 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c109
+ bl_0_109 br_0_109 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c109
+ bl_0_109 br_0_109 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c109
+ bl_0_109 br_0_109 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c109
+ bl_0_109 br_0_109 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c110
+ bl_0_110 br_0_110 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c110
+ bl_0_110 br_0_110 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c110
+ bl_0_110 br_0_110 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c110
+ bl_0_110 br_0_110 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c110
+ bl_0_110 br_0_110 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c110
+ bl_0_110 br_0_110 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c110
+ bl_0_110 br_0_110 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c110
+ bl_0_110 br_0_110 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c110
+ bl_0_110 br_0_110 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c110
+ bl_0_110 br_0_110 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c110
+ bl_0_110 br_0_110 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c110
+ bl_0_110 br_0_110 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c110
+ bl_0_110 br_0_110 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c110
+ bl_0_110 br_0_110 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c110
+ bl_0_110 br_0_110 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c110
+ bl_0_110 br_0_110 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c110
+ bl_0_110 br_0_110 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c110
+ bl_0_110 br_0_110 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c110
+ bl_0_110 br_0_110 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c110
+ bl_0_110 br_0_110 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c110
+ bl_0_110 br_0_110 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c110
+ bl_0_110 br_0_110 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c110
+ bl_0_110 br_0_110 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c110
+ bl_0_110 br_0_110 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c110
+ bl_0_110 br_0_110 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c110
+ bl_0_110 br_0_110 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c110
+ bl_0_110 br_0_110 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c110
+ bl_0_110 br_0_110 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c110
+ bl_0_110 br_0_110 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c110
+ bl_0_110 br_0_110 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c110
+ bl_0_110 br_0_110 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c110
+ bl_0_110 br_0_110 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c110
+ bl_0_110 br_0_110 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c110
+ bl_0_110 br_0_110 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c110
+ bl_0_110 br_0_110 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c110
+ bl_0_110 br_0_110 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c110
+ bl_0_110 br_0_110 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c110
+ bl_0_110 br_0_110 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c110
+ bl_0_110 br_0_110 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c110
+ bl_0_110 br_0_110 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c110
+ bl_0_110 br_0_110 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c110
+ bl_0_110 br_0_110 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c110
+ bl_0_110 br_0_110 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c110
+ bl_0_110 br_0_110 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c111
+ bl_0_111 br_0_111 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c111
+ bl_0_111 br_0_111 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c111
+ bl_0_111 br_0_111 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c111
+ bl_0_111 br_0_111 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c111
+ bl_0_111 br_0_111 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c111
+ bl_0_111 br_0_111 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c111
+ bl_0_111 br_0_111 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c111
+ bl_0_111 br_0_111 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c111
+ bl_0_111 br_0_111 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c111
+ bl_0_111 br_0_111 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c111
+ bl_0_111 br_0_111 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c111
+ bl_0_111 br_0_111 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c111
+ bl_0_111 br_0_111 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c111
+ bl_0_111 br_0_111 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c111
+ bl_0_111 br_0_111 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c111
+ bl_0_111 br_0_111 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c111
+ bl_0_111 br_0_111 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c111
+ bl_0_111 br_0_111 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c111
+ bl_0_111 br_0_111 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c111
+ bl_0_111 br_0_111 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c111
+ bl_0_111 br_0_111 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c111
+ bl_0_111 br_0_111 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c111
+ bl_0_111 br_0_111 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c111
+ bl_0_111 br_0_111 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c111
+ bl_0_111 br_0_111 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c111
+ bl_0_111 br_0_111 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c111
+ bl_0_111 br_0_111 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c111
+ bl_0_111 br_0_111 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c111
+ bl_0_111 br_0_111 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c111
+ bl_0_111 br_0_111 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c111
+ bl_0_111 br_0_111 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c111
+ bl_0_111 br_0_111 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c111
+ bl_0_111 br_0_111 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c111
+ bl_0_111 br_0_111 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c111
+ bl_0_111 br_0_111 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c111
+ bl_0_111 br_0_111 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c111
+ bl_0_111 br_0_111 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c111
+ bl_0_111 br_0_111 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c111
+ bl_0_111 br_0_111 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c111
+ bl_0_111 br_0_111 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c111
+ bl_0_111 br_0_111 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c111
+ bl_0_111 br_0_111 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c111
+ bl_0_111 br_0_111 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c111
+ bl_0_111 br_0_111 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c112
+ bl_0_112 br_0_112 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c112
+ bl_0_112 br_0_112 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c112
+ bl_0_112 br_0_112 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c112
+ bl_0_112 br_0_112 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c112
+ bl_0_112 br_0_112 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c112
+ bl_0_112 br_0_112 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c112
+ bl_0_112 br_0_112 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c112
+ bl_0_112 br_0_112 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c112
+ bl_0_112 br_0_112 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c112
+ bl_0_112 br_0_112 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c112
+ bl_0_112 br_0_112 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c112
+ bl_0_112 br_0_112 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c112
+ bl_0_112 br_0_112 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c112
+ bl_0_112 br_0_112 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c112
+ bl_0_112 br_0_112 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c112
+ bl_0_112 br_0_112 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c112
+ bl_0_112 br_0_112 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c112
+ bl_0_112 br_0_112 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c112
+ bl_0_112 br_0_112 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c112
+ bl_0_112 br_0_112 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c112
+ bl_0_112 br_0_112 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c112
+ bl_0_112 br_0_112 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c112
+ bl_0_112 br_0_112 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c112
+ bl_0_112 br_0_112 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c112
+ bl_0_112 br_0_112 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c112
+ bl_0_112 br_0_112 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c112
+ bl_0_112 br_0_112 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c112
+ bl_0_112 br_0_112 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c112
+ bl_0_112 br_0_112 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c112
+ bl_0_112 br_0_112 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c112
+ bl_0_112 br_0_112 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c112
+ bl_0_112 br_0_112 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c112
+ bl_0_112 br_0_112 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c112
+ bl_0_112 br_0_112 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c112
+ bl_0_112 br_0_112 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c112
+ bl_0_112 br_0_112 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c112
+ bl_0_112 br_0_112 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c112
+ bl_0_112 br_0_112 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c112
+ bl_0_112 br_0_112 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c112
+ bl_0_112 br_0_112 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c112
+ bl_0_112 br_0_112 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c112
+ bl_0_112 br_0_112 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c112
+ bl_0_112 br_0_112 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c112
+ bl_0_112 br_0_112 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c113
+ bl_0_113 br_0_113 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c113
+ bl_0_113 br_0_113 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c113
+ bl_0_113 br_0_113 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c113
+ bl_0_113 br_0_113 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c113
+ bl_0_113 br_0_113 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c113
+ bl_0_113 br_0_113 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c113
+ bl_0_113 br_0_113 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c113
+ bl_0_113 br_0_113 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c113
+ bl_0_113 br_0_113 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c113
+ bl_0_113 br_0_113 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c113
+ bl_0_113 br_0_113 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c113
+ bl_0_113 br_0_113 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c113
+ bl_0_113 br_0_113 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c113
+ bl_0_113 br_0_113 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c113
+ bl_0_113 br_0_113 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c113
+ bl_0_113 br_0_113 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c113
+ bl_0_113 br_0_113 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c113
+ bl_0_113 br_0_113 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c113
+ bl_0_113 br_0_113 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c113
+ bl_0_113 br_0_113 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c113
+ bl_0_113 br_0_113 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c113
+ bl_0_113 br_0_113 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c113
+ bl_0_113 br_0_113 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c113
+ bl_0_113 br_0_113 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c113
+ bl_0_113 br_0_113 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c113
+ bl_0_113 br_0_113 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c113
+ bl_0_113 br_0_113 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c113
+ bl_0_113 br_0_113 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c113
+ bl_0_113 br_0_113 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c113
+ bl_0_113 br_0_113 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c113
+ bl_0_113 br_0_113 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c113
+ bl_0_113 br_0_113 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c113
+ bl_0_113 br_0_113 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c113
+ bl_0_113 br_0_113 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c113
+ bl_0_113 br_0_113 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c113
+ bl_0_113 br_0_113 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c113
+ bl_0_113 br_0_113 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c113
+ bl_0_113 br_0_113 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c113
+ bl_0_113 br_0_113 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c113
+ bl_0_113 br_0_113 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c113
+ bl_0_113 br_0_113 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c113
+ bl_0_113 br_0_113 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c113
+ bl_0_113 br_0_113 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c113
+ bl_0_113 br_0_113 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c114
+ bl_0_114 br_0_114 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c114
+ bl_0_114 br_0_114 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c114
+ bl_0_114 br_0_114 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c114
+ bl_0_114 br_0_114 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c114
+ bl_0_114 br_0_114 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c114
+ bl_0_114 br_0_114 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c114
+ bl_0_114 br_0_114 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c114
+ bl_0_114 br_0_114 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c114
+ bl_0_114 br_0_114 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c114
+ bl_0_114 br_0_114 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c114
+ bl_0_114 br_0_114 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c114
+ bl_0_114 br_0_114 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c114
+ bl_0_114 br_0_114 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c114
+ bl_0_114 br_0_114 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c114
+ bl_0_114 br_0_114 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c114
+ bl_0_114 br_0_114 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c114
+ bl_0_114 br_0_114 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c114
+ bl_0_114 br_0_114 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c114
+ bl_0_114 br_0_114 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c114
+ bl_0_114 br_0_114 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c114
+ bl_0_114 br_0_114 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c114
+ bl_0_114 br_0_114 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c114
+ bl_0_114 br_0_114 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c114
+ bl_0_114 br_0_114 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c114
+ bl_0_114 br_0_114 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c114
+ bl_0_114 br_0_114 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c114
+ bl_0_114 br_0_114 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c114
+ bl_0_114 br_0_114 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c114
+ bl_0_114 br_0_114 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c114
+ bl_0_114 br_0_114 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c114
+ bl_0_114 br_0_114 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c114
+ bl_0_114 br_0_114 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c114
+ bl_0_114 br_0_114 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c114
+ bl_0_114 br_0_114 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c114
+ bl_0_114 br_0_114 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c114
+ bl_0_114 br_0_114 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c114
+ bl_0_114 br_0_114 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c114
+ bl_0_114 br_0_114 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c114
+ bl_0_114 br_0_114 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c114
+ bl_0_114 br_0_114 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c114
+ bl_0_114 br_0_114 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c114
+ bl_0_114 br_0_114 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c114
+ bl_0_114 br_0_114 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c114
+ bl_0_114 br_0_114 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c115
+ bl_0_115 br_0_115 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c115
+ bl_0_115 br_0_115 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c115
+ bl_0_115 br_0_115 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c115
+ bl_0_115 br_0_115 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c115
+ bl_0_115 br_0_115 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c115
+ bl_0_115 br_0_115 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c115
+ bl_0_115 br_0_115 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c115
+ bl_0_115 br_0_115 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c115
+ bl_0_115 br_0_115 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c115
+ bl_0_115 br_0_115 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c115
+ bl_0_115 br_0_115 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c115
+ bl_0_115 br_0_115 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c115
+ bl_0_115 br_0_115 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c115
+ bl_0_115 br_0_115 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c115
+ bl_0_115 br_0_115 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c115
+ bl_0_115 br_0_115 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c115
+ bl_0_115 br_0_115 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c115
+ bl_0_115 br_0_115 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c115
+ bl_0_115 br_0_115 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c115
+ bl_0_115 br_0_115 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c115
+ bl_0_115 br_0_115 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c115
+ bl_0_115 br_0_115 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c115
+ bl_0_115 br_0_115 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c115
+ bl_0_115 br_0_115 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c115
+ bl_0_115 br_0_115 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c115
+ bl_0_115 br_0_115 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c115
+ bl_0_115 br_0_115 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c115
+ bl_0_115 br_0_115 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c115
+ bl_0_115 br_0_115 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c115
+ bl_0_115 br_0_115 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c115
+ bl_0_115 br_0_115 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c115
+ bl_0_115 br_0_115 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c115
+ bl_0_115 br_0_115 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c115
+ bl_0_115 br_0_115 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c115
+ bl_0_115 br_0_115 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c115
+ bl_0_115 br_0_115 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c115
+ bl_0_115 br_0_115 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c115
+ bl_0_115 br_0_115 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c115
+ bl_0_115 br_0_115 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c115
+ bl_0_115 br_0_115 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c115
+ bl_0_115 br_0_115 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c115
+ bl_0_115 br_0_115 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c115
+ bl_0_115 br_0_115 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c115
+ bl_0_115 br_0_115 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c116
+ bl_0_116 br_0_116 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c116
+ bl_0_116 br_0_116 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c116
+ bl_0_116 br_0_116 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c116
+ bl_0_116 br_0_116 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c116
+ bl_0_116 br_0_116 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c116
+ bl_0_116 br_0_116 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c116
+ bl_0_116 br_0_116 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c116
+ bl_0_116 br_0_116 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c116
+ bl_0_116 br_0_116 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c116
+ bl_0_116 br_0_116 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c116
+ bl_0_116 br_0_116 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c116
+ bl_0_116 br_0_116 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c116
+ bl_0_116 br_0_116 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c116
+ bl_0_116 br_0_116 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c116
+ bl_0_116 br_0_116 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c116
+ bl_0_116 br_0_116 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c116
+ bl_0_116 br_0_116 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c116
+ bl_0_116 br_0_116 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c116
+ bl_0_116 br_0_116 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c116
+ bl_0_116 br_0_116 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c116
+ bl_0_116 br_0_116 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c116
+ bl_0_116 br_0_116 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c116
+ bl_0_116 br_0_116 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c116
+ bl_0_116 br_0_116 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c116
+ bl_0_116 br_0_116 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c116
+ bl_0_116 br_0_116 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c116
+ bl_0_116 br_0_116 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c116
+ bl_0_116 br_0_116 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c116
+ bl_0_116 br_0_116 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c116
+ bl_0_116 br_0_116 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c116
+ bl_0_116 br_0_116 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c116
+ bl_0_116 br_0_116 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c116
+ bl_0_116 br_0_116 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c116
+ bl_0_116 br_0_116 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c116
+ bl_0_116 br_0_116 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c116
+ bl_0_116 br_0_116 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c116
+ bl_0_116 br_0_116 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c116
+ bl_0_116 br_0_116 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c116
+ bl_0_116 br_0_116 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c116
+ bl_0_116 br_0_116 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c116
+ bl_0_116 br_0_116 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c116
+ bl_0_116 br_0_116 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c116
+ bl_0_116 br_0_116 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c116
+ bl_0_116 br_0_116 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c117
+ bl_0_117 br_0_117 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c117
+ bl_0_117 br_0_117 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c117
+ bl_0_117 br_0_117 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c117
+ bl_0_117 br_0_117 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c117
+ bl_0_117 br_0_117 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c117
+ bl_0_117 br_0_117 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c117
+ bl_0_117 br_0_117 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c117
+ bl_0_117 br_0_117 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c117
+ bl_0_117 br_0_117 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c117
+ bl_0_117 br_0_117 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c117
+ bl_0_117 br_0_117 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c117
+ bl_0_117 br_0_117 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c117
+ bl_0_117 br_0_117 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c117
+ bl_0_117 br_0_117 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c117
+ bl_0_117 br_0_117 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c117
+ bl_0_117 br_0_117 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c117
+ bl_0_117 br_0_117 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c117
+ bl_0_117 br_0_117 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c117
+ bl_0_117 br_0_117 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c117
+ bl_0_117 br_0_117 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c117
+ bl_0_117 br_0_117 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c117
+ bl_0_117 br_0_117 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c117
+ bl_0_117 br_0_117 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c117
+ bl_0_117 br_0_117 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c117
+ bl_0_117 br_0_117 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c117
+ bl_0_117 br_0_117 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c117
+ bl_0_117 br_0_117 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c117
+ bl_0_117 br_0_117 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c117
+ bl_0_117 br_0_117 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c117
+ bl_0_117 br_0_117 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c117
+ bl_0_117 br_0_117 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c117
+ bl_0_117 br_0_117 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c117
+ bl_0_117 br_0_117 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c117
+ bl_0_117 br_0_117 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c117
+ bl_0_117 br_0_117 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c117
+ bl_0_117 br_0_117 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c117
+ bl_0_117 br_0_117 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c117
+ bl_0_117 br_0_117 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c117
+ bl_0_117 br_0_117 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c117
+ bl_0_117 br_0_117 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c117
+ bl_0_117 br_0_117 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c117
+ bl_0_117 br_0_117 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c117
+ bl_0_117 br_0_117 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c117
+ bl_0_117 br_0_117 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c118
+ bl_0_118 br_0_118 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c118
+ bl_0_118 br_0_118 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c118
+ bl_0_118 br_0_118 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c118
+ bl_0_118 br_0_118 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c118
+ bl_0_118 br_0_118 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c118
+ bl_0_118 br_0_118 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c118
+ bl_0_118 br_0_118 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c118
+ bl_0_118 br_0_118 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c118
+ bl_0_118 br_0_118 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c118
+ bl_0_118 br_0_118 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c118
+ bl_0_118 br_0_118 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c118
+ bl_0_118 br_0_118 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c118
+ bl_0_118 br_0_118 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c118
+ bl_0_118 br_0_118 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c118
+ bl_0_118 br_0_118 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c118
+ bl_0_118 br_0_118 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c118
+ bl_0_118 br_0_118 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c118
+ bl_0_118 br_0_118 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c118
+ bl_0_118 br_0_118 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c118
+ bl_0_118 br_0_118 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c118
+ bl_0_118 br_0_118 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c118
+ bl_0_118 br_0_118 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c118
+ bl_0_118 br_0_118 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c118
+ bl_0_118 br_0_118 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c118
+ bl_0_118 br_0_118 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c118
+ bl_0_118 br_0_118 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c118
+ bl_0_118 br_0_118 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c118
+ bl_0_118 br_0_118 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c118
+ bl_0_118 br_0_118 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c118
+ bl_0_118 br_0_118 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c118
+ bl_0_118 br_0_118 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c118
+ bl_0_118 br_0_118 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c118
+ bl_0_118 br_0_118 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c118
+ bl_0_118 br_0_118 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c118
+ bl_0_118 br_0_118 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c118
+ bl_0_118 br_0_118 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c118
+ bl_0_118 br_0_118 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c118
+ bl_0_118 br_0_118 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c118
+ bl_0_118 br_0_118 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c118
+ bl_0_118 br_0_118 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c118
+ bl_0_118 br_0_118 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c118
+ bl_0_118 br_0_118 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c118
+ bl_0_118 br_0_118 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c118
+ bl_0_118 br_0_118 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c119
+ bl_0_119 br_0_119 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c119
+ bl_0_119 br_0_119 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c119
+ bl_0_119 br_0_119 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c119
+ bl_0_119 br_0_119 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c119
+ bl_0_119 br_0_119 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c119
+ bl_0_119 br_0_119 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c119
+ bl_0_119 br_0_119 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c119
+ bl_0_119 br_0_119 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c119
+ bl_0_119 br_0_119 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c119
+ bl_0_119 br_0_119 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c119
+ bl_0_119 br_0_119 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c119
+ bl_0_119 br_0_119 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c119
+ bl_0_119 br_0_119 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c119
+ bl_0_119 br_0_119 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c119
+ bl_0_119 br_0_119 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c119
+ bl_0_119 br_0_119 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c119
+ bl_0_119 br_0_119 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c119
+ bl_0_119 br_0_119 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c119
+ bl_0_119 br_0_119 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c119
+ bl_0_119 br_0_119 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c119
+ bl_0_119 br_0_119 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c119
+ bl_0_119 br_0_119 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c119
+ bl_0_119 br_0_119 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c119
+ bl_0_119 br_0_119 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c119
+ bl_0_119 br_0_119 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c119
+ bl_0_119 br_0_119 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c119
+ bl_0_119 br_0_119 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c119
+ bl_0_119 br_0_119 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c119
+ bl_0_119 br_0_119 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c119
+ bl_0_119 br_0_119 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c119
+ bl_0_119 br_0_119 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c119
+ bl_0_119 br_0_119 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c119
+ bl_0_119 br_0_119 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c119
+ bl_0_119 br_0_119 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c119
+ bl_0_119 br_0_119 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c119
+ bl_0_119 br_0_119 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c119
+ bl_0_119 br_0_119 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c119
+ bl_0_119 br_0_119 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c119
+ bl_0_119 br_0_119 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c119
+ bl_0_119 br_0_119 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c119
+ bl_0_119 br_0_119 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c119
+ bl_0_119 br_0_119 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c119
+ bl_0_119 br_0_119 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c119
+ bl_0_119 br_0_119 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c120
+ bl_0_120 br_0_120 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c120
+ bl_0_120 br_0_120 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c120
+ bl_0_120 br_0_120 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c120
+ bl_0_120 br_0_120 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c120
+ bl_0_120 br_0_120 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c120
+ bl_0_120 br_0_120 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c120
+ bl_0_120 br_0_120 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c120
+ bl_0_120 br_0_120 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c120
+ bl_0_120 br_0_120 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c120
+ bl_0_120 br_0_120 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c120
+ bl_0_120 br_0_120 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c120
+ bl_0_120 br_0_120 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c120
+ bl_0_120 br_0_120 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c120
+ bl_0_120 br_0_120 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c120
+ bl_0_120 br_0_120 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c120
+ bl_0_120 br_0_120 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c120
+ bl_0_120 br_0_120 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c120
+ bl_0_120 br_0_120 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c120
+ bl_0_120 br_0_120 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c120
+ bl_0_120 br_0_120 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c120
+ bl_0_120 br_0_120 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c120
+ bl_0_120 br_0_120 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c120
+ bl_0_120 br_0_120 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c120
+ bl_0_120 br_0_120 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c120
+ bl_0_120 br_0_120 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c120
+ bl_0_120 br_0_120 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c120
+ bl_0_120 br_0_120 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c120
+ bl_0_120 br_0_120 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c120
+ bl_0_120 br_0_120 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c120
+ bl_0_120 br_0_120 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c120
+ bl_0_120 br_0_120 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c120
+ bl_0_120 br_0_120 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c120
+ bl_0_120 br_0_120 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c120
+ bl_0_120 br_0_120 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c120
+ bl_0_120 br_0_120 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c120
+ bl_0_120 br_0_120 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c120
+ bl_0_120 br_0_120 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c120
+ bl_0_120 br_0_120 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c120
+ bl_0_120 br_0_120 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c120
+ bl_0_120 br_0_120 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c120
+ bl_0_120 br_0_120 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c120
+ bl_0_120 br_0_120 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c120
+ bl_0_120 br_0_120 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c120
+ bl_0_120 br_0_120 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c121
+ bl_0_121 br_0_121 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c121
+ bl_0_121 br_0_121 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c121
+ bl_0_121 br_0_121 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c121
+ bl_0_121 br_0_121 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c121
+ bl_0_121 br_0_121 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c121
+ bl_0_121 br_0_121 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c121
+ bl_0_121 br_0_121 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c121
+ bl_0_121 br_0_121 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c121
+ bl_0_121 br_0_121 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c121
+ bl_0_121 br_0_121 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c121
+ bl_0_121 br_0_121 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c121
+ bl_0_121 br_0_121 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c121
+ bl_0_121 br_0_121 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c121
+ bl_0_121 br_0_121 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c121
+ bl_0_121 br_0_121 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c121
+ bl_0_121 br_0_121 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c121
+ bl_0_121 br_0_121 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c121
+ bl_0_121 br_0_121 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c121
+ bl_0_121 br_0_121 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c121
+ bl_0_121 br_0_121 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c121
+ bl_0_121 br_0_121 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c121
+ bl_0_121 br_0_121 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c121
+ bl_0_121 br_0_121 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c121
+ bl_0_121 br_0_121 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c121
+ bl_0_121 br_0_121 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c121
+ bl_0_121 br_0_121 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c121
+ bl_0_121 br_0_121 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c121
+ bl_0_121 br_0_121 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c121
+ bl_0_121 br_0_121 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c121
+ bl_0_121 br_0_121 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c121
+ bl_0_121 br_0_121 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c121
+ bl_0_121 br_0_121 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c121
+ bl_0_121 br_0_121 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c121
+ bl_0_121 br_0_121 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c121
+ bl_0_121 br_0_121 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c121
+ bl_0_121 br_0_121 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c121
+ bl_0_121 br_0_121 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c121
+ bl_0_121 br_0_121 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c121
+ bl_0_121 br_0_121 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c121
+ bl_0_121 br_0_121 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c121
+ bl_0_121 br_0_121 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c121
+ bl_0_121 br_0_121 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c121
+ bl_0_121 br_0_121 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c121
+ bl_0_121 br_0_121 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c122
+ bl_0_122 br_0_122 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c122
+ bl_0_122 br_0_122 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c122
+ bl_0_122 br_0_122 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c122
+ bl_0_122 br_0_122 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c122
+ bl_0_122 br_0_122 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c122
+ bl_0_122 br_0_122 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c122
+ bl_0_122 br_0_122 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c122
+ bl_0_122 br_0_122 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c122
+ bl_0_122 br_0_122 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c122
+ bl_0_122 br_0_122 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c122
+ bl_0_122 br_0_122 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c122
+ bl_0_122 br_0_122 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c122
+ bl_0_122 br_0_122 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c122
+ bl_0_122 br_0_122 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c122
+ bl_0_122 br_0_122 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c122
+ bl_0_122 br_0_122 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c122
+ bl_0_122 br_0_122 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c122
+ bl_0_122 br_0_122 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c122
+ bl_0_122 br_0_122 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c122
+ bl_0_122 br_0_122 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c122
+ bl_0_122 br_0_122 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c122
+ bl_0_122 br_0_122 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c122
+ bl_0_122 br_0_122 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c122
+ bl_0_122 br_0_122 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c122
+ bl_0_122 br_0_122 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c122
+ bl_0_122 br_0_122 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c122
+ bl_0_122 br_0_122 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c122
+ bl_0_122 br_0_122 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c122
+ bl_0_122 br_0_122 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c122
+ bl_0_122 br_0_122 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c122
+ bl_0_122 br_0_122 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c122
+ bl_0_122 br_0_122 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c122
+ bl_0_122 br_0_122 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c122
+ bl_0_122 br_0_122 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c122
+ bl_0_122 br_0_122 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c122
+ bl_0_122 br_0_122 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c122
+ bl_0_122 br_0_122 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c122
+ bl_0_122 br_0_122 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c122
+ bl_0_122 br_0_122 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c122
+ bl_0_122 br_0_122 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c122
+ bl_0_122 br_0_122 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c122
+ bl_0_122 br_0_122 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c122
+ bl_0_122 br_0_122 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c122
+ bl_0_122 br_0_122 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c123
+ bl_0_123 br_0_123 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c123
+ bl_0_123 br_0_123 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c123
+ bl_0_123 br_0_123 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c123
+ bl_0_123 br_0_123 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c123
+ bl_0_123 br_0_123 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c123
+ bl_0_123 br_0_123 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c123
+ bl_0_123 br_0_123 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c123
+ bl_0_123 br_0_123 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c123
+ bl_0_123 br_0_123 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c123
+ bl_0_123 br_0_123 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c123
+ bl_0_123 br_0_123 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c123
+ bl_0_123 br_0_123 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c123
+ bl_0_123 br_0_123 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c123
+ bl_0_123 br_0_123 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c123
+ bl_0_123 br_0_123 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c123
+ bl_0_123 br_0_123 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c123
+ bl_0_123 br_0_123 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c123
+ bl_0_123 br_0_123 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c123
+ bl_0_123 br_0_123 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c123
+ bl_0_123 br_0_123 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c123
+ bl_0_123 br_0_123 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c123
+ bl_0_123 br_0_123 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c123
+ bl_0_123 br_0_123 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c123
+ bl_0_123 br_0_123 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c123
+ bl_0_123 br_0_123 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c123
+ bl_0_123 br_0_123 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c123
+ bl_0_123 br_0_123 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c123
+ bl_0_123 br_0_123 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c123
+ bl_0_123 br_0_123 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c123
+ bl_0_123 br_0_123 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c123
+ bl_0_123 br_0_123 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c123
+ bl_0_123 br_0_123 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c123
+ bl_0_123 br_0_123 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c123
+ bl_0_123 br_0_123 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c123
+ bl_0_123 br_0_123 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c123
+ bl_0_123 br_0_123 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c123
+ bl_0_123 br_0_123 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c123
+ bl_0_123 br_0_123 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c123
+ bl_0_123 br_0_123 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c123
+ bl_0_123 br_0_123 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c123
+ bl_0_123 br_0_123 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c123
+ bl_0_123 br_0_123 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c123
+ bl_0_123 br_0_123 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c123
+ bl_0_123 br_0_123 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c124
+ bl_0_124 br_0_124 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c124
+ bl_0_124 br_0_124 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c124
+ bl_0_124 br_0_124 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c124
+ bl_0_124 br_0_124 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c124
+ bl_0_124 br_0_124 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c124
+ bl_0_124 br_0_124 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c124
+ bl_0_124 br_0_124 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c124
+ bl_0_124 br_0_124 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c124
+ bl_0_124 br_0_124 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c124
+ bl_0_124 br_0_124 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c124
+ bl_0_124 br_0_124 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c124
+ bl_0_124 br_0_124 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c124
+ bl_0_124 br_0_124 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c124
+ bl_0_124 br_0_124 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c124
+ bl_0_124 br_0_124 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c124
+ bl_0_124 br_0_124 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c124
+ bl_0_124 br_0_124 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c124
+ bl_0_124 br_0_124 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c124
+ bl_0_124 br_0_124 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c124
+ bl_0_124 br_0_124 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c124
+ bl_0_124 br_0_124 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c124
+ bl_0_124 br_0_124 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c124
+ bl_0_124 br_0_124 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c124
+ bl_0_124 br_0_124 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c124
+ bl_0_124 br_0_124 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c124
+ bl_0_124 br_0_124 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c124
+ bl_0_124 br_0_124 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c124
+ bl_0_124 br_0_124 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c124
+ bl_0_124 br_0_124 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c124
+ bl_0_124 br_0_124 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c124
+ bl_0_124 br_0_124 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c124
+ bl_0_124 br_0_124 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c124
+ bl_0_124 br_0_124 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c124
+ bl_0_124 br_0_124 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c124
+ bl_0_124 br_0_124 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c124
+ bl_0_124 br_0_124 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c124
+ bl_0_124 br_0_124 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c124
+ bl_0_124 br_0_124 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c124
+ bl_0_124 br_0_124 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c124
+ bl_0_124 br_0_124 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c124
+ bl_0_124 br_0_124 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c124
+ bl_0_124 br_0_124 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c124
+ bl_0_124 br_0_124 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c124
+ bl_0_124 br_0_124 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c125
+ bl_0_125 br_0_125 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c125
+ bl_0_125 br_0_125 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c125
+ bl_0_125 br_0_125 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c125
+ bl_0_125 br_0_125 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c125
+ bl_0_125 br_0_125 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c125
+ bl_0_125 br_0_125 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c125
+ bl_0_125 br_0_125 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c125
+ bl_0_125 br_0_125 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c125
+ bl_0_125 br_0_125 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c125
+ bl_0_125 br_0_125 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c125
+ bl_0_125 br_0_125 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c125
+ bl_0_125 br_0_125 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c125
+ bl_0_125 br_0_125 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c125
+ bl_0_125 br_0_125 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c125
+ bl_0_125 br_0_125 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c125
+ bl_0_125 br_0_125 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c125
+ bl_0_125 br_0_125 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c125
+ bl_0_125 br_0_125 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c125
+ bl_0_125 br_0_125 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c125
+ bl_0_125 br_0_125 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c125
+ bl_0_125 br_0_125 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c125
+ bl_0_125 br_0_125 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c125
+ bl_0_125 br_0_125 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c125
+ bl_0_125 br_0_125 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c125
+ bl_0_125 br_0_125 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c125
+ bl_0_125 br_0_125 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c125
+ bl_0_125 br_0_125 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c125
+ bl_0_125 br_0_125 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c125
+ bl_0_125 br_0_125 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c125
+ bl_0_125 br_0_125 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c125
+ bl_0_125 br_0_125 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c125
+ bl_0_125 br_0_125 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c125
+ bl_0_125 br_0_125 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c125
+ bl_0_125 br_0_125 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c125
+ bl_0_125 br_0_125 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c125
+ bl_0_125 br_0_125 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c125
+ bl_0_125 br_0_125 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c125
+ bl_0_125 br_0_125 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c125
+ bl_0_125 br_0_125 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c125
+ bl_0_125 br_0_125 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c125
+ bl_0_125 br_0_125 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c125
+ bl_0_125 br_0_125 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c125
+ bl_0_125 br_0_125 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c125
+ bl_0_125 br_0_125 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c126
+ bl_0_126 br_0_126 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c126
+ bl_0_126 br_0_126 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c126
+ bl_0_126 br_0_126 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c126
+ bl_0_126 br_0_126 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c126
+ bl_0_126 br_0_126 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c126
+ bl_0_126 br_0_126 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c126
+ bl_0_126 br_0_126 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c126
+ bl_0_126 br_0_126 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c126
+ bl_0_126 br_0_126 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c126
+ bl_0_126 br_0_126 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c126
+ bl_0_126 br_0_126 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c126
+ bl_0_126 br_0_126 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c126
+ bl_0_126 br_0_126 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c126
+ bl_0_126 br_0_126 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c126
+ bl_0_126 br_0_126 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c126
+ bl_0_126 br_0_126 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c126
+ bl_0_126 br_0_126 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c126
+ bl_0_126 br_0_126 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c126
+ bl_0_126 br_0_126 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c126
+ bl_0_126 br_0_126 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c126
+ bl_0_126 br_0_126 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c126
+ bl_0_126 br_0_126 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c126
+ bl_0_126 br_0_126 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c126
+ bl_0_126 br_0_126 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c126
+ bl_0_126 br_0_126 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c126
+ bl_0_126 br_0_126 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c126
+ bl_0_126 br_0_126 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c126
+ bl_0_126 br_0_126 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c126
+ bl_0_126 br_0_126 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c126
+ bl_0_126 br_0_126 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c126
+ bl_0_126 br_0_126 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c126
+ bl_0_126 br_0_126 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c126
+ bl_0_126 br_0_126 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c126
+ bl_0_126 br_0_126 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c126
+ bl_0_126 br_0_126 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c126
+ bl_0_126 br_0_126 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c126
+ bl_0_126 br_0_126 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c126
+ bl_0_126 br_0_126 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c126
+ bl_0_126 br_0_126 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c126
+ bl_0_126 br_0_126 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c126
+ bl_0_126 br_0_126 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c126
+ bl_0_126 br_0_126 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c126
+ bl_0_126 br_0_126 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c126
+ bl_0_126 br_0_126 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c127
+ bl_0_127 br_0_127 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c127
+ bl_0_127 br_0_127 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c127
+ bl_0_127 br_0_127 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c127
+ bl_0_127 br_0_127 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c127
+ bl_0_127 br_0_127 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c127
+ bl_0_127 br_0_127 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c127
+ bl_0_127 br_0_127 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c127
+ bl_0_127 br_0_127 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c127
+ bl_0_127 br_0_127 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c127
+ bl_0_127 br_0_127 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c127
+ bl_0_127 br_0_127 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c127
+ bl_0_127 br_0_127 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c127
+ bl_0_127 br_0_127 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c127
+ bl_0_127 br_0_127 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c127
+ bl_0_127 br_0_127 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c127
+ bl_0_127 br_0_127 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c127
+ bl_0_127 br_0_127 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c127
+ bl_0_127 br_0_127 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c127
+ bl_0_127 br_0_127 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c127
+ bl_0_127 br_0_127 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c127
+ bl_0_127 br_0_127 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c127
+ bl_0_127 br_0_127 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c127
+ bl_0_127 br_0_127 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c127
+ bl_0_127 br_0_127 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c127
+ bl_0_127 br_0_127 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c127
+ bl_0_127 br_0_127 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c127
+ bl_0_127 br_0_127 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c127
+ bl_0_127 br_0_127 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c127
+ bl_0_127 br_0_127 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c127
+ bl_0_127 br_0_127 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c127
+ bl_0_127 br_0_127 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c127
+ bl_0_127 br_0_127 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c127
+ bl_0_127 br_0_127 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c127
+ bl_0_127 br_0_127 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c127
+ bl_0_127 br_0_127 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c127
+ bl_0_127 br_0_127 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c127
+ bl_0_127 br_0_127 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c127
+ bl_0_127 br_0_127 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c127
+ bl_0_127 br_0_127 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c127
+ bl_0_127 br_0_127 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c127
+ bl_0_127 br_0_127 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c127
+ bl_0_127 br_0_127 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c127
+ bl_0_127 br_0_127 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c127
+ bl_0_127 br_0_127 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c128
+ bl_0_128 br_0_128 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c128
+ bl_0_128 br_0_128 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c128
+ bl_0_128 br_0_128 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c128
+ bl_0_128 br_0_128 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c128
+ bl_0_128 br_0_128 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c128
+ bl_0_128 br_0_128 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c128
+ bl_0_128 br_0_128 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c128
+ bl_0_128 br_0_128 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c128
+ bl_0_128 br_0_128 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c128
+ bl_0_128 br_0_128 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c128
+ bl_0_128 br_0_128 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c128
+ bl_0_128 br_0_128 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c128
+ bl_0_128 br_0_128 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c128
+ bl_0_128 br_0_128 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c128
+ bl_0_128 br_0_128 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c128
+ bl_0_128 br_0_128 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c128
+ bl_0_128 br_0_128 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c128
+ bl_0_128 br_0_128 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c128
+ bl_0_128 br_0_128 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c128
+ bl_0_128 br_0_128 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c128
+ bl_0_128 br_0_128 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c128
+ bl_0_128 br_0_128 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c128
+ bl_0_128 br_0_128 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c128
+ bl_0_128 br_0_128 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c128
+ bl_0_128 br_0_128 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c128
+ bl_0_128 br_0_128 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c128
+ bl_0_128 br_0_128 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c128
+ bl_0_128 br_0_128 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c128
+ bl_0_128 br_0_128 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c128
+ bl_0_128 br_0_128 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c128
+ bl_0_128 br_0_128 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c128
+ bl_0_128 br_0_128 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c128
+ bl_0_128 br_0_128 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c128
+ bl_0_128 br_0_128 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c128
+ bl_0_128 br_0_128 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c128
+ bl_0_128 br_0_128 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c128
+ bl_0_128 br_0_128 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c128
+ bl_0_128 br_0_128 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c128
+ bl_0_128 br_0_128 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c128
+ bl_0_128 br_0_128 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c128
+ bl_0_128 br_0_128 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c128
+ bl_0_128 br_0_128 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c128
+ bl_0_128 br_0_128 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c128
+ bl_0_128 br_0_128 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c129
+ bl_0_129 br_0_129 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c129
+ bl_0_129 br_0_129 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c129
+ bl_0_129 br_0_129 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c129
+ bl_0_129 br_0_129 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c129
+ bl_0_129 br_0_129 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c129
+ bl_0_129 br_0_129 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c129
+ bl_0_129 br_0_129 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c129
+ bl_0_129 br_0_129 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c129
+ bl_0_129 br_0_129 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c129
+ bl_0_129 br_0_129 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c129
+ bl_0_129 br_0_129 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c129
+ bl_0_129 br_0_129 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c129
+ bl_0_129 br_0_129 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c129
+ bl_0_129 br_0_129 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c129
+ bl_0_129 br_0_129 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c129
+ bl_0_129 br_0_129 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c129
+ bl_0_129 br_0_129 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c129
+ bl_0_129 br_0_129 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c129
+ bl_0_129 br_0_129 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c129
+ bl_0_129 br_0_129 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c129
+ bl_0_129 br_0_129 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c129
+ bl_0_129 br_0_129 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c129
+ bl_0_129 br_0_129 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c129
+ bl_0_129 br_0_129 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c129
+ bl_0_129 br_0_129 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c129
+ bl_0_129 br_0_129 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c129
+ bl_0_129 br_0_129 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c129
+ bl_0_129 br_0_129 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c129
+ bl_0_129 br_0_129 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c129
+ bl_0_129 br_0_129 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c129
+ bl_0_129 br_0_129 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c129
+ bl_0_129 br_0_129 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c129
+ bl_0_129 br_0_129 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c129
+ bl_0_129 br_0_129 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c129
+ bl_0_129 br_0_129 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c129
+ bl_0_129 br_0_129 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c129
+ bl_0_129 br_0_129 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c129
+ bl_0_129 br_0_129 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c129
+ bl_0_129 br_0_129 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c129
+ bl_0_129 br_0_129 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c129
+ bl_0_129 br_0_129 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c129
+ bl_0_129 br_0_129 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c129
+ bl_0_129 br_0_129 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c129
+ bl_0_129 br_0_129 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c130
+ bl_0_130 br_0_130 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c130
+ bl_0_130 br_0_130 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c130
+ bl_0_130 br_0_130 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c130
+ bl_0_130 br_0_130 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c130
+ bl_0_130 br_0_130 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c130
+ bl_0_130 br_0_130 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c130
+ bl_0_130 br_0_130 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c130
+ bl_0_130 br_0_130 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c130
+ bl_0_130 br_0_130 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c130
+ bl_0_130 br_0_130 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c130
+ bl_0_130 br_0_130 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c130
+ bl_0_130 br_0_130 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c130
+ bl_0_130 br_0_130 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c130
+ bl_0_130 br_0_130 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c130
+ bl_0_130 br_0_130 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c130
+ bl_0_130 br_0_130 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c130
+ bl_0_130 br_0_130 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c130
+ bl_0_130 br_0_130 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c130
+ bl_0_130 br_0_130 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c130
+ bl_0_130 br_0_130 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c130
+ bl_0_130 br_0_130 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c130
+ bl_0_130 br_0_130 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c130
+ bl_0_130 br_0_130 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c130
+ bl_0_130 br_0_130 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c130
+ bl_0_130 br_0_130 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c130
+ bl_0_130 br_0_130 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c130
+ bl_0_130 br_0_130 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c130
+ bl_0_130 br_0_130 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c130
+ bl_0_130 br_0_130 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c130
+ bl_0_130 br_0_130 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c130
+ bl_0_130 br_0_130 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c130
+ bl_0_130 br_0_130 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c130
+ bl_0_130 br_0_130 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c130
+ bl_0_130 br_0_130 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c130
+ bl_0_130 br_0_130 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c130
+ bl_0_130 br_0_130 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c130
+ bl_0_130 br_0_130 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c130
+ bl_0_130 br_0_130 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c130
+ bl_0_130 br_0_130 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c130
+ bl_0_130 br_0_130 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c130
+ bl_0_130 br_0_130 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c130
+ bl_0_130 br_0_130 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c130
+ bl_0_130 br_0_130 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c130
+ bl_0_130 br_0_130 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c131
+ bl_0_131 br_0_131 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c131
+ bl_0_131 br_0_131 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c131
+ bl_0_131 br_0_131 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c131
+ bl_0_131 br_0_131 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c131
+ bl_0_131 br_0_131 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c131
+ bl_0_131 br_0_131 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c131
+ bl_0_131 br_0_131 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c131
+ bl_0_131 br_0_131 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c131
+ bl_0_131 br_0_131 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c131
+ bl_0_131 br_0_131 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c131
+ bl_0_131 br_0_131 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c131
+ bl_0_131 br_0_131 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c131
+ bl_0_131 br_0_131 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c131
+ bl_0_131 br_0_131 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c131
+ bl_0_131 br_0_131 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c131
+ bl_0_131 br_0_131 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c131
+ bl_0_131 br_0_131 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c131
+ bl_0_131 br_0_131 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c131
+ bl_0_131 br_0_131 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c131
+ bl_0_131 br_0_131 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c131
+ bl_0_131 br_0_131 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c131
+ bl_0_131 br_0_131 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c131
+ bl_0_131 br_0_131 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c131
+ bl_0_131 br_0_131 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c131
+ bl_0_131 br_0_131 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c131
+ bl_0_131 br_0_131 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c131
+ bl_0_131 br_0_131 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c131
+ bl_0_131 br_0_131 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c131
+ bl_0_131 br_0_131 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c131
+ bl_0_131 br_0_131 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c131
+ bl_0_131 br_0_131 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c131
+ bl_0_131 br_0_131 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c131
+ bl_0_131 br_0_131 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c131
+ bl_0_131 br_0_131 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c131
+ bl_0_131 br_0_131 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c131
+ bl_0_131 br_0_131 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c131
+ bl_0_131 br_0_131 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c131
+ bl_0_131 br_0_131 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c131
+ bl_0_131 br_0_131 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c131
+ bl_0_131 br_0_131 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c131
+ bl_0_131 br_0_131 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c131
+ bl_0_131 br_0_131 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c131
+ bl_0_131 br_0_131 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c131
+ bl_0_131 br_0_131 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c132
+ bl_0_132 br_0_132 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c132
+ bl_0_132 br_0_132 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c132
+ bl_0_132 br_0_132 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c132
+ bl_0_132 br_0_132 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c132
+ bl_0_132 br_0_132 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c132
+ bl_0_132 br_0_132 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c132
+ bl_0_132 br_0_132 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c132
+ bl_0_132 br_0_132 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c132
+ bl_0_132 br_0_132 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c132
+ bl_0_132 br_0_132 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c132
+ bl_0_132 br_0_132 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c132
+ bl_0_132 br_0_132 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c132
+ bl_0_132 br_0_132 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c132
+ bl_0_132 br_0_132 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c132
+ bl_0_132 br_0_132 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c132
+ bl_0_132 br_0_132 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c132
+ bl_0_132 br_0_132 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c132
+ bl_0_132 br_0_132 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c132
+ bl_0_132 br_0_132 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c132
+ bl_0_132 br_0_132 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c132
+ bl_0_132 br_0_132 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c132
+ bl_0_132 br_0_132 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c132
+ bl_0_132 br_0_132 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c132
+ bl_0_132 br_0_132 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c132
+ bl_0_132 br_0_132 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c132
+ bl_0_132 br_0_132 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c132
+ bl_0_132 br_0_132 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c132
+ bl_0_132 br_0_132 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c132
+ bl_0_132 br_0_132 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c132
+ bl_0_132 br_0_132 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c132
+ bl_0_132 br_0_132 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c132
+ bl_0_132 br_0_132 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c132
+ bl_0_132 br_0_132 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c132
+ bl_0_132 br_0_132 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c132
+ bl_0_132 br_0_132 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c132
+ bl_0_132 br_0_132 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c132
+ bl_0_132 br_0_132 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c132
+ bl_0_132 br_0_132 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c132
+ bl_0_132 br_0_132 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c132
+ bl_0_132 br_0_132 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c132
+ bl_0_132 br_0_132 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c132
+ bl_0_132 br_0_132 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c132
+ bl_0_132 br_0_132 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c132
+ bl_0_132 br_0_132 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c133
+ bl_0_133 br_0_133 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c133
+ bl_0_133 br_0_133 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c133
+ bl_0_133 br_0_133 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c133
+ bl_0_133 br_0_133 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c133
+ bl_0_133 br_0_133 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c133
+ bl_0_133 br_0_133 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c133
+ bl_0_133 br_0_133 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c133
+ bl_0_133 br_0_133 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c133
+ bl_0_133 br_0_133 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c133
+ bl_0_133 br_0_133 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c133
+ bl_0_133 br_0_133 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c133
+ bl_0_133 br_0_133 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c133
+ bl_0_133 br_0_133 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c133
+ bl_0_133 br_0_133 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c133
+ bl_0_133 br_0_133 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c133
+ bl_0_133 br_0_133 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c133
+ bl_0_133 br_0_133 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c133
+ bl_0_133 br_0_133 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c133
+ bl_0_133 br_0_133 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c133
+ bl_0_133 br_0_133 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c133
+ bl_0_133 br_0_133 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c133
+ bl_0_133 br_0_133 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c133
+ bl_0_133 br_0_133 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c133
+ bl_0_133 br_0_133 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c133
+ bl_0_133 br_0_133 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c133
+ bl_0_133 br_0_133 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c133
+ bl_0_133 br_0_133 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c133
+ bl_0_133 br_0_133 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c133
+ bl_0_133 br_0_133 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c133
+ bl_0_133 br_0_133 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c133
+ bl_0_133 br_0_133 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c133
+ bl_0_133 br_0_133 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c133
+ bl_0_133 br_0_133 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c133
+ bl_0_133 br_0_133 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c133
+ bl_0_133 br_0_133 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c133
+ bl_0_133 br_0_133 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c133
+ bl_0_133 br_0_133 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c133
+ bl_0_133 br_0_133 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c133
+ bl_0_133 br_0_133 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c133
+ bl_0_133 br_0_133 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c133
+ bl_0_133 br_0_133 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c133
+ bl_0_133 br_0_133 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c133
+ bl_0_133 br_0_133 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c133
+ bl_0_133 br_0_133 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c134
+ bl_0_134 br_0_134 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c134
+ bl_0_134 br_0_134 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c134
+ bl_0_134 br_0_134 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c134
+ bl_0_134 br_0_134 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c134
+ bl_0_134 br_0_134 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c134
+ bl_0_134 br_0_134 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c134
+ bl_0_134 br_0_134 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c134
+ bl_0_134 br_0_134 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c134
+ bl_0_134 br_0_134 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c134
+ bl_0_134 br_0_134 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c134
+ bl_0_134 br_0_134 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c134
+ bl_0_134 br_0_134 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c134
+ bl_0_134 br_0_134 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c134
+ bl_0_134 br_0_134 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c134
+ bl_0_134 br_0_134 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c134
+ bl_0_134 br_0_134 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c134
+ bl_0_134 br_0_134 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c134
+ bl_0_134 br_0_134 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c134
+ bl_0_134 br_0_134 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c134
+ bl_0_134 br_0_134 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c134
+ bl_0_134 br_0_134 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c134
+ bl_0_134 br_0_134 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c134
+ bl_0_134 br_0_134 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c134
+ bl_0_134 br_0_134 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c134
+ bl_0_134 br_0_134 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c134
+ bl_0_134 br_0_134 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c134
+ bl_0_134 br_0_134 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c134
+ bl_0_134 br_0_134 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c134
+ bl_0_134 br_0_134 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c134
+ bl_0_134 br_0_134 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c134
+ bl_0_134 br_0_134 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c134
+ bl_0_134 br_0_134 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c134
+ bl_0_134 br_0_134 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c134
+ bl_0_134 br_0_134 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c134
+ bl_0_134 br_0_134 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c134
+ bl_0_134 br_0_134 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c134
+ bl_0_134 br_0_134 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c134
+ bl_0_134 br_0_134 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c134
+ bl_0_134 br_0_134 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c134
+ bl_0_134 br_0_134 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c134
+ bl_0_134 br_0_134 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c134
+ bl_0_134 br_0_134 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c134
+ bl_0_134 br_0_134 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c134
+ bl_0_134 br_0_134 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c135
+ bl_0_135 br_0_135 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c135
+ bl_0_135 br_0_135 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c135
+ bl_0_135 br_0_135 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c135
+ bl_0_135 br_0_135 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c135
+ bl_0_135 br_0_135 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c135
+ bl_0_135 br_0_135 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c135
+ bl_0_135 br_0_135 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c135
+ bl_0_135 br_0_135 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c135
+ bl_0_135 br_0_135 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c135
+ bl_0_135 br_0_135 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c135
+ bl_0_135 br_0_135 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c135
+ bl_0_135 br_0_135 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c135
+ bl_0_135 br_0_135 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c135
+ bl_0_135 br_0_135 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c135
+ bl_0_135 br_0_135 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c135
+ bl_0_135 br_0_135 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c135
+ bl_0_135 br_0_135 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c135
+ bl_0_135 br_0_135 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c135
+ bl_0_135 br_0_135 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c135
+ bl_0_135 br_0_135 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c135
+ bl_0_135 br_0_135 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c135
+ bl_0_135 br_0_135 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c135
+ bl_0_135 br_0_135 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c135
+ bl_0_135 br_0_135 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c135
+ bl_0_135 br_0_135 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c135
+ bl_0_135 br_0_135 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c135
+ bl_0_135 br_0_135 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c135
+ bl_0_135 br_0_135 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c135
+ bl_0_135 br_0_135 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c135
+ bl_0_135 br_0_135 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c135
+ bl_0_135 br_0_135 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c135
+ bl_0_135 br_0_135 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c135
+ bl_0_135 br_0_135 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c135
+ bl_0_135 br_0_135 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c135
+ bl_0_135 br_0_135 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c135
+ bl_0_135 br_0_135 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c135
+ bl_0_135 br_0_135 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c135
+ bl_0_135 br_0_135 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c135
+ bl_0_135 br_0_135 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c135
+ bl_0_135 br_0_135 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c135
+ bl_0_135 br_0_135 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c135
+ bl_0_135 br_0_135 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c135
+ bl_0_135 br_0_135 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c135
+ bl_0_135 br_0_135 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c136
+ bl_0_136 br_0_136 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c136
+ bl_0_136 br_0_136 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c136
+ bl_0_136 br_0_136 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c136
+ bl_0_136 br_0_136 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c136
+ bl_0_136 br_0_136 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c136
+ bl_0_136 br_0_136 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c136
+ bl_0_136 br_0_136 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c136
+ bl_0_136 br_0_136 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c136
+ bl_0_136 br_0_136 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c136
+ bl_0_136 br_0_136 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c136
+ bl_0_136 br_0_136 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c136
+ bl_0_136 br_0_136 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c136
+ bl_0_136 br_0_136 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c136
+ bl_0_136 br_0_136 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c136
+ bl_0_136 br_0_136 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c136
+ bl_0_136 br_0_136 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c136
+ bl_0_136 br_0_136 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c136
+ bl_0_136 br_0_136 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c136
+ bl_0_136 br_0_136 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c136
+ bl_0_136 br_0_136 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c136
+ bl_0_136 br_0_136 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c136
+ bl_0_136 br_0_136 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c136
+ bl_0_136 br_0_136 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c136
+ bl_0_136 br_0_136 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c136
+ bl_0_136 br_0_136 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c136
+ bl_0_136 br_0_136 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c136
+ bl_0_136 br_0_136 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c136
+ bl_0_136 br_0_136 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c136
+ bl_0_136 br_0_136 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c136
+ bl_0_136 br_0_136 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c136
+ bl_0_136 br_0_136 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c136
+ bl_0_136 br_0_136 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c136
+ bl_0_136 br_0_136 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c136
+ bl_0_136 br_0_136 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c136
+ bl_0_136 br_0_136 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c136
+ bl_0_136 br_0_136 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c136
+ bl_0_136 br_0_136 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c136
+ bl_0_136 br_0_136 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c136
+ bl_0_136 br_0_136 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c136
+ bl_0_136 br_0_136 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c136
+ bl_0_136 br_0_136 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c136
+ bl_0_136 br_0_136 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c136
+ bl_0_136 br_0_136 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c136
+ bl_0_136 br_0_136 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c137
+ bl_0_137 br_0_137 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c137
+ bl_0_137 br_0_137 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c137
+ bl_0_137 br_0_137 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c137
+ bl_0_137 br_0_137 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c137
+ bl_0_137 br_0_137 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c137
+ bl_0_137 br_0_137 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c137
+ bl_0_137 br_0_137 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c137
+ bl_0_137 br_0_137 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c137
+ bl_0_137 br_0_137 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c137
+ bl_0_137 br_0_137 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c137
+ bl_0_137 br_0_137 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c137
+ bl_0_137 br_0_137 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c137
+ bl_0_137 br_0_137 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c137
+ bl_0_137 br_0_137 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c137
+ bl_0_137 br_0_137 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c137
+ bl_0_137 br_0_137 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c137
+ bl_0_137 br_0_137 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c137
+ bl_0_137 br_0_137 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c137
+ bl_0_137 br_0_137 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c137
+ bl_0_137 br_0_137 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c137
+ bl_0_137 br_0_137 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c137
+ bl_0_137 br_0_137 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c137
+ bl_0_137 br_0_137 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c137
+ bl_0_137 br_0_137 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c137
+ bl_0_137 br_0_137 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c137
+ bl_0_137 br_0_137 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c137
+ bl_0_137 br_0_137 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c137
+ bl_0_137 br_0_137 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c137
+ bl_0_137 br_0_137 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c137
+ bl_0_137 br_0_137 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c137
+ bl_0_137 br_0_137 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c137
+ bl_0_137 br_0_137 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c137
+ bl_0_137 br_0_137 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c137
+ bl_0_137 br_0_137 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c137
+ bl_0_137 br_0_137 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c137
+ bl_0_137 br_0_137 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c137
+ bl_0_137 br_0_137 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c137
+ bl_0_137 br_0_137 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c137
+ bl_0_137 br_0_137 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c137
+ bl_0_137 br_0_137 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c137
+ bl_0_137 br_0_137 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c137
+ bl_0_137 br_0_137 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c137
+ bl_0_137 br_0_137 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c137
+ bl_0_137 br_0_137 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c138
+ bl_0_138 br_0_138 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c138
+ bl_0_138 br_0_138 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c138
+ bl_0_138 br_0_138 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c138
+ bl_0_138 br_0_138 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c138
+ bl_0_138 br_0_138 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c138
+ bl_0_138 br_0_138 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c138
+ bl_0_138 br_0_138 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c138
+ bl_0_138 br_0_138 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c138
+ bl_0_138 br_0_138 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c138
+ bl_0_138 br_0_138 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c138
+ bl_0_138 br_0_138 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c138
+ bl_0_138 br_0_138 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c138
+ bl_0_138 br_0_138 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c138
+ bl_0_138 br_0_138 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c138
+ bl_0_138 br_0_138 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c138
+ bl_0_138 br_0_138 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c138
+ bl_0_138 br_0_138 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c138
+ bl_0_138 br_0_138 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c138
+ bl_0_138 br_0_138 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c138
+ bl_0_138 br_0_138 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c138
+ bl_0_138 br_0_138 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c138
+ bl_0_138 br_0_138 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c138
+ bl_0_138 br_0_138 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c138
+ bl_0_138 br_0_138 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c138
+ bl_0_138 br_0_138 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c138
+ bl_0_138 br_0_138 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c138
+ bl_0_138 br_0_138 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c138
+ bl_0_138 br_0_138 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c138
+ bl_0_138 br_0_138 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c138
+ bl_0_138 br_0_138 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c138
+ bl_0_138 br_0_138 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c138
+ bl_0_138 br_0_138 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c138
+ bl_0_138 br_0_138 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c138
+ bl_0_138 br_0_138 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c138
+ bl_0_138 br_0_138 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c138
+ bl_0_138 br_0_138 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c138
+ bl_0_138 br_0_138 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c138
+ bl_0_138 br_0_138 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c138
+ bl_0_138 br_0_138 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c138
+ bl_0_138 br_0_138 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c138
+ bl_0_138 br_0_138 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c138
+ bl_0_138 br_0_138 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c138
+ bl_0_138 br_0_138 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c138
+ bl_0_138 br_0_138 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c139
+ bl_0_139 br_0_139 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c139
+ bl_0_139 br_0_139 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c139
+ bl_0_139 br_0_139 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c139
+ bl_0_139 br_0_139 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c139
+ bl_0_139 br_0_139 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c139
+ bl_0_139 br_0_139 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c139
+ bl_0_139 br_0_139 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c139
+ bl_0_139 br_0_139 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c139
+ bl_0_139 br_0_139 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c139
+ bl_0_139 br_0_139 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c139
+ bl_0_139 br_0_139 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c139
+ bl_0_139 br_0_139 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c139
+ bl_0_139 br_0_139 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c139
+ bl_0_139 br_0_139 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c139
+ bl_0_139 br_0_139 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c139
+ bl_0_139 br_0_139 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c139
+ bl_0_139 br_0_139 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c139
+ bl_0_139 br_0_139 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c139
+ bl_0_139 br_0_139 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c139
+ bl_0_139 br_0_139 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c139
+ bl_0_139 br_0_139 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c139
+ bl_0_139 br_0_139 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c139
+ bl_0_139 br_0_139 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c139
+ bl_0_139 br_0_139 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c139
+ bl_0_139 br_0_139 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c139
+ bl_0_139 br_0_139 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c139
+ bl_0_139 br_0_139 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c139
+ bl_0_139 br_0_139 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c139
+ bl_0_139 br_0_139 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c139
+ bl_0_139 br_0_139 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c139
+ bl_0_139 br_0_139 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c139
+ bl_0_139 br_0_139 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c139
+ bl_0_139 br_0_139 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c139
+ bl_0_139 br_0_139 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c139
+ bl_0_139 br_0_139 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c139
+ bl_0_139 br_0_139 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c139
+ bl_0_139 br_0_139 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c139
+ bl_0_139 br_0_139 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c139
+ bl_0_139 br_0_139 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c139
+ bl_0_139 br_0_139 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c139
+ bl_0_139 br_0_139 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c139
+ bl_0_139 br_0_139 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c139
+ bl_0_139 br_0_139 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c139
+ bl_0_139 br_0_139 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c140
+ bl_0_140 br_0_140 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c140
+ bl_0_140 br_0_140 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c140
+ bl_0_140 br_0_140 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c140
+ bl_0_140 br_0_140 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c140
+ bl_0_140 br_0_140 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c140
+ bl_0_140 br_0_140 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c140
+ bl_0_140 br_0_140 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c140
+ bl_0_140 br_0_140 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c140
+ bl_0_140 br_0_140 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c140
+ bl_0_140 br_0_140 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c140
+ bl_0_140 br_0_140 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c140
+ bl_0_140 br_0_140 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c140
+ bl_0_140 br_0_140 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c140
+ bl_0_140 br_0_140 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c140
+ bl_0_140 br_0_140 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c140
+ bl_0_140 br_0_140 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c140
+ bl_0_140 br_0_140 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c140
+ bl_0_140 br_0_140 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c140
+ bl_0_140 br_0_140 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c140
+ bl_0_140 br_0_140 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c140
+ bl_0_140 br_0_140 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c140
+ bl_0_140 br_0_140 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c140
+ bl_0_140 br_0_140 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c140
+ bl_0_140 br_0_140 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c140
+ bl_0_140 br_0_140 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c140
+ bl_0_140 br_0_140 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c140
+ bl_0_140 br_0_140 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c140
+ bl_0_140 br_0_140 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c140
+ bl_0_140 br_0_140 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c140
+ bl_0_140 br_0_140 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c140
+ bl_0_140 br_0_140 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c140
+ bl_0_140 br_0_140 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c140
+ bl_0_140 br_0_140 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c140
+ bl_0_140 br_0_140 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c140
+ bl_0_140 br_0_140 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c140
+ bl_0_140 br_0_140 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c140
+ bl_0_140 br_0_140 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c140
+ bl_0_140 br_0_140 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c140
+ bl_0_140 br_0_140 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c140
+ bl_0_140 br_0_140 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c140
+ bl_0_140 br_0_140 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c140
+ bl_0_140 br_0_140 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c140
+ bl_0_140 br_0_140 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c140
+ bl_0_140 br_0_140 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c141
+ bl_0_141 br_0_141 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c141
+ bl_0_141 br_0_141 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c141
+ bl_0_141 br_0_141 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c141
+ bl_0_141 br_0_141 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c141
+ bl_0_141 br_0_141 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c141
+ bl_0_141 br_0_141 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c141
+ bl_0_141 br_0_141 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c141
+ bl_0_141 br_0_141 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c141
+ bl_0_141 br_0_141 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c141
+ bl_0_141 br_0_141 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c141
+ bl_0_141 br_0_141 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c141
+ bl_0_141 br_0_141 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c141
+ bl_0_141 br_0_141 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c141
+ bl_0_141 br_0_141 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c141
+ bl_0_141 br_0_141 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c141
+ bl_0_141 br_0_141 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c141
+ bl_0_141 br_0_141 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c141
+ bl_0_141 br_0_141 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c141
+ bl_0_141 br_0_141 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c141
+ bl_0_141 br_0_141 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c141
+ bl_0_141 br_0_141 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c141
+ bl_0_141 br_0_141 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c141
+ bl_0_141 br_0_141 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c141
+ bl_0_141 br_0_141 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c141
+ bl_0_141 br_0_141 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c141
+ bl_0_141 br_0_141 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c141
+ bl_0_141 br_0_141 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c141
+ bl_0_141 br_0_141 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c141
+ bl_0_141 br_0_141 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c141
+ bl_0_141 br_0_141 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c141
+ bl_0_141 br_0_141 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c141
+ bl_0_141 br_0_141 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c141
+ bl_0_141 br_0_141 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c141
+ bl_0_141 br_0_141 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c141
+ bl_0_141 br_0_141 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c141
+ bl_0_141 br_0_141 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c141
+ bl_0_141 br_0_141 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c141
+ bl_0_141 br_0_141 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c141
+ bl_0_141 br_0_141 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c141
+ bl_0_141 br_0_141 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c141
+ bl_0_141 br_0_141 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c141
+ bl_0_141 br_0_141 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c141
+ bl_0_141 br_0_141 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c141
+ bl_0_141 br_0_141 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c142
+ bl_0_142 br_0_142 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c142
+ bl_0_142 br_0_142 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c142
+ bl_0_142 br_0_142 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c142
+ bl_0_142 br_0_142 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c142
+ bl_0_142 br_0_142 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c142
+ bl_0_142 br_0_142 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c142
+ bl_0_142 br_0_142 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c142
+ bl_0_142 br_0_142 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c142
+ bl_0_142 br_0_142 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c142
+ bl_0_142 br_0_142 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c142
+ bl_0_142 br_0_142 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c142
+ bl_0_142 br_0_142 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c142
+ bl_0_142 br_0_142 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c142
+ bl_0_142 br_0_142 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c142
+ bl_0_142 br_0_142 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c142
+ bl_0_142 br_0_142 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c142
+ bl_0_142 br_0_142 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c142
+ bl_0_142 br_0_142 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c142
+ bl_0_142 br_0_142 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c142
+ bl_0_142 br_0_142 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c142
+ bl_0_142 br_0_142 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c142
+ bl_0_142 br_0_142 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c142
+ bl_0_142 br_0_142 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c142
+ bl_0_142 br_0_142 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c142
+ bl_0_142 br_0_142 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c142
+ bl_0_142 br_0_142 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c142
+ bl_0_142 br_0_142 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c142
+ bl_0_142 br_0_142 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c142
+ bl_0_142 br_0_142 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c142
+ bl_0_142 br_0_142 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c142
+ bl_0_142 br_0_142 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c142
+ bl_0_142 br_0_142 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c142
+ bl_0_142 br_0_142 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c142
+ bl_0_142 br_0_142 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c142
+ bl_0_142 br_0_142 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c142
+ bl_0_142 br_0_142 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c142
+ bl_0_142 br_0_142 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c142
+ bl_0_142 br_0_142 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c142
+ bl_0_142 br_0_142 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c142
+ bl_0_142 br_0_142 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c142
+ bl_0_142 br_0_142 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c142
+ bl_0_142 br_0_142 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c142
+ bl_0_142 br_0_142 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c142
+ bl_0_142 br_0_142 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c143
+ bl_0_143 br_0_143 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c143
+ bl_0_143 br_0_143 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c143
+ bl_0_143 br_0_143 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c143
+ bl_0_143 br_0_143 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c143
+ bl_0_143 br_0_143 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c143
+ bl_0_143 br_0_143 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c143
+ bl_0_143 br_0_143 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c143
+ bl_0_143 br_0_143 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c143
+ bl_0_143 br_0_143 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c143
+ bl_0_143 br_0_143 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c143
+ bl_0_143 br_0_143 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c143
+ bl_0_143 br_0_143 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c143
+ bl_0_143 br_0_143 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c143
+ bl_0_143 br_0_143 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c143
+ bl_0_143 br_0_143 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c143
+ bl_0_143 br_0_143 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c143
+ bl_0_143 br_0_143 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c143
+ bl_0_143 br_0_143 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c143
+ bl_0_143 br_0_143 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c143
+ bl_0_143 br_0_143 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c143
+ bl_0_143 br_0_143 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c143
+ bl_0_143 br_0_143 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c143
+ bl_0_143 br_0_143 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c143
+ bl_0_143 br_0_143 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c143
+ bl_0_143 br_0_143 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c143
+ bl_0_143 br_0_143 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c143
+ bl_0_143 br_0_143 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c143
+ bl_0_143 br_0_143 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c143
+ bl_0_143 br_0_143 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c143
+ bl_0_143 br_0_143 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c143
+ bl_0_143 br_0_143 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c143
+ bl_0_143 br_0_143 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c143
+ bl_0_143 br_0_143 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c143
+ bl_0_143 br_0_143 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c143
+ bl_0_143 br_0_143 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c143
+ bl_0_143 br_0_143 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c143
+ bl_0_143 br_0_143 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c143
+ bl_0_143 br_0_143 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c143
+ bl_0_143 br_0_143 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c143
+ bl_0_143 br_0_143 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c143
+ bl_0_143 br_0_143 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c143
+ bl_0_143 br_0_143 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c143
+ bl_0_143 br_0_143 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c143
+ bl_0_143 br_0_143 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c144
+ bl_0_144 br_0_144 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c144
+ bl_0_144 br_0_144 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c144
+ bl_0_144 br_0_144 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c144
+ bl_0_144 br_0_144 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c144
+ bl_0_144 br_0_144 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c144
+ bl_0_144 br_0_144 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c144
+ bl_0_144 br_0_144 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c144
+ bl_0_144 br_0_144 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c144
+ bl_0_144 br_0_144 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c144
+ bl_0_144 br_0_144 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c144
+ bl_0_144 br_0_144 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c144
+ bl_0_144 br_0_144 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c144
+ bl_0_144 br_0_144 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c144
+ bl_0_144 br_0_144 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c144
+ bl_0_144 br_0_144 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c144
+ bl_0_144 br_0_144 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c144
+ bl_0_144 br_0_144 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c144
+ bl_0_144 br_0_144 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c144
+ bl_0_144 br_0_144 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c144
+ bl_0_144 br_0_144 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c144
+ bl_0_144 br_0_144 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c144
+ bl_0_144 br_0_144 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c144
+ bl_0_144 br_0_144 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c144
+ bl_0_144 br_0_144 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c144
+ bl_0_144 br_0_144 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c144
+ bl_0_144 br_0_144 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c144
+ bl_0_144 br_0_144 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c144
+ bl_0_144 br_0_144 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c144
+ bl_0_144 br_0_144 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c144
+ bl_0_144 br_0_144 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c144
+ bl_0_144 br_0_144 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c144
+ bl_0_144 br_0_144 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c144
+ bl_0_144 br_0_144 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c144
+ bl_0_144 br_0_144 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c144
+ bl_0_144 br_0_144 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c144
+ bl_0_144 br_0_144 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c144
+ bl_0_144 br_0_144 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c144
+ bl_0_144 br_0_144 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c144
+ bl_0_144 br_0_144 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c144
+ bl_0_144 br_0_144 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c144
+ bl_0_144 br_0_144 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c144
+ bl_0_144 br_0_144 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c144
+ bl_0_144 br_0_144 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c144
+ bl_0_144 br_0_144 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c145
+ bl_0_145 br_0_145 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c145
+ bl_0_145 br_0_145 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c145
+ bl_0_145 br_0_145 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c145
+ bl_0_145 br_0_145 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c145
+ bl_0_145 br_0_145 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c145
+ bl_0_145 br_0_145 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c145
+ bl_0_145 br_0_145 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c145
+ bl_0_145 br_0_145 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c145
+ bl_0_145 br_0_145 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c145
+ bl_0_145 br_0_145 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c145
+ bl_0_145 br_0_145 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c145
+ bl_0_145 br_0_145 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c145
+ bl_0_145 br_0_145 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c145
+ bl_0_145 br_0_145 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c145
+ bl_0_145 br_0_145 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c145
+ bl_0_145 br_0_145 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c145
+ bl_0_145 br_0_145 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c145
+ bl_0_145 br_0_145 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c145
+ bl_0_145 br_0_145 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c145
+ bl_0_145 br_0_145 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c145
+ bl_0_145 br_0_145 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c145
+ bl_0_145 br_0_145 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c145
+ bl_0_145 br_0_145 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c145
+ bl_0_145 br_0_145 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c145
+ bl_0_145 br_0_145 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c145
+ bl_0_145 br_0_145 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c145
+ bl_0_145 br_0_145 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c145
+ bl_0_145 br_0_145 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c145
+ bl_0_145 br_0_145 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c145
+ bl_0_145 br_0_145 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c145
+ bl_0_145 br_0_145 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c145
+ bl_0_145 br_0_145 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c145
+ bl_0_145 br_0_145 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c145
+ bl_0_145 br_0_145 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c145
+ bl_0_145 br_0_145 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c145
+ bl_0_145 br_0_145 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c145
+ bl_0_145 br_0_145 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c145
+ bl_0_145 br_0_145 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c145
+ bl_0_145 br_0_145 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c145
+ bl_0_145 br_0_145 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c145
+ bl_0_145 br_0_145 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c145
+ bl_0_145 br_0_145 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c145
+ bl_0_145 br_0_145 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c145
+ bl_0_145 br_0_145 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c146
+ bl_0_146 br_0_146 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c146
+ bl_0_146 br_0_146 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c146
+ bl_0_146 br_0_146 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c146
+ bl_0_146 br_0_146 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c146
+ bl_0_146 br_0_146 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c146
+ bl_0_146 br_0_146 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c146
+ bl_0_146 br_0_146 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c146
+ bl_0_146 br_0_146 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c146
+ bl_0_146 br_0_146 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c146
+ bl_0_146 br_0_146 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c146
+ bl_0_146 br_0_146 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c146
+ bl_0_146 br_0_146 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c146
+ bl_0_146 br_0_146 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c146
+ bl_0_146 br_0_146 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c146
+ bl_0_146 br_0_146 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c146
+ bl_0_146 br_0_146 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c146
+ bl_0_146 br_0_146 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c146
+ bl_0_146 br_0_146 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c146
+ bl_0_146 br_0_146 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c146
+ bl_0_146 br_0_146 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c146
+ bl_0_146 br_0_146 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c146
+ bl_0_146 br_0_146 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c146
+ bl_0_146 br_0_146 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c146
+ bl_0_146 br_0_146 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c146
+ bl_0_146 br_0_146 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c146
+ bl_0_146 br_0_146 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c146
+ bl_0_146 br_0_146 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c146
+ bl_0_146 br_0_146 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c146
+ bl_0_146 br_0_146 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c146
+ bl_0_146 br_0_146 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c146
+ bl_0_146 br_0_146 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c146
+ bl_0_146 br_0_146 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c146
+ bl_0_146 br_0_146 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c146
+ bl_0_146 br_0_146 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c146
+ bl_0_146 br_0_146 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c146
+ bl_0_146 br_0_146 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c146
+ bl_0_146 br_0_146 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c146
+ bl_0_146 br_0_146 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c146
+ bl_0_146 br_0_146 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c146
+ bl_0_146 br_0_146 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c146
+ bl_0_146 br_0_146 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c146
+ bl_0_146 br_0_146 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c146
+ bl_0_146 br_0_146 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c146
+ bl_0_146 br_0_146 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c147
+ bl_0_147 br_0_147 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c147
+ bl_0_147 br_0_147 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c147
+ bl_0_147 br_0_147 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c147
+ bl_0_147 br_0_147 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c147
+ bl_0_147 br_0_147 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c147
+ bl_0_147 br_0_147 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c147
+ bl_0_147 br_0_147 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c147
+ bl_0_147 br_0_147 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c147
+ bl_0_147 br_0_147 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c147
+ bl_0_147 br_0_147 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c147
+ bl_0_147 br_0_147 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c147
+ bl_0_147 br_0_147 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c147
+ bl_0_147 br_0_147 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c147
+ bl_0_147 br_0_147 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c147
+ bl_0_147 br_0_147 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c147
+ bl_0_147 br_0_147 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c147
+ bl_0_147 br_0_147 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c147
+ bl_0_147 br_0_147 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c147
+ bl_0_147 br_0_147 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c147
+ bl_0_147 br_0_147 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c147
+ bl_0_147 br_0_147 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c147
+ bl_0_147 br_0_147 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c147
+ bl_0_147 br_0_147 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c147
+ bl_0_147 br_0_147 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c147
+ bl_0_147 br_0_147 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c147
+ bl_0_147 br_0_147 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c147
+ bl_0_147 br_0_147 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c147
+ bl_0_147 br_0_147 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c147
+ bl_0_147 br_0_147 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c147
+ bl_0_147 br_0_147 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c147
+ bl_0_147 br_0_147 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c147
+ bl_0_147 br_0_147 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c147
+ bl_0_147 br_0_147 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c147
+ bl_0_147 br_0_147 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c147
+ bl_0_147 br_0_147 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c147
+ bl_0_147 br_0_147 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c147
+ bl_0_147 br_0_147 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c147
+ bl_0_147 br_0_147 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c147
+ bl_0_147 br_0_147 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c147
+ bl_0_147 br_0_147 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c147
+ bl_0_147 br_0_147 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c147
+ bl_0_147 br_0_147 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c147
+ bl_0_147 br_0_147 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c147
+ bl_0_147 br_0_147 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c148
+ bl_0_148 br_0_148 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c148
+ bl_0_148 br_0_148 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c148
+ bl_0_148 br_0_148 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c148
+ bl_0_148 br_0_148 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c148
+ bl_0_148 br_0_148 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c148
+ bl_0_148 br_0_148 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c148
+ bl_0_148 br_0_148 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c148
+ bl_0_148 br_0_148 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c148
+ bl_0_148 br_0_148 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c148
+ bl_0_148 br_0_148 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c148
+ bl_0_148 br_0_148 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c148
+ bl_0_148 br_0_148 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c148
+ bl_0_148 br_0_148 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c148
+ bl_0_148 br_0_148 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c148
+ bl_0_148 br_0_148 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c148
+ bl_0_148 br_0_148 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c148
+ bl_0_148 br_0_148 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c148
+ bl_0_148 br_0_148 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c148
+ bl_0_148 br_0_148 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c148
+ bl_0_148 br_0_148 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c148
+ bl_0_148 br_0_148 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c148
+ bl_0_148 br_0_148 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c148
+ bl_0_148 br_0_148 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c148
+ bl_0_148 br_0_148 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c148
+ bl_0_148 br_0_148 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c148
+ bl_0_148 br_0_148 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c148
+ bl_0_148 br_0_148 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c148
+ bl_0_148 br_0_148 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c148
+ bl_0_148 br_0_148 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c148
+ bl_0_148 br_0_148 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c148
+ bl_0_148 br_0_148 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c148
+ bl_0_148 br_0_148 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c148
+ bl_0_148 br_0_148 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c148
+ bl_0_148 br_0_148 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c148
+ bl_0_148 br_0_148 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c148
+ bl_0_148 br_0_148 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c148
+ bl_0_148 br_0_148 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c148
+ bl_0_148 br_0_148 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c148
+ bl_0_148 br_0_148 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c148
+ bl_0_148 br_0_148 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c148
+ bl_0_148 br_0_148 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c148
+ bl_0_148 br_0_148 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c148
+ bl_0_148 br_0_148 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c148
+ bl_0_148 br_0_148 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c149
+ bl_0_149 br_0_149 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c149
+ bl_0_149 br_0_149 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c149
+ bl_0_149 br_0_149 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c149
+ bl_0_149 br_0_149 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c149
+ bl_0_149 br_0_149 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c149
+ bl_0_149 br_0_149 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c149
+ bl_0_149 br_0_149 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c149
+ bl_0_149 br_0_149 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c149
+ bl_0_149 br_0_149 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c149
+ bl_0_149 br_0_149 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c149
+ bl_0_149 br_0_149 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c149
+ bl_0_149 br_0_149 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c149
+ bl_0_149 br_0_149 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c149
+ bl_0_149 br_0_149 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c149
+ bl_0_149 br_0_149 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c149
+ bl_0_149 br_0_149 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c149
+ bl_0_149 br_0_149 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c149
+ bl_0_149 br_0_149 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c149
+ bl_0_149 br_0_149 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c149
+ bl_0_149 br_0_149 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c149
+ bl_0_149 br_0_149 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c149
+ bl_0_149 br_0_149 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c149
+ bl_0_149 br_0_149 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c149
+ bl_0_149 br_0_149 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c149
+ bl_0_149 br_0_149 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c149
+ bl_0_149 br_0_149 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c149
+ bl_0_149 br_0_149 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c149
+ bl_0_149 br_0_149 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c149
+ bl_0_149 br_0_149 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c149
+ bl_0_149 br_0_149 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c149
+ bl_0_149 br_0_149 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c149
+ bl_0_149 br_0_149 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c149
+ bl_0_149 br_0_149 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c149
+ bl_0_149 br_0_149 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c149
+ bl_0_149 br_0_149 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c149
+ bl_0_149 br_0_149 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c149
+ bl_0_149 br_0_149 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c149
+ bl_0_149 br_0_149 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c149
+ bl_0_149 br_0_149 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c149
+ bl_0_149 br_0_149 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c149
+ bl_0_149 br_0_149 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c149
+ bl_0_149 br_0_149 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c149
+ bl_0_149 br_0_149 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c149
+ bl_0_149 br_0_149 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c150
+ bl_0_150 br_0_150 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c150
+ bl_0_150 br_0_150 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c150
+ bl_0_150 br_0_150 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c150
+ bl_0_150 br_0_150 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c150
+ bl_0_150 br_0_150 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c150
+ bl_0_150 br_0_150 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c150
+ bl_0_150 br_0_150 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c150
+ bl_0_150 br_0_150 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c150
+ bl_0_150 br_0_150 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c150
+ bl_0_150 br_0_150 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c150
+ bl_0_150 br_0_150 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c150
+ bl_0_150 br_0_150 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c150
+ bl_0_150 br_0_150 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c150
+ bl_0_150 br_0_150 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c150
+ bl_0_150 br_0_150 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c150
+ bl_0_150 br_0_150 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c150
+ bl_0_150 br_0_150 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c150
+ bl_0_150 br_0_150 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c150
+ bl_0_150 br_0_150 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c150
+ bl_0_150 br_0_150 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c150
+ bl_0_150 br_0_150 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c150
+ bl_0_150 br_0_150 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c150
+ bl_0_150 br_0_150 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c150
+ bl_0_150 br_0_150 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c150
+ bl_0_150 br_0_150 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c150
+ bl_0_150 br_0_150 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c150
+ bl_0_150 br_0_150 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c150
+ bl_0_150 br_0_150 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c150
+ bl_0_150 br_0_150 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c150
+ bl_0_150 br_0_150 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c150
+ bl_0_150 br_0_150 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c150
+ bl_0_150 br_0_150 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c150
+ bl_0_150 br_0_150 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c150
+ bl_0_150 br_0_150 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c150
+ bl_0_150 br_0_150 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c150
+ bl_0_150 br_0_150 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c150
+ bl_0_150 br_0_150 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c150
+ bl_0_150 br_0_150 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c150
+ bl_0_150 br_0_150 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c150
+ bl_0_150 br_0_150 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c150
+ bl_0_150 br_0_150 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c150
+ bl_0_150 br_0_150 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c150
+ bl_0_150 br_0_150 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c150
+ bl_0_150 br_0_150 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c151
+ bl_0_151 br_0_151 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c151
+ bl_0_151 br_0_151 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c151
+ bl_0_151 br_0_151 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c151
+ bl_0_151 br_0_151 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c151
+ bl_0_151 br_0_151 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c151
+ bl_0_151 br_0_151 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c151
+ bl_0_151 br_0_151 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c151
+ bl_0_151 br_0_151 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c151
+ bl_0_151 br_0_151 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c151
+ bl_0_151 br_0_151 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c151
+ bl_0_151 br_0_151 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c151
+ bl_0_151 br_0_151 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c151
+ bl_0_151 br_0_151 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c151
+ bl_0_151 br_0_151 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c151
+ bl_0_151 br_0_151 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c151
+ bl_0_151 br_0_151 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c151
+ bl_0_151 br_0_151 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c151
+ bl_0_151 br_0_151 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c151
+ bl_0_151 br_0_151 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c151
+ bl_0_151 br_0_151 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c151
+ bl_0_151 br_0_151 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c151
+ bl_0_151 br_0_151 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c151
+ bl_0_151 br_0_151 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c151
+ bl_0_151 br_0_151 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c151
+ bl_0_151 br_0_151 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c151
+ bl_0_151 br_0_151 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c151
+ bl_0_151 br_0_151 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c151
+ bl_0_151 br_0_151 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c151
+ bl_0_151 br_0_151 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c151
+ bl_0_151 br_0_151 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c151
+ bl_0_151 br_0_151 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c151
+ bl_0_151 br_0_151 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c151
+ bl_0_151 br_0_151 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c151
+ bl_0_151 br_0_151 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c151
+ bl_0_151 br_0_151 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c151
+ bl_0_151 br_0_151 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c151
+ bl_0_151 br_0_151 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c151
+ bl_0_151 br_0_151 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c151
+ bl_0_151 br_0_151 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c151
+ bl_0_151 br_0_151 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c151
+ bl_0_151 br_0_151 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c151
+ bl_0_151 br_0_151 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c151
+ bl_0_151 br_0_151 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c151
+ bl_0_151 br_0_151 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c152
+ bl_0_152 br_0_152 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c152
+ bl_0_152 br_0_152 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c152
+ bl_0_152 br_0_152 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c152
+ bl_0_152 br_0_152 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c152
+ bl_0_152 br_0_152 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c152
+ bl_0_152 br_0_152 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c152
+ bl_0_152 br_0_152 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c152
+ bl_0_152 br_0_152 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c152
+ bl_0_152 br_0_152 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c152
+ bl_0_152 br_0_152 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c152
+ bl_0_152 br_0_152 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c152
+ bl_0_152 br_0_152 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c152
+ bl_0_152 br_0_152 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c152
+ bl_0_152 br_0_152 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c152
+ bl_0_152 br_0_152 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c152
+ bl_0_152 br_0_152 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c152
+ bl_0_152 br_0_152 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c152
+ bl_0_152 br_0_152 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c152
+ bl_0_152 br_0_152 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c152
+ bl_0_152 br_0_152 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c152
+ bl_0_152 br_0_152 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c152
+ bl_0_152 br_0_152 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c152
+ bl_0_152 br_0_152 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c152
+ bl_0_152 br_0_152 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c152
+ bl_0_152 br_0_152 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c152
+ bl_0_152 br_0_152 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c152
+ bl_0_152 br_0_152 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c152
+ bl_0_152 br_0_152 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c152
+ bl_0_152 br_0_152 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c152
+ bl_0_152 br_0_152 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c152
+ bl_0_152 br_0_152 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c152
+ bl_0_152 br_0_152 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c152
+ bl_0_152 br_0_152 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c152
+ bl_0_152 br_0_152 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c152
+ bl_0_152 br_0_152 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c152
+ bl_0_152 br_0_152 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c152
+ bl_0_152 br_0_152 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c152
+ bl_0_152 br_0_152 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c152
+ bl_0_152 br_0_152 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c152
+ bl_0_152 br_0_152 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c152
+ bl_0_152 br_0_152 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c152
+ bl_0_152 br_0_152 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c152
+ bl_0_152 br_0_152 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c152
+ bl_0_152 br_0_152 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c153
+ bl_0_153 br_0_153 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c153
+ bl_0_153 br_0_153 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c153
+ bl_0_153 br_0_153 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c153
+ bl_0_153 br_0_153 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c153
+ bl_0_153 br_0_153 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c153
+ bl_0_153 br_0_153 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c153
+ bl_0_153 br_0_153 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c153
+ bl_0_153 br_0_153 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c153
+ bl_0_153 br_0_153 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c153
+ bl_0_153 br_0_153 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c153
+ bl_0_153 br_0_153 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c153
+ bl_0_153 br_0_153 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c153
+ bl_0_153 br_0_153 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c153
+ bl_0_153 br_0_153 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c153
+ bl_0_153 br_0_153 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c153
+ bl_0_153 br_0_153 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c153
+ bl_0_153 br_0_153 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c153
+ bl_0_153 br_0_153 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c153
+ bl_0_153 br_0_153 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c153
+ bl_0_153 br_0_153 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c153
+ bl_0_153 br_0_153 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c153
+ bl_0_153 br_0_153 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c153
+ bl_0_153 br_0_153 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c153
+ bl_0_153 br_0_153 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c153
+ bl_0_153 br_0_153 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c153
+ bl_0_153 br_0_153 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c153
+ bl_0_153 br_0_153 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c153
+ bl_0_153 br_0_153 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c153
+ bl_0_153 br_0_153 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c153
+ bl_0_153 br_0_153 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c153
+ bl_0_153 br_0_153 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c153
+ bl_0_153 br_0_153 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c153
+ bl_0_153 br_0_153 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c153
+ bl_0_153 br_0_153 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c153
+ bl_0_153 br_0_153 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c153
+ bl_0_153 br_0_153 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c153
+ bl_0_153 br_0_153 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c153
+ bl_0_153 br_0_153 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c153
+ bl_0_153 br_0_153 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c153
+ bl_0_153 br_0_153 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c153
+ bl_0_153 br_0_153 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c153
+ bl_0_153 br_0_153 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c153
+ bl_0_153 br_0_153 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c153
+ bl_0_153 br_0_153 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c154
+ bl_0_154 br_0_154 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c154
+ bl_0_154 br_0_154 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c154
+ bl_0_154 br_0_154 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c154
+ bl_0_154 br_0_154 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c154
+ bl_0_154 br_0_154 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c154
+ bl_0_154 br_0_154 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c154
+ bl_0_154 br_0_154 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c154
+ bl_0_154 br_0_154 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c154
+ bl_0_154 br_0_154 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c154
+ bl_0_154 br_0_154 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c154
+ bl_0_154 br_0_154 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c154
+ bl_0_154 br_0_154 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c154
+ bl_0_154 br_0_154 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c154
+ bl_0_154 br_0_154 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c154
+ bl_0_154 br_0_154 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c154
+ bl_0_154 br_0_154 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c154
+ bl_0_154 br_0_154 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c154
+ bl_0_154 br_0_154 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c154
+ bl_0_154 br_0_154 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c154
+ bl_0_154 br_0_154 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c154
+ bl_0_154 br_0_154 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c154
+ bl_0_154 br_0_154 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c154
+ bl_0_154 br_0_154 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c154
+ bl_0_154 br_0_154 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c154
+ bl_0_154 br_0_154 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c154
+ bl_0_154 br_0_154 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c154
+ bl_0_154 br_0_154 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c154
+ bl_0_154 br_0_154 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c154
+ bl_0_154 br_0_154 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c154
+ bl_0_154 br_0_154 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c154
+ bl_0_154 br_0_154 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c154
+ bl_0_154 br_0_154 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c154
+ bl_0_154 br_0_154 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c154
+ bl_0_154 br_0_154 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c154
+ bl_0_154 br_0_154 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c154
+ bl_0_154 br_0_154 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c154
+ bl_0_154 br_0_154 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c154
+ bl_0_154 br_0_154 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c154
+ bl_0_154 br_0_154 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c154
+ bl_0_154 br_0_154 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c154
+ bl_0_154 br_0_154 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c154
+ bl_0_154 br_0_154 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c154
+ bl_0_154 br_0_154 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c154
+ bl_0_154 br_0_154 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c155
+ bl_0_155 br_0_155 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c155
+ bl_0_155 br_0_155 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c155
+ bl_0_155 br_0_155 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c155
+ bl_0_155 br_0_155 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c155
+ bl_0_155 br_0_155 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c155
+ bl_0_155 br_0_155 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c155
+ bl_0_155 br_0_155 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c155
+ bl_0_155 br_0_155 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c155
+ bl_0_155 br_0_155 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c155
+ bl_0_155 br_0_155 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c155
+ bl_0_155 br_0_155 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c155
+ bl_0_155 br_0_155 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c155
+ bl_0_155 br_0_155 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c155
+ bl_0_155 br_0_155 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c155
+ bl_0_155 br_0_155 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c155
+ bl_0_155 br_0_155 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c155
+ bl_0_155 br_0_155 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c155
+ bl_0_155 br_0_155 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c155
+ bl_0_155 br_0_155 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c155
+ bl_0_155 br_0_155 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c155
+ bl_0_155 br_0_155 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c155
+ bl_0_155 br_0_155 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c155
+ bl_0_155 br_0_155 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c155
+ bl_0_155 br_0_155 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c155
+ bl_0_155 br_0_155 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c155
+ bl_0_155 br_0_155 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c155
+ bl_0_155 br_0_155 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c155
+ bl_0_155 br_0_155 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c155
+ bl_0_155 br_0_155 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c155
+ bl_0_155 br_0_155 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c155
+ bl_0_155 br_0_155 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c155
+ bl_0_155 br_0_155 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c155
+ bl_0_155 br_0_155 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c155
+ bl_0_155 br_0_155 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c155
+ bl_0_155 br_0_155 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c155
+ bl_0_155 br_0_155 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c155
+ bl_0_155 br_0_155 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c155
+ bl_0_155 br_0_155 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c155
+ bl_0_155 br_0_155 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c155
+ bl_0_155 br_0_155 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c155
+ bl_0_155 br_0_155 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c155
+ bl_0_155 br_0_155 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c155
+ bl_0_155 br_0_155 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c155
+ bl_0_155 br_0_155 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c156
+ bl_0_156 br_0_156 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c156
+ bl_0_156 br_0_156 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c156
+ bl_0_156 br_0_156 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c156
+ bl_0_156 br_0_156 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c156
+ bl_0_156 br_0_156 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c156
+ bl_0_156 br_0_156 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c156
+ bl_0_156 br_0_156 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c156
+ bl_0_156 br_0_156 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c156
+ bl_0_156 br_0_156 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c156
+ bl_0_156 br_0_156 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c156
+ bl_0_156 br_0_156 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c156
+ bl_0_156 br_0_156 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c156
+ bl_0_156 br_0_156 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c156
+ bl_0_156 br_0_156 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c156
+ bl_0_156 br_0_156 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c156
+ bl_0_156 br_0_156 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c156
+ bl_0_156 br_0_156 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c156
+ bl_0_156 br_0_156 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c156
+ bl_0_156 br_0_156 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c156
+ bl_0_156 br_0_156 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c156
+ bl_0_156 br_0_156 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c156
+ bl_0_156 br_0_156 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c156
+ bl_0_156 br_0_156 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c156
+ bl_0_156 br_0_156 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c156
+ bl_0_156 br_0_156 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c156
+ bl_0_156 br_0_156 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c156
+ bl_0_156 br_0_156 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c156
+ bl_0_156 br_0_156 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c156
+ bl_0_156 br_0_156 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c156
+ bl_0_156 br_0_156 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c156
+ bl_0_156 br_0_156 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c156
+ bl_0_156 br_0_156 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c156
+ bl_0_156 br_0_156 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c156
+ bl_0_156 br_0_156 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c156
+ bl_0_156 br_0_156 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c156
+ bl_0_156 br_0_156 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c156
+ bl_0_156 br_0_156 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c156
+ bl_0_156 br_0_156 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c156
+ bl_0_156 br_0_156 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c156
+ bl_0_156 br_0_156 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c156
+ bl_0_156 br_0_156 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c156
+ bl_0_156 br_0_156 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c156
+ bl_0_156 br_0_156 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c156
+ bl_0_156 br_0_156 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c157
+ bl_0_157 br_0_157 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c157
+ bl_0_157 br_0_157 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c157
+ bl_0_157 br_0_157 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c157
+ bl_0_157 br_0_157 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c157
+ bl_0_157 br_0_157 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c157
+ bl_0_157 br_0_157 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c157
+ bl_0_157 br_0_157 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c157
+ bl_0_157 br_0_157 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c157
+ bl_0_157 br_0_157 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c157
+ bl_0_157 br_0_157 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c157
+ bl_0_157 br_0_157 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c157
+ bl_0_157 br_0_157 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c157
+ bl_0_157 br_0_157 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c157
+ bl_0_157 br_0_157 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c157
+ bl_0_157 br_0_157 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c157
+ bl_0_157 br_0_157 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c157
+ bl_0_157 br_0_157 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c157
+ bl_0_157 br_0_157 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c157
+ bl_0_157 br_0_157 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c157
+ bl_0_157 br_0_157 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c157
+ bl_0_157 br_0_157 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c157
+ bl_0_157 br_0_157 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c157
+ bl_0_157 br_0_157 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c157
+ bl_0_157 br_0_157 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c157
+ bl_0_157 br_0_157 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c157
+ bl_0_157 br_0_157 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c157
+ bl_0_157 br_0_157 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c157
+ bl_0_157 br_0_157 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c157
+ bl_0_157 br_0_157 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c157
+ bl_0_157 br_0_157 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c157
+ bl_0_157 br_0_157 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c157
+ bl_0_157 br_0_157 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c157
+ bl_0_157 br_0_157 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c157
+ bl_0_157 br_0_157 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c157
+ bl_0_157 br_0_157 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c157
+ bl_0_157 br_0_157 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c157
+ bl_0_157 br_0_157 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c157
+ bl_0_157 br_0_157 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c157
+ bl_0_157 br_0_157 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c157
+ bl_0_157 br_0_157 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c157
+ bl_0_157 br_0_157 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c157
+ bl_0_157 br_0_157 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c157
+ bl_0_157 br_0_157 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c157
+ bl_0_157 br_0_157 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c158
+ bl_0_158 br_0_158 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c158
+ bl_0_158 br_0_158 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c158
+ bl_0_158 br_0_158 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c158
+ bl_0_158 br_0_158 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c158
+ bl_0_158 br_0_158 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c158
+ bl_0_158 br_0_158 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c158
+ bl_0_158 br_0_158 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c158
+ bl_0_158 br_0_158 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c158
+ bl_0_158 br_0_158 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c158
+ bl_0_158 br_0_158 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c158
+ bl_0_158 br_0_158 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c158
+ bl_0_158 br_0_158 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c158
+ bl_0_158 br_0_158 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c158
+ bl_0_158 br_0_158 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c158
+ bl_0_158 br_0_158 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c158
+ bl_0_158 br_0_158 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c158
+ bl_0_158 br_0_158 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c158
+ bl_0_158 br_0_158 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c158
+ bl_0_158 br_0_158 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c158
+ bl_0_158 br_0_158 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c158
+ bl_0_158 br_0_158 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c158
+ bl_0_158 br_0_158 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c158
+ bl_0_158 br_0_158 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c158
+ bl_0_158 br_0_158 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c158
+ bl_0_158 br_0_158 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c158
+ bl_0_158 br_0_158 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c158
+ bl_0_158 br_0_158 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c158
+ bl_0_158 br_0_158 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c158
+ bl_0_158 br_0_158 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c158
+ bl_0_158 br_0_158 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c158
+ bl_0_158 br_0_158 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c158
+ bl_0_158 br_0_158 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c158
+ bl_0_158 br_0_158 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c158
+ bl_0_158 br_0_158 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c158
+ bl_0_158 br_0_158 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c158
+ bl_0_158 br_0_158 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c158
+ bl_0_158 br_0_158 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c158
+ bl_0_158 br_0_158 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c158
+ bl_0_158 br_0_158 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c158
+ bl_0_158 br_0_158 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c158
+ bl_0_158 br_0_158 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c158
+ bl_0_158 br_0_158 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c158
+ bl_0_158 br_0_158 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c158
+ bl_0_158 br_0_158 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c159
+ bl_0_159 br_0_159 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c159
+ bl_0_159 br_0_159 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c159
+ bl_0_159 br_0_159 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c159
+ bl_0_159 br_0_159 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c159
+ bl_0_159 br_0_159 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c159
+ bl_0_159 br_0_159 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c159
+ bl_0_159 br_0_159 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c159
+ bl_0_159 br_0_159 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c159
+ bl_0_159 br_0_159 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c159
+ bl_0_159 br_0_159 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c159
+ bl_0_159 br_0_159 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c159
+ bl_0_159 br_0_159 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c159
+ bl_0_159 br_0_159 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c159
+ bl_0_159 br_0_159 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c159
+ bl_0_159 br_0_159 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c159
+ bl_0_159 br_0_159 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c159
+ bl_0_159 br_0_159 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c159
+ bl_0_159 br_0_159 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c159
+ bl_0_159 br_0_159 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c159
+ bl_0_159 br_0_159 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c159
+ bl_0_159 br_0_159 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c159
+ bl_0_159 br_0_159 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c159
+ bl_0_159 br_0_159 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c159
+ bl_0_159 br_0_159 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c159
+ bl_0_159 br_0_159 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c159
+ bl_0_159 br_0_159 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c159
+ bl_0_159 br_0_159 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c159
+ bl_0_159 br_0_159 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c159
+ bl_0_159 br_0_159 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c159
+ bl_0_159 br_0_159 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c159
+ bl_0_159 br_0_159 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c159
+ bl_0_159 br_0_159 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c159
+ bl_0_159 br_0_159 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c159
+ bl_0_159 br_0_159 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c159
+ bl_0_159 br_0_159 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c159
+ bl_0_159 br_0_159 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c159
+ bl_0_159 br_0_159 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c159
+ bl_0_159 br_0_159 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c159
+ bl_0_159 br_0_159 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c159
+ bl_0_159 br_0_159 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c159
+ bl_0_159 br_0_159 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c159
+ bl_0_159 br_0_159 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c159
+ bl_0_159 br_0_159 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c159
+ bl_0_159 br_0_159 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c160
+ bl_0_160 br_0_160 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c160
+ bl_0_160 br_0_160 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c160
+ bl_0_160 br_0_160 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c160
+ bl_0_160 br_0_160 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c160
+ bl_0_160 br_0_160 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c160
+ bl_0_160 br_0_160 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c160
+ bl_0_160 br_0_160 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c160
+ bl_0_160 br_0_160 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c160
+ bl_0_160 br_0_160 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c160
+ bl_0_160 br_0_160 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c160
+ bl_0_160 br_0_160 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c160
+ bl_0_160 br_0_160 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c160
+ bl_0_160 br_0_160 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c160
+ bl_0_160 br_0_160 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c160
+ bl_0_160 br_0_160 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c160
+ bl_0_160 br_0_160 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c160
+ bl_0_160 br_0_160 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c160
+ bl_0_160 br_0_160 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c160
+ bl_0_160 br_0_160 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c160
+ bl_0_160 br_0_160 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c160
+ bl_0_160 br_0_160 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c160
+ bl_0_160 br_0_160 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c160
+ bl_0_160 br_0_160 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c160
+ bl_0_160 br_0_160 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c160
+ bl_0_160 br_0_160 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c160
+ bl_0_160 br_0_160 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c160
+ bl_0_160 br_0_160 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c160
+ bl_0_160 br_0_160 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c160
+ bl_0_160 br_0_160 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c160
+ bl_0_160 br_0_160 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c160
+ bl_0_160 br_0_160 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c160
+ bl_0_160 br_0_160 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c160
+ bl_0_160 br_0_160 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c160
+ bl_0_160 br_0_160 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c160
+ bl_0_160 br_0_160 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c160
+ bl_0_160 br_0_160 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c160
+ bl_0_160 br_0_160 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c160
+ bl_0_160 br_0_160 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c160
+ bl_0_160 br_0_160 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c160
+ bl_0_160 br_0_160 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c160
+ bl_0_160 br_0_160 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c160
+ bl_0_160 br_0_160 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c160
+ bl_0_160 br_0_160 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c160
+ bl_0_160 br_0_160 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c161
+ bl_0_161 br_0_161 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c161
+ bl_0_161 br_0_161 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c161
+ bl_0_161 br_0_161 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c161
+ bl_0_161 br_0_161 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c161
+ bl_0_161 br_0_161 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c161
+ bl_0_161 br_0_161 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c161
+ bl_0_161 br_0_161 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c161
+ bl_0_161 br_0_161 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c161
+ bl_0_161 br_0_161 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c161
+ bl_0_161 br_0_161 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c161
+ bl_0_161 br_0_161 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c161
+ bl_0_161 br_0_161 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c161
+ bl_0_161 br_0_161 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c161
+ bl_0_161 br_0_161 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c161
+ bl_0_161 br_0_161 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c161
+ bl_0_161 br_0_161 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c161
+ bl_0_161 br_0_161 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c161
+ bl_0_161 br_0_161 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c161
+ bl_0_161 br_0_161 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c161
+ bl_0_161 br_0_161 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c161
+ bl_0_161 br_0_161 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c161
+ bl_0_161 br_0_161 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c161
+ bl_0_161 br_0_161 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c161
+ bl_0_161 br_0_161 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c161
+ bl_0_161 br_0_161 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c161
+ bl_0_161 br_0_161 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c161
+ bl_0_161 br_0_161 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c161
+ bl_0_161 br_0_161 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c161
+ bl_0_161 br_0_161 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c161
+ bl_0_161 br_0_161 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c161
+ bl_0_161 br_0_161 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c161
+ bl_0_161 br_0_161 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c161
+ bl_0_161 br_0_161 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c161
+ bl_0_161 br_0_161 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c161
+ bl_0_161 br_0_161 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c161
+ bl_0_161 br_0_161 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c161
+ bl_0_161 br_0_161 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c161
+ bl_0_161 br_0_161 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c161
+ bl_0_161 br_0_161 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c161
+ bl_0_161 br_0_161 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c161
+ bl_0_161 br_0_161 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c161
+ bl_0_161 br_0_161 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c161
+ bl_0_161 br_0_161 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c161
+ bl_0_161 br_0_161 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c162
+ bl_0_162 br_0_162 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c162
+ bl_0_162 br_0_162 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c162
+ bl_0_162 br_0_162 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c162
+ bl_0_162 br_0_162 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c162
+ bl_0_162 br_0_162 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c162
+ bl_0_162 br_0_162 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c162
+ bl_0_162 br_0_162 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c162
+ bl_0_162 br_0_162 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c162
+ bl_0_162 br_0_162 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c162
+ bl_0_162 br_0_162 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c162
+ bl_0_162 br_0_162 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c162
+ bl_0_162 br_0_162 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c162
+ bl_0_162 br_0_162 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c162
+ bl_0_162 br_0_162 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c162
+ bl_0_162 br_0_162 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c162
+ bl_0_162 br_0_162 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c162
+ bl_0_162 br_0_162 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c162
+ bl_0_162 br_0_162 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c162
+ bl_0_162 br_0_162 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c162
+ bl_0_162 br_0_162 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c162
+ bl_0_162 br_0_162 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c162
+ bl_0_162 br_0_162 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c162
+ bl_0_162 br_0_162 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c162
+ bl_0_162 br_0_162 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c162
+ bl_0_162 br_0_162 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c162
+ bl_0_162 br_0_162 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c162
+ bl_0_162 br_0_162 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c162
+ bl_0_162 br_0_162 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c162
+ bl_0_162 br_0_162 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c162
+ bl_0_162 br_0_162 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c162
+ bl_0_162 br_0_162 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c162
+ bl_0_162 br_0_162 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c162
+ bl_0_162 br_0_162 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c162
+ bl_0_162 br_0_162 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c162
+ bl_0_162 br_0_162 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c162
+ bl_0_162 br_0_162 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c162
+ bl_0_162 br_0_162 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c162
+ bl_0_162 br_0_162 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c162
+ bl_0_162 br_0_162 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c162
+ bl_0_162 br_0_162 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c162
+ bl_0_162 br_0_162 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c162
+ bl_0_162 br_0_162 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c162
+ bl_0_162 br_0_162 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c162
+ bl_0_162 br_0_162 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c163
+ bl_0_163 br_0_163 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c163
+ bl_0_163 br_0_163 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c163
+ bl_0_163 br_0_163 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c163
+ bl_0_163 br_0_163 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c163
+ bl_0_163 br_0_163 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c163
+ bl_0_163 br_0_163 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c163
+ bl_0_163 br_0_163 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c163
+ bl_0_163 br_0_163 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c163
+ bl_0_163 br_0_163 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c163
+ bl_0_163 br_0_163 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c163
+ bl_0_163 br_0_163 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c163
+ bl_0_163 br_0_163 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c163
+ bl_0_163 br_0_163 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c163
+ bl_0_163 br_0_163 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c163
+ bl_0_163 br_0_163 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c163
+ bl_0_163 br_0_163 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c163
+ bl_0_163 br_0_163 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c163
+ bl_0_163 br_0_163 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c163
+ bl_0_163 br_0_163 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c163
+ bl_0_163 br_0_163 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c163
+ bl_0_163 br_0_163 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c163
+ bl_0_163 br_0_163 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c163
+ bl_0_163 br_0_163 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c163
+ bl_0_163 br_0_163 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c163
+ bl_0_163 br_0_163 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c163
+ bl_0_163 br_0_163 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c163
+ bl_0_163 br_0_163 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c163
+ bl_0_163 br_0_163 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c163
+ bl_0_163 br_0_163 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c163
+ bl_0_163 br_0_163 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c163
+ bl_0_163 br_0_163 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c163
+ bl_0_163 br_0_163 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c163
+ bl_0_163 br_0_163 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c163
+ bl_0_163 br_0_163 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c163
+ bl_0_163 br_0_163 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c163
+ bl_0_163 br_0_163 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c163
+ bl_0_163 br_0_163 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c163
+ bl_0_163 br_0_163 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c163
+ bl_0_163 br_0_163 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c163
+ bl_0_163 br_0_163 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c163
+ bl_0_163 br_0_163 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c163
+ bl_0_163 br_0_163 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c163
+ bl_0_163 br_0_163 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c163
+ bl_0_163 br_0_163 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c164
+ bl_0_164 br_0_164 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c164
+ bl_0_164 br_0_164 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c164
+ bl_0_164 br_0_164 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c164
+ bl_0_164 br_0_164 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c164
+ bl_0_164 br_0_164 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c164
+ bl_0_164 br_0_164 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c164
+ bl_0_164 br_0_164 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c164
+ bl_0_164 br_0_164 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c164
+ bl_0_164 br_0_164 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c164
+ bl_0_164 br_0_164 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c164
+ bl_0_164 br_0_164 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c164
+ bl_0_164 br_0_164 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c164
+ bl_0_164 br_0_164 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c164
+ bl_0_164 br_0_164 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c164
+ bl_0_164 br_0_164 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c164
+ bl_0_164 br_0_164 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c164
+ bl_0_164 br_0_164 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c164
+ bl_0_164 br_0_164 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c164
+ bl_0_164 br_0_164 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c164
+ bl_0_164 br_0_164 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c164
+ bl_0_164 br_0_164 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c164
+ bl_0_164 br_0_164 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c164
+ bl_0_164 br_0_164 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c164
+ bl_0_164 br_0_164 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c164
+ bl_0_164 br_0_164 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c164
+ bl_0_164 br_0_164 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c164
+ bl_0_164 br_0_164 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c164
+ bl_0_164 br_0_164 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c164
+ bl_0_164 br_0_164 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c164
+ bl_0_164 br_0_164 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c164
+ bl_0_164 br_0_164 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c164
+ bl_0_164 br_0_164 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c164
+ bl_0_164 br_0_164 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c164
+ bl_0_164 br_0_164 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c164
+ bl_0_164 br_0_164 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c164
+ bl_0_164 br_0_164 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c164
+ bl_0_164 br_0_164 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c164
+ bl_0_164 br_0_164 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c164
+ bl_0_164 br_0_164 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c164
+ bl_0_164 br_0_164 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c164
+ bl_0_164 br_0_164 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c164
+ bl_0_164 br_0_164 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c164
+ bl_0_164 br_0_164 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c164
+ bl_0_164 br_0_164 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c165
+ bl_0_165 br_0_165 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c165
+ bl_0_165 br_0_165 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c165
+ bl_0_165 br_0_165 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c165
+ bl_0_165 br_0_165 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c165
+ bl_0_165 br_0_165 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c165
+ bl_0_165 br_0_165 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c165
+ bl_0_165 br_0_165 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c165
+ bl_0_165 br_0_165 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c165
+ bl_0_165 br_0_165 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c165
+ bl_0_165 br_0_165 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c165
+ bl_0_165 br_0_165 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c165
+ bl_0_165 br_0_165 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c165
+ bl_0_165 br_0_165 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c165
+ bl_0_165 br_0_165 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c165
+ bl_0_165 br_0_165 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c165
+ bl_0_165 br_0_165 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c165
+ bl_0_165 br_0_165 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c165
+ bl_0_165 br_0_165 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c165
+ bl_0_165 br_0_165 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c165
+ bl_0_165 br_0_165 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c165
+ bl_0_165 br_0_165 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c165
+ bl_0_165 br_0_165 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c165
+ bl_0_165 br_0_165 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c165
+ bl_0_165 br_0_165 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c165
+ bl_0_165 br_0_165 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c165
+ bl_0_165 br_0_165 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c165
+ bl_0_165 br_0_165 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c165
+ bl_0_165 br_0_165 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c165
+ bl_0_165 br_0_165 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c165
+ bl_0_165 br_0_165 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c165
+ bl_0_165 br_0_165 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c165
+ bl_0_165 br_0_165 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c165
+ bl_0_165 br_0_165 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c165
+ bl_0_165 br_0_165 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c165
+ bl_0_165 br_0_165 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c165
+ bl_0_165 br_0_165 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c165
+ bl_0_165 br_0_165 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c165
+ bl_0_165 br_0_165 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c165
+ bl_0_165 br_0_165 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c165
+ bl_0_165 br_0_165 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c165
+ bl_0_165 br_0_165 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c165
+ bl_0_165 br_0_165 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c165
+ bl_0_165 br_0_165 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c165
+ bl_0_165 br_0_165 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c166
+ bl_0_166 br_0_166 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c166
+ bl_0_166 br_0_166 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c166
+ bl_0_166 br_0_166 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c166
+ bl_0_166 br_0_166 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c166
+ bl_0_166 br_0_166 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c166
+ bl_0_166 br_0_166 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c166
+ bl_0_166 br_0_166 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c166
+ bl_0_166 br_0_166 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c166
+ bl_0_166 br_0_166 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c166
+ bl_0_166 br_0_166 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c166
+ bl_0_166 br_0_166 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c166
+ bl_0_166 br_0_166 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c166
+ bl_0_166 br_0_166 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c166
+ bl_0_166 br_0_166 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c166
+ bl_0_166 br_0_166 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c166
+ bl_0_166 br_0_166 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c166
+ bl_0_166 br_0_166 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c166
+ bl_0_166 br_0_166 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c166
+ bl_0_166 br_0_166 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c166
+ bl_0_166 br_0_166 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c166
+ bl_0_166 br_0_166 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c166
+ bl_0_166 br_0_166 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c166
+ bl_0_166 br_0_166 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c166
+ bl_0_166 br_0_166 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c166
+ bl_0_166 br_0_166 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c166
+ bl_0_166 br_0_166 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c166
+ bl_0_166 br_0_166 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c166
+ bl_0_166 br_0_166 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c166
+ bl_0_166 br_0_166 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c166
+ bl_0_166 br_0_166 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c166
+ bl_0_166 br_0_166 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c166
+ bl_0_166 br_0_166 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c166
+ bl_0_166 br_0_166 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c166
+ bl_0_166 br_0_166 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c166
+ bl_0_166 br_0_166 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c166
+ bl_0_166 br_0_166 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c166
+ bl_0_166 br_0_166 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c166
+ bl_0_166 br_0_166 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c166
+ bl_0_166 br_0_166 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c166
+ bl_0_166 br_0_166 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c166
+ bl_0_166 br_0_166 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c166
+ bl_0_166 br_0_166 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c166
+ bl_0_166 br_0_166 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c166
+ bl_0_166 br_0_166 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c167
+ bl_0_167 br_0_167 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c167
+ bl_0_167 br_0_167 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c167
+ bl_0_167 br_0_167 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c167
+ bl_0_167 br_0_167 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c167
+ bl_0_167 br_0_167 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c167
+ bl_0_167 br_0_167 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c167
+ bl_0_167 br_0_167 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c167
+ bl_0_167 br_0_167 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c167
+ bl_0_167 br_0_167 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c167
+ bl_0_167 br_0_167 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c167
+ bl_0_167 br_0_167 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c167
+ bl_0_167 br_0_167 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c167
+ bl_0_167 br_0_167 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c167
+ bl_0_167 br_0_167 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c167
+ bl_0_167 br_0_167 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c167
+ bl_0_167 br_0_167 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c167
+ bl_0_167 br_0_167 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c167
+ bl_0_167 br_0_167 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c167
+ bl_0_167 br_0_167 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c167
+ bl_0_167 br_0_167 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c167
+ bl_0_167 br_0_167 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c167
+ bl_0_167 br_0_167 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c167
+ bl_0_167 br_0_167 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c167
+ bl_0_167 br_0_167 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c167
+ bl_0_167 br_0_167 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c167
+ bl_0_167 br_0_167 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c167
+ bl_0_167 br_0_167 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c167
+ bl_0_167 br_0_167 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c167
+ bl_0_167 br_0_167 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c167
+ bl_0_167 br_0_167 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c167
+ bl_0_167 br_0_167 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c167
+ bl_0_167 br_0_167 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c167
+ bl_0_167 br_0_167 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c167
+ bl_0_167 br_0_167 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c167
+ bl_0_167 br_0_167 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c167
+ bl_0_167 br_0_167 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c167
+ bl_0_167 br_0_167 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c167
+ bl_0_167 br_0_167 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c167
+ bl_0_167 br_0_167 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c167
+ bl_0_167 br_0_167 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c167
+ bl_0_167 br_0_167 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c167
+ bl_0_167 br_0_167 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c167
+ bl_0_167 br_0_167 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c167
+ bl_0_167 br_0_167 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c168
+ bl_0_168 br_0_168 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c168
+ bl_0_168 br_0_168 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c168
+ bl_0_168 br_0_168 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c168
+ bl_0_168 br_0_168 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c168
+ bl_0_168 br_0_168 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c168
+ bl_0_168 br_0_168 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c168
+ bl_0_168 br_0_168 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c168
+ bl_0_168 br_0_168 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c168
+ bl_0_168 br_0_168 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c168
+ bl_0_168 br_0_168 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c168
+ bl_0_168 br_0_168 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c168
+ bl_0_168 br_0_168 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c168
+ bl_0_168 br_0_168 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c168
+ bl_0_168 br_0_168 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c168
+ bl_0_168 br_0_168 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c168
+ bl_0_168 br_0_168 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c168
+ bl_0_168 br_0_168 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c168
+ bl_0_168 br_0_168 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c168
+ bl_0_168 br_0_168 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c168
+ bl_0_168 br_0_168 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c168
+ bl_0_168 br_0_168 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c168
+ bl_0_168 br_0_168 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c168
+ bl_0_168 br_0_168 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c168
+ bl_0_168 br_0_168 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c168
+ bl_0_168 br_0_168 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c168
+ bl_0_168 br_0_168 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c168
+ bl_0_168 br_0_168 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c168
+ bl_0_168 br_0_168 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c168
+ bl_0_168 br_0_168 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c168
+ bl_0_168 br_0_168 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c168
+ bl_0_168 br_0_168 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c168
+ bl_0_168 br_0_168 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c168
+ bl_0_168 br_0_168 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c168
+ bl_0_168 br_0_168 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c168
+ bl_0_168 br_0_168 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c168
+ bl_0_168 br_0_168 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c168
+ bl_0_168 br_0_168 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c168
+ bl_0_168 br_0_168 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c168
+ bl_0_168 br_0_168 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c168
+ bl_0_168 br_0_168 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c168
+ bl_0_168 br_0_168 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c168
+ bl_0_168 br_0_168 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c168
+ bl_0_168 br_0_168 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c168
+ bl_0_168 br_0_168 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c169
+ bl_0_169 br_0_169 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c169
+ bl_0_169 br_0_169 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c169
+ bl_0_169 br_0_169 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c169
+ bl_0_169 br_0_169 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c169
+ bl_0_169 br_0_169 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c169
+ bl_0_169 br_0_169 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c169
+ bl_0_169 br_0_169 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c169
+ bl_0_169 br_0_169 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c169
+ bl_0_169 br_0_169 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c169
+ bl_0_169 br_0_169 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c169
+ bl_0_169 br_0_169 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c169
+ bl_0_169 br_0_169 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c169
+ bl_0_169 br_0_169 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c169
+ bl_0_169 br_0_169 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c169
+ bl_0_169 br_0_169 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c169
+ bl_0_169 br_0_169 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c169
+ bl_0_169 br_0_169 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c169
+ bl_0_169 br_0_169 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c169
+ bl_0_169 br_0_169 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c169
+ bl_0_169 br_0_169 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c169
+ bl_0_169 br_0_169 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c169
+ bl_0_169 br_0_169 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c169
+ bl_0_169 br_0_169 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c169
+ bl_0_169 br_0_169 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c169
+ bl_0_169 br_0_169 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c169
+ bl_0_169 br_0_169 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c169
+ bl_0_169 br_0_169 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c169
+ bl_0_169 br_0_169 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c169
+ bl_0_169 br_0_169 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c169
+ bl_0_169 br_0_169 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c169
+ bl_0_169 br_0_169 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c169
+ bl_0_169 br_0_169 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c169
+ bl_0_169 br_0_169 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c169
+ bl_0_169 br_0_169 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c169
+ bl_0_169 br_0_169 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c169
+ bl_0_169 br_0_169 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c169
+ bl_0_169 br_0_169 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c169
+ bl_0_169 br_0_169 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c169
+ bl_0_169 br_0_169 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c169
+ bl_0_169 br_0_169 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c169
+ bl_0_169 br_0_169 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c169
+ bl_0_169 br_0_169 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c169
+ bl_0_169 br_0_169 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c169
+ bl_0_169 br_0_169 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c170
+ bl_0_170 br_0_170 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c170
+ bl_0_170 br_0_170 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c170
+ bl_0_170 br_0_170 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c170
+ bl_0_170 br_0_170 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c170
+ bl_0_170 br_0_170 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c170
+ bl_0_170 br_0_170 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c170
+ bl_0_170 br_0_170 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c170
+ bl_0_170 br_0_170 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c170
+ bl_0_170 br_0_170 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c170
+ bl_0_170 br_0_170 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c170
+ bl_0_170 br_0_170 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c170
+ bl_0_170 br_0_170 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c170
+ bl_0_170 br_0_170 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c170
+ bl_0_170 br_0_170 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c170
+ bl_0_170 br_0_170 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c170
+ bl_0_170 br_0_170 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c170
+ bl_0_170 br_0_170 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c170
+ bl_0_170 br_0_170 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c170
+ bl_0_170 br_0_170 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c170
+ bl_0_170 br_0_170 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c170
+ bl_0_170 br_0_170 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c170
+ bl_0_170 br_0_170 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c170
+ bl_0_170 br_0_170 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c170
+ bl_0_170 br_0_170 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c170
+ bl_0_170 br_0_170 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c170
+ bl_0_170 br_0_170 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c170
+ bl_0_170 br_0_170 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c170
+ bl_0_170 br_0_170 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c170
+ bl_0_170 br_0_170 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c170
+ bl_0_170 br_0_170 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c170
+ bl_0_170 br_0_170 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c170
+ bl_0_170 br_0_170 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c170
+ bl_0_170 br_0_170 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c170
+ bl_0_170 br_0_170 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c170
+ bl_0_170 br_0_170 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c170
+ bl_0_170 br_0_170 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c170
+ bl_0_170 br_0_170 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c170
+ bl_0_170 br_0_170 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c170
+ bl_0_170 br_0_170 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c170
+ bl_0_170 br_0_170 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c170
+ bl_0_170 br_0_170 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c170
+ bl_0_170 br_0_170 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c170
+ bl_0_170 br_0_170 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c170
+ bl_0_170 br_0_170 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c171
+ bl_0_171 br_0_171 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c171
+ bl_0_171 br_0_171 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c171
+ bl_0_171 br_0_171 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c171
+ bl_0_171 br_0_171 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c171
+ bl_0_171 br_0_171 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c171
+ bl_0_171 br_0_171 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c171
+ bl_0_171 br_0_171 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c171
+ bl_0_171 br_0_171 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c171
+ bl_0_171 br_0_171 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c171
+ bl_0_171 br_0_171 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c171
+ bl_0_171 br_0_171 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c171
+ bl_0_171 br_0_171 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c171
+ bl_0_171 br_0_171 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c171
+ bl_0_171 br_0_171 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c171
+ bl_0_171 br_0_171 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c171
+ bl_0_171 br_0_171 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c171
+ bl_0_171 br_0_171 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c171
+ bl_0_171 br_0_171 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c171
+ bl_0_171 br_0_171 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c171
+ bl_0_171 br_0_171 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c171
+ bl_0_171 br_0_171 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c171
+ bl_0_171 br_0_171 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c171
+ bl_0_171 br_0_171 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c171
+ bl_0_171 br_0_171 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c171
+ bl_0_171 br_0_171 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c171
+ bl_0_171 br_0_171 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c171
+ bl_0_171 br_0_171 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c171
+ bl_0_171 br_0_171 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c171
+ bl_0_171 br_0_171 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c171
+ bl_0_171 br_0_171 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c171
+ bl_0_171 br_0_171 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c171
+ bl_0_171 br_0_171 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c171
+ bl_0_171 br_0_171 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c171
+ bl_0_171 br_0_171 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c171
+ bl_0_171 br_0_171 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c171
+ bl_0_171 br_0_171 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c171
+ bl_0_171 br_0_171 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c171
+ bl_0_171 br_0_171 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c171
+ bl_0_171 br_0_171 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c171
+ bl_0_171 br_0_171 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c171
+ bl_0_171 br_0_171 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c171
+ bl_0_171 br_0_171 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c171
+ bl_0_171 br_0_171 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c171
+ bl_0_171 br_0_171 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c172
+ bl_0_172 br_0_172 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c172
+ bl_0_172 br_0_172 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c172
+ bl_0_172 br_0_172 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c172
+ bl_0_172 br_0_172 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c172
+ bl_0_172 br_0_172 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c172
+ bl_0_172 br_0_172 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c172
+ bl_0_172 br_0_172 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c172
+ bl_0_172 br_0_172 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c172
+ bl_0_172 br_0_172 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c172
+ bl_0_172 br_0_172 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c172
+ bl_0_172 br_0_172 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c172
+ bl_0_172 br_0_172 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c172
+ bl_0_172 br_0_172 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c172
+ bl_0_172 br_0_172 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c172
+ bl_0_172 br_0_172 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c172
+ bl_0_172 br_0_172 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c172
+ bl_0_172 br_0_172 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c172
+ bl_0_172 br_0_172 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c172
+ bl_0_172 br_0_172 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c172
+ bl_0_172 br_0_172 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c172
+ bl_0_172 br_0_172 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c172
+ bl_0_172 br_0_172 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c172
+ bl_0_172 br_0_172 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c172
+ bl_0_172 br_0_172 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c172
+ bl_0_172 br_0_172 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c172
+ bl_0_172 br_0_172 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c172
+ bl_0_172 br_0_172 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c172
+ bl_0_172 br_0_172 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c172
+ bl_0_172 br_0_172 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c172
+ bl_0_172 br_0_172 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c172
+ bl_0_172 br_0_172 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c172
+ bl_0_172 br_0_172 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c172
+ bl_0_172 br_0_172 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c172
+ bl_0_172 br_0_172 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c172
+ bl_0_172 br_0_172 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c172
+ bl_0_172 br_0_172 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c172
+ bl_0_172 br_0_172 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c172
+ bl_0_172 br_0_172 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c172
+ bl_0_172 br_0_172 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c172
+ bl_0_172 br_0_172 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c172
+ bl_0_172 br_0_172 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c172
+ bl_0_172 br_0_172 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c172
+ bl_0_172 br_0_172 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c172
+ bl_0_172 br_0_172 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c173
+ bl_0_173 br_0_173 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c173
+ bl_0_173 br_0_173 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c173
+ bl_0_173 br_0_173 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c173
+ bl_0_173 br_0_173 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c173
+ bl_0_173 br_0_173 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c173
+ bl_0_173 br_0_173 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c173
+ bl_0_173 br_0_173 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c173
+ bl_0_173 br_0_173 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c173
+ bl_0_173 br_0_173 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c173
+ bl_0_173 br_0_173 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c173
+ bl_0_173 br_0_173 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c173
+ bl_0_173 br_0_173 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c173
+ bl_0_173 br_0_173 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c173
+ bl_0_173 br_0_173 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c173
+ bl_0_173 br_0_173 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c173
+ bl_0_173 br_0_173 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c173
+ bl_0_173 br_0_173 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c173
+ bl_0_173 br_0_173 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c173
+ bl_0_173 br_0_173 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c173
+ bl_0_173 br_0_173 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c173
+ bl_0_173 br_0_173 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c173
+ bl_0_173 br_0_173 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c173
+ bl_0_173 br_0_173 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c173
+ bl_0_173 br_0_173 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c173
+ bl_0_173 br_0_173 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c173
+ bl_0_173 br_0_173 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c173
+ bl_0_173 br_0_173 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c173
+ bl_0_173 br_0_173 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c173
+ bl_0_173 br_0_173 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c173
+ bl_0_173 br_0_173 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c173
+ bl_0_173 br_0_173 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c173
+ bl_0_173 br_0_173 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c173
+ bl_0_173 br_0_173 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c173
+ bl_0_173 br_0_173 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c173
+ bl_0_173 br_0_173 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c173
+ bl_0_173 br_0_173 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c173
+ bl_0_173 br_0_173 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c173
+ bl_0_173 br_0_173 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c173
+ bl_0_173 br_0_173 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c173
+ bl_0_173 br_0_173 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c173
+ bl_0_173 br_0_173 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c173
+ bl_0_173 br_0_173 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c173
+ bl_0_173 br_0_173 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c173
+ bl_0_173 br_0_173 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c174
+ bl_0_174 br_0_174 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c174
+ bl_0_174 br_0_174 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c174
+ bl_0_174 br_0_174 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c174
+ bl_0_174 br_0_174 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c174
+ bl_0_174 br_0_174 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c174
+ bl_0_174 br_0_174 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c174
+ bl_0_174 br_0_174 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c174
+ bl_0_174 br_0_174 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c174
+ bl_0_174 br_0_174 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c174
+ bl_0_174 br_0_174 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c174
+ bl_0_174 br_0_174 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c174
+ bl_0_174 br_0_174 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c174
+ bl_0_174 br_0_174 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c174
+ bl_0_174 br_0_174 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c174
+ bl_0_174 br_0_174 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c174
+ bl_0_174 br_0_174 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c174
+ bl_0_174 br_0_174 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c174
+ bl_0_174 br_0_174 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c174
+ bl_0_174 br_0_174 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c174
+ bl_0_174 br_0_174 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c174
+ bl_0_174 br_0_174 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c174
+ bl_0_174 br_0_174 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c174
+ bl_0_174 br_0_174 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c174
+ bl_0_174 br_0_174 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c174
+ bl_0_174 br_0_174 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c174
+ bl_0_174 br_0_174 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c174
+ bl_0_174 br_0_174 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c174
+ bl_0_174 br_0_174 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c174
+ bl_0_174 br_0_174 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c174
+ bl_0_174 br_0_174 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c174
+ bl_0_174 br_0_174 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c174
+ bl_0_174 br_0_174 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c174
+ bl_0_174 br_0_174 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c174
+ bl_0_174 br_0_174 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c174
+ bl_0_174 br_0_174 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c174
+ bl_0_174 br_0_174 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c174
+ bl_0_174 br_0_174 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c174
+ bl_0_174 br_0_174 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c174
+ bl_0_174 br_0_174 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c174
+ bl_0_174 br_0_174 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c174
+ bl_0_174 br_0_174 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c174
+ bl_0_174 br_0_174 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c174
+ bl_0_174 br_0_174 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c174
+ bl_0_174 br_0_174 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c175
+ bl_0_175 br_0_175 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c175
+ bl_0_175 br_0_175 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c175
+ bl_0_175 br_0_175 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c175
+ bl_0_175 br_0_175 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c175
+ bl_0_175 br_0_175 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c175
+ bl_0_175 br_0_175 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c175
+ bl_0_175 br_0_175 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c175
+ bl_0_175 br_0_175 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c175
+ bl_0_175 br_0_175 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c175
+ bl_0_175 br_0_175 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c175
+ bl_0_175 br_0_175 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c175
+ bl_0_175 br_0_175 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c175
+ bl_0_175 br_0_175 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c175
+ bl_0_175 br_0_175 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c175
+ bl_0_175 br_0_175 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c175
+ bl_0_175 br_0_175 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c175
+ bl_0_175 br_0_175 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c175
+ bl_0_175 br_0_175 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c175
+ bl_0_175 br_0_175 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c175
+ bl_0_175 br_0_175 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c175
+ bl_0_175 br_0_175 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c175
+ bl_0_175 br_0_175 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c175
+ bl_0_175 br_0_175 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c175
+ bl_0_175 br_0_175 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c175
+ bl_0_175 br_0_175 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c175
+ bl_0_175 br_0_175 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c175
+ bl_0_175 br_0_175 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c175
+ bl_0_175 br_0_175 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c175
+ bl_0_175 br_0_175 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c175
+ bl_0_175 br_0_175 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c175
+ bl_0_175 br_0_175 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c175
+ bl_0_175 br_0_175 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c175
+ bl_0_175 br_0_175 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c175
+ bl_0_175 br_0_175 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c175
+ bl_0_175 br_0_175 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c175
+ bl_0_175 br_0_175 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c175
+ bl_0_175 br_0_175 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c175
+ bl_0_175 br_0_175 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c175
+ bl_0_175 br_0_175 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c175
+ bl_0_175 br_0_175 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c175
+ bl_0_175 br_0_175 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c175
+ bl_0_175 br_0_175 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c175
+ bl_0_175 br_0_175 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c175
+ bl_0_175 br_0_175 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c176
+ bl_0_176 br_0_176 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c176
+ bl_0_176 br_0_176 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c176
+ bl_0_176 br_0_176 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c176
+ bl_0_176 br_0_176 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c176
+ bl_0_176 br_0_176 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c176
+ bl_0_176 br_0_176 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c176
+ bl_0_176 br_0_176 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c176
+ bl_0_176 br_0_176 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c176
+ bl_0_176 br_0_176 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c176
+ bl_0_176 br_0_176 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c176
+ bl_0_176 br_0_176 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c176
+ bl_0_176 br_0_176 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c176
+ bl_0_176 br_0_176 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c176
+ bl_0_176 br_0_176 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c176
+ bl_0_176 br_0_176 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c176
+ bl_0_176 br_0_176 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c176
+ bl_0_176 br_0_176 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c176
+ bl_0_176 br_0_176 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c176
+ bl_0_176 br_0_176 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c176
+ bl_0_176 br_0_176 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c176
+ bl_0_176 br_0_176 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c176
+ bl_0_176 br_0_176 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c176
+ bl_0_176 br_0_176 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c176
+ bl_0_176 br_0_176 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c176
+ bl_0_176 br_0_176 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c176
+ bl_0_176 br_0_176 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c176
+ bl_0_176 br_0_176 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c176
+ bl_0_176 br_0_176 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c176
+ bl_0_176 br_0_176 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c176
+ bl_0_176 br_0_176 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c176
+ bl_0_176 br_0_176 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c176
+ bl_0_176 br_0_176 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c176
+ bl_0_176 br_0_176 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c176
+ bl_0_176 br_0_176 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c176
+ bl_0_176 br_0_176 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c176
+ bl_0_176 br_0_176 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c176
+ bl_0_176 br_0_176 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c176
+ bl_0_176 br_0_176 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c176
+ bl_0_176 br_0_176 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c176
+ bl_0_176 br_0_176 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c176
+ bl_0_176 br_0_176 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c176
+ bl_0_176 br_0_176 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c176
+ bl_0_176 br_0_176 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c176
+ bl_0_176 br_0_176 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c177
+ bl_0_177 br_0_177 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c177
+ bl_0_177 br_0_177 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c177
+ bl_0_177 br_0_177 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c177
+ bl_0_177 br_0_177 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c177
+ bl_0_177 br_0_177 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c177
+ bl_0_177 br_0_177 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c177
+ bl_0_177 br_0_177 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c177
+ bl_0_177 br_0_177 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c177
+ bl_0_177 br_0_177 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c177
+ bl_0_177 br_0_177 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c177
+ bl_0_177 br_0_177 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c177
+ bl_0_177 br_0_177 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c177
+ bl_0_177 br_0_177 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c177
+ bl_0_177 br_0_177 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c177
+ bl_0_177 br_0_177 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c177
+ bl_0_177 br_0_177 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c177
+ bl_0_177 br_0_177 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c177
+ bl_0_177 br_0_177 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c177
+ bl_0_177 br_0_177 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c177
+ bl_0_177 br_0_177 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c177
+ bl_0_177 br_0_177 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c177
+ bl_0_177 br_0_177 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c177
+ bl_0_177 br_0_177 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c177
+ bl_0_177 br_0_177 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c177
+ bl_0_177 br_0_177 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c177
+ bl_0_177 br_0_177 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c177
+ bl_0_177 br_0_177 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c177
+ bl_0_177 br_0_177 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c177
+ bl_0_177 br_0_177 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c177
+ bl_0_177 br_0_177 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c177
+ bl_0_177 br_0_177 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c177
+ bl_0_177 br_0_177 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c177
+ bl_0_177 br_0_177 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c177
+ bl_0_177 br_0_177 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c177
+ bl_0_177 br_0_177 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c177
+ bl_0_177 br_0_177 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c177
+ bl_0_177 br_0_177 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c177
+ bl_0_177 br_0_177 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c177
+ bl_0_177 br_0_177 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c177
+ bl_0_177 br_0_177 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c177
+ bl_0_177 br_0_177 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c177
+ bl_0_177 br_0_177 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c177
+ bl_0_177 br_0_177 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c177
+ bl_0_177 br_0_177 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c178
+ bl_0_178 br_0_178 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c178
+ bl_0_178 br_0_178 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c178
+ bl_0_178 br_0_178 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c178
+ bl_0_178 br_0_178 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c178
+ bl_0_178 br_0_178 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c178
+ bl_0_178 br_0_178 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c178
+ bl_0_178 br_0_178 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c178
+ bl_0_178 br_0_178 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c178
+ bl_0_178 br_0_178 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c178
+ bl_0_178 br_0_178 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c178
+ bl_0_178 br_0_178 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c178
+ bl_0_178 br_0_178 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c178
+ bl_0_178 br_0_178 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c178
+ bl_0_178 br_0_178 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c178
+ bl_0_178 br_0_178 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c178
+ bl_0_178 br_0_178 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c178
+ bl_0_178 br_0_178 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c178
+ bl_0_178 br_0_178 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c178
+ bl_0_178 br_0_178 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c178
+ bl_0_178 br_0_178 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c178
+ bl_0_178 br_0_178 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c178
+ bl_0_178 br_0_178 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c178
+ bl_0_178 br_0_178 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c178
+ bl_0_178 br_0_178 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c178
+ bl_0_178 br_0_178 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c178
+ bl_0_178 br_0_178 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c178
+ bl_0_178 br_0_178 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c178
+ bl_0_178 br_0_178 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c178
+ bl_0_178 br_0_178 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c178
+ bl_0_178 br_0_178 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c178
+ bl_0_178 br_0_178 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c178
+ bl_0_178 br_0_178 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c178
+ bl_0_178 br_0_178 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c178
+ bl_0_178 br_0_178 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c178
+ bl_0_178 br_0_178 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c178
+ bl_0_178 br_0_178 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c178
+ bl_0_178 br_0_178 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c178
+ bl_0_178 br_0_178 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c178
+ bl_0_178 br_0_178 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c178
+ bl_0_178 br_0_178 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c178
+ bl_0_178 br_0_178 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c178
+ bl_0_178 br_0_178 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c178
+ bl_0_178 br_0_178 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c178
+ bl_0_178 br_0_178 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c179
+ bl_0_179 br_0_179 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c179
+ bl_0_179 br_0_179 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c179
+ bl_0_179 br_0_179 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c179
+ bl_0_179 br_0_179 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c179
+ bl_0_179 br_0_179 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c179
+ bl_0_179 br_0_179 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c179
+ bl_0_179 br_0_179 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c179
+ bl_0_179 br_0_179 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c179
+ bl_0_179 br_0_179 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c179
+ bl_0_179 br_0_179 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c179
+ bl_0_179 br_0_179 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c179
+ bl_0_179 br_0_179 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c179
+ bl_0_179 br_0_179 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c179
+ bl_0_179 br_0_179 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c179
+ bl_0_179 br_0_179 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c179
+ bl_0_179 br_0_179 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c179
+ bl_0_179 br_0_179 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c179
+ bl_0_179 br_0_179 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c179
+ bl_0_179 br_0_179 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c179
+ bl_0_179 br_0_179 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c179
+ bl_0_179 br_0_179 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c179
+ bl_0_179 br_0_179 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c179
+ bl_0_179 br_0_179 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c179
+ bl_0_179 br_0_179 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c179
+ bl_0_179 br_0_179 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c179
+ bl_0_179 br_0_179 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c179
+ bl_0_179 br_0_179 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c179
+ bl_0_179 br_0_179 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c179
+ bl_0_179 br_0_179 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c179
+ bl_0_179 br_0_179 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c179
+ bl_0_179 br_0_179 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c179
+ bl_0_179 br_0_179 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c179
+ bl_0_179 br_0_179 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c179
+ bl_0_179 br_0_179 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c179
+ bl_0_179 br_0_179 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c179
+ bl_0_179 br_0_179 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c179
+ bl_0_179 br_0_179 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c179
+ bl_0_179 br_0_179 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c179
+ bl_0_179 br_0_179 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c179
+ bl_0_179 br_0_179 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c179
+ bl_0_179 br_0_179 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c179
+ bl_0_179 br_0_179 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c179
+ bl_0_179 br_0_179 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c179
+ bl_0_179 br_0_179 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c180
+ bl_0_180 br_0_180 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c180
+ bl_0_180 br_0_180 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c180
+ bl_0_180 br_0_180 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c180
+ bl_0_180 br_0_180 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c180
+ bl_0_180 br_0_180 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c180
+ bl_0_180 br_0_180 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c180
+ bl_0_180 br_0_180 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c180
+ bl_0_180 br_0_180 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c180
+ bl_0_180 br_0_180 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c180
+ bl_0_180 br_0_180 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c180
+ bl_0_180 br_0_180 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c180
+ bl_0_180 br_0_180 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c180
+ bl_0_180 br_0_180 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c180
+ bl_0_180 br_0_180 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c180
+ bl_0_180 br_0_180 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c180
+ bl_0_180 br_0_180 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c180
+ bl_0_180 br_0_180 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c180
+ bl_0_180 br_0_180 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c180
+ bl_0_180 br_0_180 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c180
+ bl_0_180 br_0_180 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c180
+ bl_0_180 br_0_180 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c180
+ bl_0_180 br_0_180 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c180
+ bl_0_180 br_0_180 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c180
+ bl_0_180 br_0_180 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c180
+ bl_0_180 br_0_180 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c180
+ bl_0_180 br_0_180 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c180
+ bl_0_180 br_0_180 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c180
+ bl_0_180 br_0_180 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c180
+ bl_0_180 br_0_180 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c180
+ bl_0_180 br_0_180 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c180
+ bl_0_180 br_0_180 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c180
+ bl_0_180 br_0_180 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c180
+ bl_0_180 br_0_180 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c180
+ bl_0_180 br_0_180 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c180
+ bl_0_180 br_0_180 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c180
+ bl_0_180 br_0_180 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c180
+ bl_0_180 br_0_180 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c180
+ bl_0_180 br_0_180 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c180
+ bl_0_180 br_0_180 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c180
+ bl_0_180 br_0_180 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c180
+ bl_0_180 br_0_180 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c180
+ bl_0_180 br_0_180 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c180
+ bl_0_180 br_0_180 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c180
+ bl_0_180 br_0_180 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c181
+ bl_0_181 br_0_181 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c181
+ bl_0_181 br_0_181 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c181
+ bl_0_181 br_0_181 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c181
+ bl_0_181 br_0_181 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c181
+ bl_0_181 br_0_181 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c181
+ bl_0_181 br_0_181 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c181
+ bl_0_181 br_0_181 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c181
+ bl_0_181 br_0_181 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c181
+ bl_0_181 br_0_181 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c181
+ bl_0_181 br_0_181 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c181
+ bl_0_181 br_0_181 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c181
+ bl_0_181 br_0_181 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c181
+ bl_0_181 br_0_181 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c181
+ bl_0_181 br_0_181 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c181
+ bl_0_181 br_0_181 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c181
+ bl_0_181 br_0_181 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c181
+ bl_0_181 br_0_181 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c181
+ bl_0_181 br_0_181 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c181
+ bl_0_181 br_0_181 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c181
+ bl_0_181 br_0_181 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c181
+ bl_0_181 br_0_181 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c181
+ bl_0_181 br_0_181 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c181
+ bl_0_181 br_0_181 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c181
+ bl_0_181 br_0_181 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c181
+ bl_0_181 br_0_181 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c181
+ bl_0_181 br_0_181 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c181
+ bl_0_181 br_0_181 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c181
+ bl_0_181 br_0_181 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c181
+ bl_0_181 br_0_181 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c181
+ bl_0_181 br_0_181 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c181
+ bl_0_181 br_0_181 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c181
+ bl_0_181 br_0_181 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c181
+ bl_0_181 br_0_181 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c181
+ bl_0_181 br_0_181 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c181
+ bl_0_181 br_0_181 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c181
+ bl_0_181 br_0_181 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c181
+ bl_0_181 br_0_181 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c181
+ bl_0_181 br_0_181 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c181
+ bl_0_181 br_0_181 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c181
+ bl_0_181 br_0_181 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c181
+ bl_0_181 br_0_181 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c181
+ bl_0_181 br_0_181 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c181
+ bl_0_181 br_0_181 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c181
+ bl_0_181 br_0_181 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c182
+ bl_0_182 br_0_182 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c182
+ bl_0_182 br_0_182 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c182
+ bl_0_182 br_0_182 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c182
+ bl_0_182 br_0_182 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c182
+ bl_0_182 br_0_182 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c182
+ bl_0_182 br_0_182 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c182
+ bl_0_182 br_0_182 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c182
+ bl_0_182 br_0_182 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c182
+ bl_0_182 br_0_182 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c182
+ bl_0_182 br_0_182 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c182
+ bl_0_182 br_0_182 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c182
+ bl_0_182 br_0_182 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c182
+ bl_0_182 br_0_182 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c182
+ bl_0_182 br_0_182 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c182
+ bl_0_182 br_0_182 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c182
+ bl_0_182 br_0_182 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c182
+ bl_0_182 br_0_182 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c182
+ bl_0_182 br_0_182 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c182
+ bl_0_182 br_0_182 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c182
+ bl_0_182 br_0_182 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c182
+ bl_0_182 br_0_182 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c182
+ bl_0_182 br_0_182 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c182
+ bl_0_182 br_0_182 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c182
+ bl_0_182 br_0_182 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c182
+ bl_0_182 br_0_182 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c182
+ bl_0_182 br_0_182 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c182
+ bl_0_182 br_0_182 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c182
+ bl_0_182 br_0_182 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c182
+ bl_0_182 br_0_182 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c182
+ bl_0_182 br_0_182 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c182
+ bl_0_182 br_0_182 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c182
+ bl_0_182 br_0_182 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c182
+ bl_0_182 br_0_182 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c182
+ bl_0_182 br_0_182 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c182
+ bl_0_182 br_0_182 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c182
+ bl_0_182 br_0_182 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c182
+ bl_0_182 br_0_182 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c182
+ bl_0_182 br_0_182 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c182
+ bl_0_182 br_0_182 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c182
+ bl_0_182 br_0_182 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c182
+ bl_0_182 br_0_182 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c182
+ bl_0_182 br_0_182 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c182
+ bl_0_182 br_0_182 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c182
+ bl_0_182 br_0_182 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c183
+ bl_0_183 br_0_183 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c183
+ bl_0_183 br_0_183 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c183
+ bl_0_183 br_0_183 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c183
+ bl_0_183 br_0_183 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c183
+ bl_0_183 br_0_183 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c183
+ bl_0_183 br_0_183 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c183
+ bl_0_183 br_0_183 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c183
+ bl_0_183 br_0_183 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c183
+ bl_0_183 br_0_183 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c183
+ bl_0_183 br_0_183 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c183
+ bl_0_183 br_0_183 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c183
+ bl_0_183 br_0_183 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c183
+ bl_0_183 br_0_183 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c183
+ bl_0_183 br_0_183 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c183
+ bl_0_183 br_0_183 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c183
+ bl_0_183 br_0_183 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c183
+ bl_0_183 br_0_183 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c183
+ bl_0_183 br_0_183 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c183
+ bl_0_183 br_0_183 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c183
+ bl_0_183 br_0_183 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c183
+ bl_0_183 br_0_183 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c183
+ bl_0_183 br_0_183 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c183
+ bl_0_183 br_0_183 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c183
+ bl_0_183 br_0_183 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c183
+ bl_0_183 br_0_183 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c183
+ bl_0_183 br_0_183 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c183
+ bl_0_183 br_0_183 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c183
+ bl_0_183 br_0_183 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c183
+ bl_0_183 br_0_183 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c183
+ bl_0_183 br_0_183 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c183
+ bl_0_183 br_0_183 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c183
+ bl_0_183 br_0_183 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c183
+ bl_0_183 br_0_183 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c183
+ bl_0_183 br_0_183 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c183
+ bl_0_183 br_0_183 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c183
+ bl_0_183 br_0_183 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c183
+ bl_0_183 br_0_183 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c183
+ bl_0_183 br_0_183 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c183
+ bl_0_183 br_0_183 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c183
+ bl_0_183 br_0_183 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c183
+ bl_0_183 br_0_183 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c183
+ bl_0_183 br_0_183 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c183
+ bl_0_183 br_0_183 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c183
+ bl_0_183 br_0_183 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c184
+ bl_0_184 br_0_184 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c184
+ bl_0_184 br_0_184 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c184
+ bl_0_184 br_0_184 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c184
+ bl_0_184 br_0_184 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c184
+ bl_0_184 br_0_184 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c184
+ bl_0_184 br_0_184 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c184
+ bl_0_184 br_0_184 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c184
+ bl_0_184 br_0_184 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c184
+ bl_0_184 br_0_184 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c184
+ bl_0_184 br_0_184 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c184
+ bl_0_184 br_0_184 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c184
+ bl_0_184 br_0_184 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c184
+ bl_0_184 br_0_184 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c184
+ bl_0_184 br_0_184 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c184
+ bl_0_184 br_0_184 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c184
+ bl_0_184 br_0_184 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c184
+ bl_0_184 br_0_184 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c184
+ bl_0_184 br_0_184 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c184
+ bl_0_184 br_0_184 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c184
+ bl_0_184 br_0_184 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c184
+ bl_0_184 br_0_184 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c184
+ bl_0_184 br_0_184 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c184
+ bl_0_184 br_0_184 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c184
+ bl_0_184 br_0_184 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c184
+ bl_0_184 br_0_184 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c184
+ bl_0_184 br_0_184 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c184
+ bl_0_184 br_0_184 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c184
+ bl_0_184 br_0_184 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c184
+ bl_0_184 br_0_184 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c184
+ bl_0_184 br_0_184 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c184
+ bl_0_184 br_0_184 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c184
+ bl_0_184 br_0_184 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c184
+ bl_0_184 br_0_184 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c184
+ bl_0_184 br_0_184 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c184
+ bl_0_184 br_0_184 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c184
+ bl_0_184 br_0_184 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c184
+ bl_0_184 br_0_184 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c184
+ bl_0_184 br_0_184 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c184
+ bl_0_184 br_0_184 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c184
+ bl_0_184 br_0_184 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c184
+ bl_0_184 br_0_184 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c184
+ bl_0_184 br_0_184 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c184
+ bl_0_184 br_0_184 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c184
+ bl_0_184 br_0_184 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c185
+ bl_0_185 br_0_185 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c185
+ bl_0_185 br_0_185 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c185
+ bl_0_185 br_0_185 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c185
+ bl_0_185 br_0_185 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c185
+ bl_0_185 br_0_185 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c185
+ bl_0_185 br_0_185 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c185
+ bl_0_185 br_0_185 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c185
+ bl_0_185 br_0_185 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c185
+ bl_0_185 br_0_185 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c185
+ bl_0_185 br_0_185 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c185
+ bl_0_185 br_0_185 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c185
+ bl_0_185 br_0_185 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c185
+ bl_0_185 br_0_185 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c185
+ bl_0_185 br_0_185 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c185
+ bl_0_185 br_0_185 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c185
+ bl_0_185 br_0_185 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c185
+ bl_0_185 br_0_185 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c185
+ bl_0_185 br_0_185 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c185
+ bl_0_185 br_0_185 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c185
+ bl_0_185 br_0_185 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c185
+ bl_0_185 br_0_185 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c185
+ bl_0_185 br_0_185 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c185
+ bl_0_185 br_0_185 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c185
+ bl_0_185 br_0_185 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c185
+ bl_0_185 br_0_185 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c185
+ bl_0_185 br_0_185 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c185
+ bl_0_185 br_0_185 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c185
+ bl_0_185 br_0_185 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c185
+ bl_0_185 br_0_185 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c185
+ bl_0_185 br_0_185 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c185
+ bl_0_185 br_0_185 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c185
+ bl_0_185 br_0_185 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c185
+ bl_0_185 br_0_185 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c185
+ bl_0_185 br_0_185 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c185
+ bl_0_185 br_0_185 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c185
+ bl_0_185 br_0_185 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c185
+ bl_0_185 br_0_185 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c185
+ bl_0_185 br_0_185 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c185
+ bl_0_185 br_0_185 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c185
+ bl_0_185 br_0_185 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c185
+ bl_0_185 br_0_185 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c185
+ bl_0_185 br_0_185 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c185
+ bl_0_185 br_0_185 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c185
+ bl_0_185 br_0_185 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c186
+ bl_0_186 br_0_186 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c186
+ bl_0_186 br_0_186 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c186
+ bl_0_186 br_0_186 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c186
+ bl_0_186 br_0_186 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c186
+ bl_0_186 br_0_186 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c186
+ bl_0_186 br_0_186 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c186
+ bl_0_186 br_0_186 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c186
+ bl_0_186 br_0_186 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c186
+ bl_0_186 br_0_186 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c186
+ bl_0_186 br_0_186 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c186
+ bl_0_186 br_0_186 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c186
+ bl_0_186 br_0_186 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c186
+ bl_0_186 br_0_186 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c186
+ bl_0_186 br_0_186 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c186
+ bl_0_186 br_0_186 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c186
+ bl_0_186 br_0_186 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c186
+ bl_0_186 br_0_186 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c186
+ bl_0_186 br_0_186 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c186
+ bl_0_186 br_0_186 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c186
+ bl_0_186 br_0_186 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c186
+ bl_0_186 br_0_186 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c186
+ bl_0_186 br_0_186 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c186
+ bl_0_186 br_0_186 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c186
+ bl_0_186 br_0_186 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c186
+ bl_0_186 br_0_186 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c186
+ bl_0_186 br_0_186 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c186
+ bl_0_186 br_0_186 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c186
+ bl_0_186 br_0_186 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c186
+ bl_0_186 br_0_186 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c186
+ bl_0_186 br_0_186 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c186
+ bl_0_186 br_0_186 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c186
+ bl_0_186 br_0_186 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c186
+ bl_0_186 br_0_186 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c186
+ bl_0_186 br_0_186 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c186
+ bl_0_186 br_0_186 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c186
+ bl_0_186 br_0_186 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c186
+ bl_0_186 br_0_186 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c186
+ bl_0_186 br_0_186 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c186
+ bl_0_186 br_0_186 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c186
+ bl_0_186 br_0_186 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c186
+ bl_0_186 br_0_186 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c186
+ bl_0_186 br_0_186 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c186
+ bl_0_186 br_0_186 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c186
+ bl_0_186 br_0_186 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c187
+ bl_0_187 br_0_187 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c187
+ bl_0_187 br_0_187 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c187
+ bl_0_187 br_0_187 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c187
+ bl_0_187 br_0_187 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c187
+ bl_0_187 br_0_187 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c187
+ bl_0_187 br_0_187 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c187
+ bl_0_187 br_0_187 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c187
+ bl_0_187 br_0_187 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c187
+ bl_0_187 br_0_187 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c187
+ bl_0_187 br_0_187 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c187
+ bl_0_187 br_0_187 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c187
+ bl_0_187 br_0_187 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c187
+ bl_0_187 br_0_187 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c187
+ bl_0_187 br_0_187 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c187
+ bl_0_187 br_0_187 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c187
+ bl_0_187 br_0_187 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c187
+ bl_0_187 br_0_187 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c187
+ bl_0_187 br_0_187 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c187
+ bl_0_187 br_0_187 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c187
+ bl_0_187 br_0_187 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c187
+ bl_0_187 br_0_187 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c187
+ bl_0_187 br_0_187 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c187
+ bl_0_187 br_0_187 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c187
+ bl_0_187 br_0_187 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c187
+ bl_0_187 br_0_187 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c187
+ bl_0_187 br_0_187 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c187
+ bl_0_187 br_0_187 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c187
+ bl_0_187 br_0_187 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c187
+ bl_0_187 br_0_187 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c187
+ bl_0_187 br_0_187 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c187
+ bl_0_187 br_0_187 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c187
+ bl_0_187 br_0_187 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c187
+ bl_0_187 br_0_187 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c187
+ bl_0_187 br_0_187 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c187
+ bl_0_187 br_0_187 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c187
+ bl_0_187 br_0_187 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c187
+ bl_0_187 br_0_187 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c187
+ bl_0_187 br_0_187 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c187
+ bl_0_187 br_0_187 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c187
+ bl_0_187 br_0_187 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c187
+ bl_0_187 br_0_187 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c187
+ bl_0_187 br_0_187 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c187
+ bl_0_187 br_0_187 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c187
+ bl_0_187 br_0_187 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c188
+ bl_0_188 br_0_188 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c188
+ bl_0_188 br_0_188 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c188
+ bl_0_188 br_0_188 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c188
+ bl_0_188 br_0_188 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c188
+ bl_0_188 br_0_188 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c188
+ bl_0_188 br_0_188 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c188
+ bl_0_188 br_0_188 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c188
+ bl_0_188 br_0_188 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c188
+ bl_0_188 br_0_188 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c188
+ bl_0_188 br_0_188 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c188
+ bl_0_188 br_0_188 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c188
+ bl_0_188 br_0_188 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c188
+ bl_0_188 br_0_188 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c188
+ bl_0_188 br_0_188 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c188
+ bl_0_188 br_0_188 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c188
+ bl_0_188 br_0_188 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c188
+ bl_0_188 br_0_188 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c188
+ bl_0_188 br_0_188 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c188
+ bl_0_188 br_0_188 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c188
+ bl_0_188 br_0_188 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c188
+ bl_0_188 br_0_188 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c188
+ bl_0_188 br_0_188 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c188
+ bl_0_188 br_0_188 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c188
+ bl_0_188 br_0_188 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c188
+ bl_0_188 br_0_188 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c188
+ bl_0_188 br_0_188 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c188
+ bl_0_188 br_0_188 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c188
+ bl_0_188 br_0_188 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c188
+ bl_0_188 br_0_188 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c188
+ bl_0_188 br_0_188 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c188
+ bl_0_188 br_0_188 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c188
+ bl_0_188 br_0_188 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c188
+ bl_0_188 br_0_188 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c188
+ bl_0_188 br_0_188 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c188
+ bl_0_188 br_0_188 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c188
+ bl_0_188 br_0_188 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c188
+ bl_0_188 br_0_188 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c188
+ bl_0_188 br_0_188 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c188
+ bl_0_188 br_0_188 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c188
+ bl_0_188 br_0_188 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c188
+ bl_0_188 br_0_188 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c188
+ bl_0_188 br_0_188 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c188
+ bl_0_188 br_0_188 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c188
+ bl_0_188 br_0_188 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c189
+ bl_0_189 br_0_189 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c189
+ bl_0_189 br_0_189 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c189
+ bl_0_189 br_0_189 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c189
+ bl_0_189 br_0_189 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c189
+ bl_0_189 br_0_189 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c189
+ bl_0_189 br_0_189 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c189
+ bl_0_189 br_0_189 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c189
+ bl_0_189 br_0_189 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c189
+ bl_0_189 br_0_189 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c189
+ bl_0_189 br_0_189 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c189
+ bl_0_189 br_0_189 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c189
+ bl_0_189 br_0_189 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c189
+ bl_0_189 br_0_189 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c189
+ bl_0_189 br_0_189 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c189
+ bl_0_189 br_0_189 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c189
+ bl_0_189 br_0_189 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c189
+ bl_0_189 br_0_189 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c189
+ bl_0_189 br_0_189 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c189
+ bl_0_189 br_0_189 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c189
+ bl_0_189 br_0_189 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c189
+ bl_0_189 br_0_189 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c189
+ bl_0_189 br_0_189 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c189
+ bl_0_189 br_0_189 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c189
+ bl_0_189 br_0_189 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c189
+ bl_0_189 br_0_189 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c189
+ bl_0_189 br_0_189 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c189
+ bl_0_189 br_0_189 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c189
+ bl_0_189 br_0_189 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c189
+ bl_0_189 br_0_189 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c189
+ bl_0_189 br_0_189 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c189
+ bl_0_189 br_0_189 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c189
+ bl_0_189 br_0_189 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c189
+ bl_0_189 br_0_189 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c189
+ bl_0_189 br_0_189 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c189
+ bl_0_189 br_0_189 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c189
+ bl_0_189 br_0_189 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c189
+ bl_0_189 br_0_189 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c189
+ bl_0_189 br_0_189 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c189
+ bl_0_189 br_0_189 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c189
+ bl_0_189 br_0_189 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c189
+ bl_0_189 br_0_189 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c189
+ bl_0_189 br_0_189 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c189
+ bl_0_189 br_0_189 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c189
+ bl_0_189 br_0_189 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c190
+ bl_0_190 br_0_190 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c190
+ bl_0_190 br_0_190 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c190
+ bl_0_190 br_0_190 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c190
+ bl_0_190 br_0_190 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c190
+ bl_0_190 br_0_190 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c190
+ bl_0_190 br_0_190 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c190
+ bl_0_190 br_0_190 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c190
+ bl_0_190 br_0_190 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c190
+ bl_0_190 br_0_190 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c190
+ bl_0_190 br_0_190 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c190
+ bl_0_190 br_0_190 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c190
+ bl_0_190 br_0_190 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c190
+ bl_0_190 br_0_190 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c190
+ bl_0_190 br_0_190 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c190
+ bl_0_190 br_0_190 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c190
+ bl_0_190 br_0_190 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c190
+ bl_0_190 br_0_190 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c190
+ bl_0_190 br_0_190 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c190
+ bl_0_190 br_0_190 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c190
+ bl_0_190 br_0_190 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c190
+ bl_0_190 br_0_190 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c190
+ bl_0_190 br_0_190 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c190
+ bl_0_190 br_0_190 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c190
+ bl_0_190 br_0_190 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c190
+ bl_0_190 br_0_190 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c190
+ bl_0_190 br_0_190 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c190
+ bl_0_190 br_0_190 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c190
+ bl_0_190 br_0_190 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c190
+ bl_0_190 br_0_190 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c190
+ bl_0_190 br_0_190 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c190
+ bl_0_190 br_0_190 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c190
+ bl_0_190 br_0_190 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c190
+ bl_0_190 br_0_190 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c190
+ bl_0_190 br_0_190 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c190
+ bl_0_190 br_0_190 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c190
+ bl_0_190 br_0_190 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c190
+ bl_0_190 br_0_190 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c190
+ bl_0_190 br_0_190 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c190
+ bl_0_190 br_0_190 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c190
+ bl_0_190 br_0_190 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c190
+ bl_0_190 br_0_190 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c190
+ bl_0_190 br_0_190 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c190
+ bl_0_190 br_0_190 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c190
+ bl_0_190 br_0_190 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c191
+ bl_0_191 br_0_191 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c191
+ bl_0_191 br_0_191 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c191
+ bl_0_191 br_0_191 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c191
+ bl_0_191 br_0_191 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c191
+ bl_0_191 br_0_191 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c191
+ bl_0_191 br_0_191 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c191
+ bl_0_191 br_0_191 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c191
+ bl_0_191 br_0_191 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c191
+ bl_0_191 br_0_191 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c191
+ bl_0_191 br_0_191 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c191
+ bl_0_191 br_0_191 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c191
+ bl_0_191 br_0_191 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c191
+ bl_0_191 br_0_191 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c191
+ bl_0_191 br_0_191 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c191
+ bl_0_191 br_0_191 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c191
+ bl_0_191 br_0_191 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c191
+ bl_0_191 br_0_191 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c191
+ bl_0_191 br_0_191 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c191
+ bl_0_191 br_0_191 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c191
+ bl_0_191 br_0_191 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c191
+ bl_0_191 br_0_191 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c191
+ bl_0_191 br_0_191 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c191
+ bl_0_191 br_0_191 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c191
+ bl_0_191 br_0_191 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c191
+ bl_0_191 br_0_191 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c191
+ bl_0_191 br_0_191 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c191
+ bl_0_191 br_0_191 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c191
+ bl_0_191 br_0_191 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c191
+ bl_0_191 br_0_191 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c191
+ bl_0_191 br_0_191 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c191
+ bl_0_191 br_0_191 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c191
+ bl_0_191 br_0_191 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c191
+ bl_0_191 br_0_191 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c191
+ bl_0_191 br_0_191 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c191
+ bl_0_191 br_0_191 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c191
+ bl_0_191 br_0_191 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c191
+ bl_0_191 br_0_191 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c191
+ bl_0_191 br_0_191 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c191
+ bl_0_191 br_0_191 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c191
+ bl_0_191 br_0_191 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c191
+ bl_0_191 br_0_191 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c191
+ bl_0_191 br_0_191 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c191
+ bl_0_191 br_0_191 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c191
+ bl_0_191 br_0_191 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c192
+ bl_0_192 br_0_192 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c192
+ bl_0_192 br_0_192 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c192
+ bl_0_192 br_0_192 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c192
+ bl_0_192 br_0_192 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c192
+ bl_0_192 br_0_192 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c192
+ bl_0_192 br_0_192 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c192
+ bl_0_192 br_0_192 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c192
+ bl_0_192 br_0_192 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c192
+ bl_0_192 br_0_192 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c192
+ bl_0_192 br_0_192 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c192
+ bl_0_192 br_0_192 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c192
+ bl_0_192 br_0_192 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c192
+ bl_0_192 br_0_192 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c192
+ bl_0_192 br_0_192 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c192
+ bl_0_192 br_0_192 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c192
+ bl_0_192 br_0_192 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c192
+ bl_0_192 br_0_192 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c192
+ bl_0_192 br_0_192 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c192
+ bl_0_192 br_0_192 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c192
+ bl_0_192 br_0_192 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c192
+ bl_0_192 br_0_192 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c192
+ bl_0_192 br_0_192 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c192
+ bl_0_192 br_0_192 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c192
+ bl_0_192 br_0_192 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c192
+ bl_0_192 br_0_192 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c192
+ bl_0_192 br_0_192 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c192
+ bl_0_192 br_0_192 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c192
+ bl_0_192 br_0_192 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c192
+ bl_0_192 br_0_192 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c192
+ bl_0_192 br_0_192 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c192
+ bl_0_192 br_0_192 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c192
+ bl_0_192 br_0_192 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c192
+ bl_0_192 br_0_192 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c192
+ bl_0_192 br_0_192 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c192
+ bl_0_192 br_0_192 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c192
+ bl_0_192 br_0_192 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c192
+ bl_0_192 br_0_192 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c192
+ bl_0_192 br_0_192 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c192
+ bl_0_192 br_0_192 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c192
+ bl_0_192 br_0_192 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c192
+ bl_0_192 br_0_192 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c192
+ bl_0_192 br_0_192 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c192
+ bl_0_192 br_0_192 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c192
+ bl_0_192 br_0_192 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c193
+ bl_0_193 br_0_193 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c193
+ bl_0_193 br_0_193 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c193
+ bl_0_193 br_0_193 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c193
+ bl_0_193 br_0_193 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c193
+ bl_0_193 br_0_193 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c193
+ bl_0_193 br_0_193 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c193
+ bl_0_193 br_0_193 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c193
+ bl_0_193 br_0_193 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c193
+ bl_0_193 br_0_193 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c193
+ bl_0_193 br_0_193 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c193
+ bl_0_193 br_0_193 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c193
+ bl_0_193 br_0_193 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c193
+ bl_0_193 br_0_193 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c193
+ bl_0_193 br_0_193 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c193
+ bl_0_193 br_0_193 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c193
+ bl_0_193 br_0_193 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c193
+ bl_0_193 br_0_193 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c193
+ bl_0_193 br_0_193 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c193
+ bl_0_193 br_0_193 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c193
+ bl_0_193 br_0_193 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c193
+ bl_0_193 br_0_193 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c193
+ bl_0_193 br_0_193 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c193
+ bl_0_193 br_0_193 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c193
+ bl_0_193 br_0_193 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c193
+ bl_0_193 br_0_193 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c193
+ bl_0_193 br_0_193 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c193
+ bl_0_193 br_0_193 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c193
+ bl_0_193 br_0_193 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c193
+ bl_0_193 br_0_193 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c193
+ bl_0_193 br_0_193 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c193
+ bl_0_193 br_0_193 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c193
+ bl_0_193 br_0_193 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c193
+ bl_0_193 br_0_193 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c193
+ bl_0_193 br_0_193 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c193
+ bl_0_193 br_0_193 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c193
+ bl_0_193 br_0_193 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c193
+ bl_0_193 br_0_193 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c193
+ bl_0_193 br_0_193 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c193
+ bl_0_193 br_0_193 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c193
+ bl_0_193 br_0_193 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c193
+ bl_0_193 br_0_193 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c193
+ bl_0_193 br_0_193 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c193
+ bl_0_193 br_0_193 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c193
+ bl_0_193 br_0_193 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c194
+ bl_0_194 br_0_194 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c194
+ bl_0_194 br_0_194 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c194
+ bl_0_194 br_0_194 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c194
+ bl_0_194 br_0_194 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c194
+ bl_0_194 br_0_194 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c194
+ bl_0_194 br_0_194 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c194
+ bl_0_194 br_0_194 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c194
+ bl_0_194 br_0_194 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c194
+ bl_0_194 br_0_194 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c194
+ bl_0_194 br_0_194 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c194
+ bl_0_194 br_0_194 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c194
+ bl_0_194 br_0_194 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c194
+ bl_0_194 br_0_194 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c194
+ bl_0_194 br_0_194 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c194
+ bl_0_194 br_0_194 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c194
+ bl_0_194 br_0_194 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c194
+ bl_0_194 br_0_194 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c194
+ bl_0_194 br_0_194 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c194
+ bl_0_194 br_0_194 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c194
+ bl_0_194 br_0_194 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c194
+ bl_0_194 br_0_194 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c194
+ bl_0_194 br_0_194 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c194
+ bl_0_194 br_0_194 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c194
+ bl_0_194 br_0_194 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c194
+ bl_0_194 br_0_194 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c194
+ bl_0_194 br_0_194 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c194
+ bl_0_194 br_0_194 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c194
+ bl_0_194 br_0_194 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c194
+ bl_0_194 br_0_194 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c194
+ bl_0_194 br_0_194 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c194
+ bl_0_194 br_0_194 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c194
+ bl_0_194 br_0_194 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c194
+ bl_0_194 br_0_194 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c194
+ bl_0_194 br_0_194 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c194
+ bl_0_194 br_0_194 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c194
+ bl_0_194 br_0_194 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c194
+ bl_0_194 br_0_194 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c194
+ bl_0_194 br_0_194 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c194
+ bl_0_194 br_0_194 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c194
+ bl_0_194 br_0_194 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c194
+ bl_0_194 br_0_194 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c194
+ bl_0_194 br_0_194 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c194
+ bl_0_194 br_0_194 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c194
+ bl_0_194 br_0_194 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c195
+ bl_0_195 br_0_195 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c195
+ bl_0_195 br_0_195 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c195
+ bl_0_195 br_0_195 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c195
+ bl_0_195 br_0_195 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c195
+ bl_0_195 br_0_195 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c195
+ bl_0_195 br_0_195 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c195
+ bl_0_195 br_0_195 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c195
+ bl_0_195 br_0_195 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c195
+ bl_0_195 br_0_195 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c195
+ bl_0_195 br_0_195 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c195
+ bl_0_195 br_0_195 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c195
+ bl_0_195 br_0_195 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c195
+ bl_0_195 br_0_195 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c195
+ bl_0_195 br_0_195 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c195
+ bl_0_195 br_0_195 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c195
+ bl_0_195 br_0_195 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c195
+ bl_0_195 br_0_195 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c195
+ bl_0_195 br_0_195 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c195
+ bl_0_195 br_0_195 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c195
+ bl_0_195 br_0_195 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c195
+ bl_0_195 br_0_195 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c195
+ bl_0_195 br_0_195 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c195
+ bl_0_195 br_0_195 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c195
+ bl_0_195 br_0_195 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c195
+ bl_0_195 br_0_195 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c195
+ bl_0_195 br_0_195 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c195
+ bl_0_195 br_0_195 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c195
+ bl_0_195 br_0_195 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c195
+ bl_0_195 br_0_195 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c195
+ bl_0_195 br_0_195 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c195
+ bl_0_195 br_0_195 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c195
+ bl_0_195 br_0_195 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c195
+ bl_0_195 br_0_195 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c195
+ bl_0_195 br_0_195 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c195
+ bl_0_195 br_0_195 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c195
+ bl_0_195 br_0_195 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c195
+ bl_0_195 br_0_195 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c195
+ bl_0_195 br_0_195 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c195
+ bl_0_195 br_0_195 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c195
+ bl_0_195 br_0_195 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c195
+ bl_0_195 br_0_195 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c195
+ bl_0_195 br_0_195 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c195
+ bl_0_195 br_0_195 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c195
+ bl_0_195 br_0_195 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c196
+ bl_0_196 br_0_196 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c196
+ bl_0_196 br_0_196 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c196
+ bl_0_196 br_0_196 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c196
+ bl_0_196 br_0_196 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c196
+ bl_0_196 br_0_196 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c196
+ bl_0_196 br_0_196 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c196
+ bl_0_196 br_0_196 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c196
+ bl_0_196 br_0_196 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c196
+ bl_0_196 br_0_196 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c196
+ bl_0_196 br_0_196 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c196
+ bl_0_196 br_0_196 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c196
+ bl_0_196 br_0_196 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c196
+ bl_0_196 br_0_196 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c196
+ bl_0_196 br_0_196 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c196
+ bl_0_196 br_0_196 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c196
+ bl_0_196 br_0_196 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c196
+ bl_0_196 br_0_196 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c196
+ bl_0_196 br_0_196 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c196
+ bl_0_196 br_0_196 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c196
+ bl_0_196 br_0_196 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c196
+ bl_0_196 br_0_196 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c196
+ bl_0_196 br_0_196 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c196
+ bl_0_196 br_0_196 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c196
+ bl_0_196 br_0_196 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c196
+ bl_0_196 br_0_196 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c196
+ bl_0_196 br_0_196 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c196
+ bl_0_196 br_0_196 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c196
+ bl_0_196 br_0_196 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c196
+ bl_0_196 br_0_196 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c196
+ bl_0_196 br_0_196 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c196
+ bl_0_196 br_0_196 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c196
+ bl_0_196 br_0_196 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c196
+ bl_0_196 br_0_196 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c196
+ bl_0_196 br_0_196 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c196
+ bl_0_196 br_0_196 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c196
+ bl_0_196 br_0_196 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c196
+ bl_0_196 br_0_196 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c196
+ bl_0_196 br_0_196 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c196
+ bl_0_196 br_0_196 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c196
+ bl_0_196 br_0_196 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c196
+ bl_0_196 br_0_196 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c196
+ bl_0_196 br_0_196 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c196
+ bl_0_196 br_0_196 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c196
+ bl_0_196 br_0_196 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c197
+ bl_0_197 br_0_197 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c197
+ bl_0_197 br_0_197 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c197
+ bl_0_197 br_0_197 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c197
+ bl_0_197 br_0_197 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c197
+ bl_0_197 br_0_197 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c197
+ bl_0_197 br_0_197 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c197
+ bl_0_197 br_0_197 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c197
+ bl_0_197 br_0_197 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c197
+ bl_0_197 br_0_197 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c197
+ bl_0_197 br_0_197 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c197
+ bl_0_197 br_0_197 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c197
+ bl_0_197 br_0_197 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c197
+ bl_0_197 br_0_197 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c197
+ bl_0_197 br_0_197 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c197
+ bl_0_197 br_0_197 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c197
+ bl_0_197 br_0_197 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c197
+ bl_0_197 br_0_197 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c197
+ bl_0_197 br_0_197 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c197
+ bl_0_197 br_0_197 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c197
+ bl_0_197 br_0_197 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c197
+ bl_0_197 br_0_197 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c197
+ bl_0_197 br_0_197 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c197
+ bl_0_197 br_0_197 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c197
+ bl_0_197 br_0_197 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c197
+ bl_0_197 br_0_197 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c197
+ bl_0_197 br_0_197 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c197
+ bl_0_197 br_0_197 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c197
+ bl_0_197 br_0_197 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c197
+ bl_0_197 br_0_197 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c197
+ bl_0_197 br_0_197 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c197
+ bl_0_197 br_0_197 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c197
+ bl_0_197 br_0_197 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c197
+ bl_0_197 br_0_197 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c197
+ bl_0_197 br_0_197 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c197
+ bl_0_197 br_0_197 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c197
+ bl_0_197 br_0_197 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c197
+ bl_0_197 br_0_197 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c197
+ bl_0_197 br_0_197 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c197
+ bl_0_197 br_0_197 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c197
+ bl_0_197 br_0_197 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c197
+ bl_0_197 br_0_197 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c197
+ bl_0_197 br_0_197 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c197
+ bl_0_197 br_0_197 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c197
+ bl_0_197 br_0_197 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c198
+ bl_0_198 br_0_198 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c198
+ bl_0_198 br_0_198 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c198
+ bl_0_198 br_0_198 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c198
+ bl_0_198 br_0_198 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c198
+ bl_0_198 br_0_198 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c198
+ bl_0_198 br_0_198 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c198
+ bl_0_198 br_0_198 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c198
+ bl_0_198 br_0_198 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c198
+ bl_0_198 br_0_198 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c198
+ bl_0_198 br_0_198 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c198
+ bl_0_198 br_0_198 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c198
+ bl_0_198 br_0_198 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c198
+ bl_0_198 br_0_198 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c198
+ bl_0_198 br_0_198 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c198
+ bl_0_198 br_0_198 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c198
+ bl_0_198 br_0_198 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c198
+ bl_0_198 br_0_198 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c198
+ bl_0_198 br_0_198 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c198
+ bl_0_198 br_0_198 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c198
+ bl_0_198 br_0_198 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c198
+ bl_0_198 br_0_198 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c198
+ bl_0_198 br_0_198 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c198
+ bl_0_198 br_0_198 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c198
+ bl_0_198 br_0_198 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c198
+ bl_0_198 br_0_198 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c198
+ bl_0_198 br_0_198 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c198
+ bl_0_198 br_0_198 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c198
+ bl_0_198 br_0_198 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c198
+ bl_0_198 br_0_198 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c198
+ bl_0_198 br_0_198 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c198
+ bl_0_198 br_0_198 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c198
+ bl_0_198 br_0_198 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c198
+ bl_0_198 br_0_198 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c198
+ bl_0_198 br_0_198 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c198
+ bl_0_198 br_0_198 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c198
+ bl_0_198 br_0_198 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c198
+ bl_0_198 br_0_198 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c198
+ bl_0_198 br_0_198 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c198
+ bl_0_198 br_0_198 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c198
+ bl_0_198 br_0_198 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c198
+ bl_0_198 br_0_198 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c198
+ bl_0_198 br_0_198 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c198
+ bl_0_198 br_0_198 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c198
+ bl_0_198 br_0_198 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c199
+ bl_0_199 br_0_199 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c199
+ bl_0_199 br_0_199 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c199
+ bl_0_199 br_0_199 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c199
+ bl_0_199 br_0_199 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c199
+ bl_0_199 br_0_199 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c199
+ bl_0_199 br_0_199 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c199
+ bl_0_199 br_0_199 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c199
+ bl_0_199 br_0_199 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c199
+ bl_0_199 br_0_199 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c199
+ bl_0_199 br_0_199 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c199
+ bl_0_199 br_0_199 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c199
+ bl_0_199 br_0_199 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c199
+ bl_0_199 br_0_199 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c199
+ bl_0_199 br_0_199 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c199
+ bl_0_199 br_0_199 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c199
+ bl_0_199 br_0_199 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c199
+ bl_0_199 br_0_199 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c199
+ bl_0_199 br_0_199 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c199
+ bl_0_199 br_0_199 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c199
+ bl_0_199 br_0_199 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c199
+ bl_0_199 br_0_199 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c199
+ bl_0_199 br_0_199 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c199
+ bl_0_199 br_0_199 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c199
+ bl_0_199 br_0_199 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c199
+ bl_0_199 br_0_199 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c199
+ bl_0_199 br_0_199 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c199
+ bl_0_199 br_0_199 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c199
+ bl_0_199 br_0_199 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c199
+ bl_0_199 br_0_199 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c199
+ bl_0_199 br_0_199 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c199
+ bl_0_199 br_0_199 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c199
+ bl_0_199 br_0_199 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c199
+ bl_0_199 br_0_199 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c199
+ bl_0_199 br_0_199 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c199
+ bl_0_199 br_0_199 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c199
+ bl_0_199 br_0_199 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c199
+ bl_0_199 br_0_199 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c199
+ bl_0_199 br_0_199 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c199
+ bl_0_199 br_0_199 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c199
+ bl_0_199 br_0_199 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c199
+ bl_0_199 br_0_199 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c199
+ bl_0_199 br_0_199 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c199
+ bl_0_199 br_0_199 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c199
+ bl_0_199 br_0_199 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c200
+ bl_0_200 br_0_200 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c200
+ bl_0_200 br_0_200 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c200
+ bl_0_200 br_0_200 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c200
+ bl_0_200 br_0_200 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c200
+ bl_0_200 br_0_200 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c200
+ bl_0_200 br_0_200 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c200
+ bl_0_200 br_0_200 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c200
+ bl_0_200 br_0_200 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c200
+ bl_0_200 br_0_200 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c200
+ bl_0_200 br_0_200 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c200
+ bl_0_200 br_0_200 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c200
+ bl_0_200 br_0_200 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c200
+ bl_0_200 br_0_200 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c200
+ bl_0_200 br_0_200 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c200
+ bl_0_200 br_0_200 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c200
+ bl_0_200 br_0_200 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c200
+ bl_0_200 br_0_200 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c200
+ bl_0_200 br_0_200 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c200
+ bl_0_200 br_0_200 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c200
+ bl_0_200 br_0_200 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c200
+ bl_0_200 br_0_200 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c200
+ bl_0_200 br_0_200 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c200
+ bl_0_200 br_0_200 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c200
+ bl_0_200 br_0_200 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c200
+ bl_0_200 br_0_200 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c200
+ bl_0_200 br_0_200 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c200
+ bl_0_200 br_0_200 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c200
+ bl_0_200 br_0_200 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c200
+ bl_0_200 br_0_200 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c200
+ bl_0_200 br_0_200 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c200
+ bl_0_200 br_0_200 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c200
+ bl_0_200 br_0_200 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c200
+ bl_0_200 br_0_200 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c200
+ bl_0_200 br_0_200 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c200
+ bl_0_200 br_0_200 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c200
+ bl_0_200 br_0_200 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c200
+ bl_0_200 br_0_200 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c200
+ bl_0_200 br_0_200 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c200
+ bl_0_200 br_0_200 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c200
+ bl_0_200 br_0_200 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c200
+ bl_0_200 br_0_200 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c200
+ bl_0_200 br_0_200 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c200
+ bl_0_200 br_0_200 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c200
+ bl_0_200 br_0_200 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c201
+ bl_0_201 br_0_201 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c201
+ bl_0_201 br_0_201 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c201
+ bl_0_201 br_0_201 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c201
+ bl_0_201 br_0_201 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c201
+ bl_0_201 br_0_201 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c201
+ bl_0_201 br_0_201 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c201
+ bl_0_201 br_0_201 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c201
+ bl_0_201 br_0_201 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c201
+ bl_0_201 br_0_201 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c201
+ bl_0_201 br_0_201 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c201
+ bl_0_201 br_0_201 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c201
+ bl_0_201 br_0_201 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c201
+ bl_0_201 br_0_201 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c201
+ bl_0_201 br_0_201 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c201
+ bl_0_201 br_0_201 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c201
+ bl_0_201 br_0_201 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c201
+ bl_0_201 br_0_201 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c201
+ bl_0_201 br_0_201 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c201
+ bl_0_201 br_0_201 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c201
+ bl_0_201 br_0_201 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c201
+ bl_0_201 br_0_201 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c201
+ bl_0_201 br_0_201 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c201
+ bl_0_201 br_0_201 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c201
+ bl_0_201 br_0_201 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c201
+ bl_0_201 br_0_201 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c201
+ bl_0_201 br_0_201 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c201
+ bl_0_201 br_0_201 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c201
+ bl_0_201 br_0_201 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c201
+ bl_0_201 br_0_201 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c201
+ bl_0_201 br_0_201 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c201
+ bl_0_201 br_0_201 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c201
+ bl_0_201 br_0_201 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c201
+ bl_0_201 br_0_201 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c201
+ bl_0_201 br_0_201 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c201
+ bl_0_201 br_0_201 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c201
+ bl_0_201 br_0_201 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c201
+ bl_0_201 br_0_201 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c201
+ bl_0_201 br_0_201 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c201
+ bl_0_201 br_0_201 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c201
+ bl_0_201 br_0_201 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c201
+ bl_0_201 br_0_201 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c201
+ bl_0_201 br_0_201 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c201
+ bl_0_201 br_0_201 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c201
+ bl_0_201 br_0_201 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c202
+ bl_0_202 br_0_202 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c202
+ bl_0_202 br_0_202 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c202
+ bl_0_202 br_0_202 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c202
+ bl_0_202 br_0_202 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c202
+ bl_0_202 br_0_202 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c202
+ bl_0_202 br_0_202 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c202
+ bl_0_202 br_0_202 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c202
+ bl_0_202 br_0_202 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c202
+ bl_0_202 br_0_202 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c202
+ bl_0_202 br_0_202 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c202
+ bl_0_202 br_0_202 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c202
+ bl_0_202 br_0_202 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c202
+ bl_0_202 br_0_202 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c202
+ bl_0_202 br_0_202 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c202
+ bl_0_202 br_0_202 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c202
+ bl_0_202 br_0_202 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c202
+ bl_0_202 br_0_202 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c202
+ bl_0_202 br_0_202 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c202
+ bl_0_202 br_0_202 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c202
+ bl_0_202 br_0_202 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c202
+ bl_0_202 br_0_202 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c202
+ bl_0_202 br_0_202 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c202
+ bl_0_202 br_0_202 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c202
+ bl_0_202 br_0_202 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c202
+ bl_0_202 br_0_202 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c202
+ bl_0_202 br_0_202 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c202
+ bl_0_202 br_0_202 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c202
+ bl_0_202 br_0_202 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c202
+ bl_0_202 br_0_202 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c202
+ bl_0_202 br_0_202 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c202
+ bl_0_202 br_0_202 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c202
+ bl_0_202 br_0_202 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c202
+ bl_0_202 br_0_202 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c202
+ bl_0_202 br_0_202 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c202
+ bl_0_202 br_0_202 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c202
+ bl_0_202 br_0_202 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c202
+ bl_0_202 br_0_202 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c202
+ bl_0_202 br_0_202 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c202
+ bl_0_202 br_0_202 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c202
+ bl_0_202 br_0_202 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c202
+ bl_0_202 br_0_202 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c202
+ bl_0_202 br_0_202 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c202
+ bl_0_202 br_0_202 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c202
+ bl_0_202 br_0_202 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c203
+ bl_0_203 br_0_203 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c203
+ bl_0_203 br_0_203 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c203
+ bl_0_203 br_0_203 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c203
+ bl_0_203 br_0_203 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c203
+ bl_0_203 br_0_203 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c203
+ bl_0_203 br_0_203 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c203
+ bl_0_203 br_0_203 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c203
+ bl_0_203 br_0_203 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c203
+ bl_0_203 br_0_203 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c203
+ bl_0_203 br_0_203 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c203
+ bl_0_203 br_0_203 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c203
+ bl_0_203 br_0_203 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c203
+ bl_0_203 br_0_203 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c203
+ bl_0_203 br_0_203 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c203
+ bl_0_203 br_0_203 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c203
+ bl_0_203 br_0_203 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c203
+ bl_0_203 br_0_203 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c203
+ bl_0_203 br_0_203 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c203
+ bl_0_203 br_0_203 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c203
+ bl_0_203 br_0_203 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c203
+ bl_0_203 br_0_203 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c203
+ bl_0_203 br_0_203 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c203
+ bl_0_203 br_0_203 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c203
+ bl_0_203 br_0_203 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c203
+ bl_0_203 br_0_203 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c203
+ bl_0_203 br_0_203 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c203
+ bl_0_203 br_0_203 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c203
+ bl_0_203 br_0_203 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c203
+ bl_0_203 br_0_203 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c203
+ bl_0_203 br_0_203 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c203
+ bl_0_203 br_0_203 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c203
+ bl_0_203 br_0_203 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c203
+ bl_0_203 br_0_203 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c203
+ bl_0_203 br_0_203 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c203
+ bl_0_203 br_0_203 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c203
+ bl_0_203 br_0_203 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c203
+ bl_0_203 br_0_203 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c203
+ bl_0_203 br_0_203 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c203
+ bl_0_203 br_0_203 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c203
+ bl_0_203 br_0_203 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c203
+ bl_0_203 br_0_203 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c203
+ bl_0_203 br_0_203 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c203
+ bl_0_203 br_0_203 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c203
+ bl_0_203 br_0_203 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c204
+ bl_0_204 br_0_204 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c204
+ bl_0_204 br_0_204 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c204
+ bl_0_204 br_0_204 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c204
+ bl_0_204 br_0_204 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c204
+ bl_0_204 br_0_204 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c204
+ bl_0_204 br_0_204 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c204
+ bl_0_204 br_0_204 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c204
+ bl_0_204 br_0_204 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c204
+ bl_0_204 br_0_204 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c204
+ bl_0_204 br_0_204 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c204
+ bl_0_204 br_0_204 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c204
+ bl_0_204 br_0_204 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c204
+ bl_0_204 br_0_204 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c204
+ bl_0_204 br_0_204 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c204
+ bl_0_204 br_0_204 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c204
+ bl_0_204 br_0_204 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c204
+ bl_0_204 br_0_204 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c204
+ bl_0_204 br_0_204 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c204
+ bl_0_204 br_0_204 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c204
+ bl_0_204 br_0_204 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c204
+ bl_0_204 br_0_204 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c204
+ bl_0_204 br_0_204 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c204
+ bl_0_204 br_0_204 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c204
+ bl_0_204 br_0_204 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c204
+ bl_0_204 br_0_204 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c204
+ bl_0_204 br_0_204 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c204
+ bl_0_204 br_0_204 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c204
+ bl_0_204 br_0_204 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c204
+ bl_0_204 br_0_204 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c204
+ bl_0_204 br_0_204 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c204
+ bl_0_204 br_0_204 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c204
+ bl_0_204 br_0_204 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c204
+ bl_0_204 br_0_204 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c204
+ bl_0_204 br_0_204 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c204
+ bl_0_204 br_0_204 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c204
+ bl_0_204 br_0_204 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c204
+ bl_0_204 br_0_204 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c204
+ bl_0_204 br_0_204 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c204
+ bl_0_204 br_0_204 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c204
+ bl_0_204 br_0_204 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c204
+ bl_0_204 br_0_204 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c204
+ bl_0_204 br_0_204 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c204
+ bl_0_204 br_0_204 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c204
+ bl_0_204 br_0_204 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c205
+ bl_0_205 br_0_205 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c205
+ bl_0_205 br_0_205 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c205
+ bl_0_205 br_0_205 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c205
+ bl_0_205 br_0_205 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c205
+ bl_0_205 br_0_205 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c205
+ bl_0_205 br_0_205 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c205
+ bl_0_205 br_0_205 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c205
+ bl_0_205 br_0_205 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c205
+ bl_0_205 br_0_205 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c205
+ bl_0_205 br_0_205 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c205
+ bl_0_205 br_0_205 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c205
+ bl_0_205 br_0_205 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c205
+ bl_0_205 br_0_205 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c205
+ bl_0_205 br_0_205 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c205
+ bl_0_205 br_0_205 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c205
+ bl_0_205 br_0_205 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c205
+ bl_0_205 br_0_205 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c205
+ bl_0_205 br_0_205 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c205
+ bl_0_205 br_0_205 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c205
+ bl_0_205 br_0_205 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c205
+ bl_0_205 br_0_205 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c205
+ bl_0_205 br_0_205 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c205
+ bl_0_205 br_0_205 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c205
+ bl_0_205 br_0_205 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c205
+ bl_0_205 br_0_205 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c205
+ bl_0_205 br_0_205 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c205
+ bl_0_205 br_0_205 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c205
+ bl_0_205 br_0_205 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c205
+ bl_0_205 br_0_205 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c205
+ bl_0_205 br_0_205 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c205
+ bl_0_205 br_0_205 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c205
+ bl_0_205 br_0_205 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c205
+ bl_0_205 br_0_205 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c205
+ bl_0_205 br_0_205 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c205
+ bl_0_205 br_0_205 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c205
+ bl_0_205 br_0_205 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c205
+ bl_0_205 br_0_205 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c205
+ bl_0_205 br_0_205 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c205
+ bl_0_205 br_0_205 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c205
+ bl_0_205 br_0_205 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c205
+ bl_0_205 br_0_205 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c205
+ bl_0_205 br_0_205 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c205
+ bl_0_205 br_0_205 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c205
+ bl_0_205 br_0_205 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c206
+ bl_0_206 br_0_206 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c206
+ bl_0_206 br_0_206 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c206
+ bl_0_206 br_0_206 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c206
+ bl_0_206 br_0_206 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c206
+ bl_0_206 br_0_206 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c206
+ bl_0_206 br_0_206 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c206
+ bl_0_206 br_0_206 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c206
+ bl_0_206 br_0_206 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c206
+ bl_0_206 br_0_206 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c206
+ bl_0_206 br_0_206 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c206
+ bl_0_206 br_0_206 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c206
+ bl_0_206 br_0_206 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c206
+ bl_0_206 br_0_206 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c206
+ bl_0_206 br_0_206 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c206
+ bl_0_206 br_0_206 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c206
+ bl_0_206 br_0_206 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c206
+ bl_0_206 br_0_206 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c206
+ bl_0_206 br_0_206 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c206
+ bl_0_206 br_0_206 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c206
+ bl_0_206 br_0_206 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c206
+ bl_0_206 br_0_206 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c206
+ bl_0_206 br_0_206 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c206
+ bl_0_206 br_0_206 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c206
+ bl_0_206 br_0_206 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c206
+ bl_0_206 br_0_206 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c206
+ bl_0_206 br_0_206 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c206
+ bl_0_206 br_0_206 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c206
+ bl_0_206 br_0_206 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c206
+ bl_0_206 br_0_206 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c206
+ bl_0_206 br_0_206 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c206
+ bl_0_206 br_0_206 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c206
+ bl_0_206 br_0_206 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c206
+ bl_0_206 br_0_206 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c206
+ bl_0_206 br_0_206 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c206
+ bl_0_206 br_0_206 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c206
+ bl_0_206 br_0_206 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c206
+ bl_0_206 br_0_206 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c206
+ bl_0_206 br_0_206 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c206
+ bl_0_206 br_0_206 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c206
+ bl_0_206 br_0_206 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c206
+ bl_0_206 br_0_206 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c206
+ bl_0_206 br_0_206 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c206
+ bl_0_206 br_0_206 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c206
+ bl_0_206 br_0_206 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c207
+ bl_0_207 br_0_207 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c207
+ bl_0_207 br_0_207 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c207
+ bl_0_207 br_0_207 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c207
+ bl_0_207 br_0_207 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c207
+ bl_0_207 br_0_207 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c207
+ bl_0_207 br_0_207 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c207
+ bl_0_207 br_0_207 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c207
+ bl_0_207 br_0_207 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c207
+ bl_0_207 br_0_207 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c207
+ bl_0_207 br_0_207 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c207
+ bl_0_207 br_0_207 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c207
+ bl_0_207 br_0_207 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c207
+ bl_0_207 br_0_207 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c207
+ bl_0_207 br_0_207 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c207
+ bl_0_207 br_0_207 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c207
+ bl_0_207 br_0_207 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c207
+ bl_0_207 br_0_207 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c207
+ bl_0_207 br_0_207 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c207
+ bl_0_207 br_0_207 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c207
+ bl_0_207 br_0_207 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c207
+ bl_0_207 br_0_207 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c207
+ bl_0_207 br_0_207 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c207
+ bl_0_207 br_0_207 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c207
+ bl_0_207 br_0_207 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c207
+ bl_0_207 br_0_207 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c207
+ bl_0_207 br_0_207 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c207
+ bl_0_207 br_0_207 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c207
+ bl_0_207 br_0_207 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c207
+ bl_0_207 br_0_207 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c207
+ bl_0_207 br_0_207 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c207
+ bl_0_207 br_0_207 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c207
+ bl_0_207 br_0_207 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c207
+ bl_0_207 br_0_207 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c207
+ bl_0_207 br_0_207 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c207
+ bl_0_207 br_0_207 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c207
+ bl_0_207 br_0_207 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c207
+ bl_0_207 br_0_207 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c207
+ bl_0_207 br_0_207 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c207
+ bl_0_207 br_0_207 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c207
+ bl_0_207 br_0_207 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c207
+ bl_0_207 br_0_207 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c207
+ bl_0_207 br_0_207 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c207
+ bl_0_207 br_0_207 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c207
+ bl_0_207 br_0_207 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c208
+ bl_0_208 br_0_208 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c208
+ bl_0_208 br_0_208 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c208
+ bl_0_208 br_0_208 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c208
+ bl_0_208 br_0_208 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c208
+ bl_0_208 br_0_208 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c208
+ bl_0_208 br_0_208 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c208
+ bl_0_208 br_0_208 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c208
+ bl_0_208 br_0_208 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c208
+ bl_0_208 br_0_208 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c208
+ bl_0_208 br_0_208 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c208
+ bl_0_208 br_0_208 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c208
+ bl_0_208 br_0_208 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c208
+ bl_0_208 br_0_208 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c208
+ bl_0_208 br_0_208 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c208
+ bl_0_208 br_0_208 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c208
+ bl_0_208 br_0_208 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c208
+ bl_0_208 br_0_208 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c208
+ bl_0_208 br_0_208 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c208
+ bl_0_208 br_0_208 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c208
+ bl_0_208 br_0_208 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c208
+ bl_0_208 br_0_208 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c208
+ bl_0_208 br_0_208 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c208
+ bl_0_208 br_0_208 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c208
+ bl_0_208 br_0_208 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c208
+ bl_0_208 br_0_208 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c208
+ bl_0_208 br_0_208 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c208
+ bl_0_208 br_0_208 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c208
+ bl_0_208 br_0_208 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c208
+ bl_0_208 br_0_208 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c208
+ bl_0_208 br_0_208 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c208
+ bl_0_208 br_0_208 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c208
+ bl_0_208 br_0_208 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c208
+ bl_0_208 br_0_208 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c208
+ bl_0_208 br_0_208 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c208
+ bl_0_208 br_0_208 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c208
+ bl_0_208 br_0_208 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c208
+ bl_0_208 br_0_208 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c208
+ bl_0_208 br_0_208 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c208
+ bl_0_208 br_0_208 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c208
+ bl_0_208 br_0_208 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c208
+ bl_0_208 br_0_208 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c208
+ bl_0_208 br_0_208 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c208
+ bl_0_208 br_0_208 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c208
+ bl_0_208 br_0_208 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c209
+ bl_0_209 br_0_209 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c209
+ bl_0_209 br_0_209 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c209
+ bl_0_209 br_0_209 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c209
+ bl_0_209 br_0_209 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c209
+ bl_0_209 br_0_209 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c209
+ bl_0_209 br_0_209 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c209
+ bl_0_209 br_0_209 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c209
+ bl_0_209 br_0_209 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c209
+ bl_0_209 br_0_209 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c209
+ bl_0_209 br_0_209 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c209
+ bl_0_209 br_0_209 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c209
+ bl_0_209 br_0_209 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c209
+ bl_0_209 br_0_209 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c209
+ bl_0_209 br_0_209 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c209
+ bl_0_209 br_0_209 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c209
+ bl_0_209 br_0_209 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c209
+ bl_0_209 br_0_209 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c209
+ bl_0_209 br_0_209 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c209
+ bl_0_209 br_0_209 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c209
+ bl_0_209 br_0_209 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c209
+ bl_0_209 br_0_209 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c209
+ bl_0_209 br_0_209 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c209
+ bl_0_209 br_0_209 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c209
+ bl_0_209 br_0_209 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c209
+ bl_0_209 br_0_209 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c209
+ bl_0_209 br_0_209 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c209
+ bl_0_209 br_0_209 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c209
+ bl_0_209 br_0_209 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c209
+ bl_0_209 br_0_209 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c209
+ bl_0_209 br_0_209 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c209
+ bl_0_209 br_0_209 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c209
+ bl_0_209 br_0_209 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c209
+ bl_0_209 br_0_209 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c209
+ bl_0_209 br_0_209 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c209
+ bl_0_209 br_0_209 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c209
+ bl_0_209 br_0_209 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c209
+ bl_0_209 br_0_209 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c209
+ bl_0_209 br_0_209 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c209
+ bl_0_209 br_0_209 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c209
+ bl_0_209 br_0_209 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c209
+ bl_0_209 br_0_209 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c209
+ bl_0_209 br_0_209 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c209
+ bl_0_209 br_0_209 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c209
+ bl_0_209 br_0_209 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c210
+ bl_0_210 br_0_210 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c210
+ bl_0_210 br_0_210 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c210
+ bl_0_210 br_0_210 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c210
+ bl_0_210 br_0_210 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c210
+ bl_0_210 br_0_210 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c210
+ bl_0_210 br_0_210 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c210
+ bl_0_210 br_0_210 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c210
+ bl_0_210 br_0_210 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c210
+ bl_0_210 br_0_210 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c210
+ bl_0_210 br_0_210 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c210
+ bl_0_210 br_0_210 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c210
+ bl_0_210 br_0_210 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c210
+ bl_0_210 br_0_210 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c210
+ bl_0_210 br_0_210 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c210
+ bl_0_210 br_0_210 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c210
+ bl_0_210 br_0_210 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c210
+ bl_0_210 br_0_210 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c210
+ bl_0_210 br_0_210 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c210
+ bl_0_210 br_0_210 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c210
+ bl_0_210 br_0_210 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c210
+ bl_0_210 br_0_210 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c210
+ bl_0_210 br_0_210 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c210
+ bl_0_210 br_0_210 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c210
+ bl_0_210 br_0_210 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c210
+ bl_0_210 br_0_210 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c210
+ bl_0_210 br_0_210 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c210
+ bl_0_210 br_0_210 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c210
+ bl_0_210 br_0_210 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c210
+ bl_0_210 br_0_210 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c210
+ bl_0_210 br_0_210 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c210
+ bl_0_210 br_0_210 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c210
+ bl_0_210 br_0_210 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c210
+ bl_0_210 br_0_210 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c210
+ bl_0_210 br_0_210 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c210
+ bl_0_210 br_0_210 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c210
+ bl_0_210 br_0_210 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c210
+ bl_0_210 br_0_210 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c210
+ bl_0_210 br_0_210 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c210
+ bl_0_210 br_0_210 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c210
+ bl_0_210 br_0_210 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c210
+ bl_0_210 br_0_210 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c210
+ bl_0_210 br_0_210 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c210
+ bl_0_210 br_0_210 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c210
+ bl_0_210 br_0_210 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c211
+ bl_0_211 br_0_211 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c211
+ bl_0_211 br_0_211 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c211
+ bl_0_211 br_0_211 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c211
+ bl_0_211 br_0_211 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c211
+ bl_0_211 br_0_211 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c211
+ bl_0_211 br_0_211 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c211
+ bl_0_211 br_0_211 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c211
+ bl_0_211 br_0_211 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c211
+ bl_0_211 br_0_211 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c211
+ bl_0_211 br_0_211 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c211
+ bl_0_211 br_0_211 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c211
+ bl_0_211 br_0_211 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c211
+ bl_0_211 br_0_211 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c211
+ bl_0_211 br_0_211 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c211
+ bl_0_211 br_0_211 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c211
+ bl_0_211 br_0_211 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c211
+ bl_0_211 br_0_211 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c211
+ bl_0_211 br_0_211 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c211
+ bl_0_211 br_0_211 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c211
+ bl_0_211 br_0_211 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c211
+ bl_0_211 br_0_211 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c211
+ bl_0_211 br_0_211 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c211
+ bl_0_211 br_0_211 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c211
+ bl_0_211 br_0_211 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c211
+ bl_0_211 br_0_211 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c211
+ bl_0_211 br_0_211 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c211
+ bl_0_211 br_0_211 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c211
+ bl_0_211 br_0_211 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c211
+ bl_0_211 br_0_211 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c211
+ bl_0_211 br_0_211 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c211
+ bl_0_211 br_0_211 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c211
+ bl_0_211 br_0_211 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c211
+ bl_0_211 br_0_211 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c211
+ bl_0_211 br_0_211 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c211
+ bl_0_211 br_0_211 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c211
+ bl_0_211 br_0_211 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c211
+ bl_0_211 br_0_211 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c211
+ bl_0_211 br_0_211 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c211
+ bl_0_211 br_0_211 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c211
+ bl_0_211 br_0_211 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c211
+ bl_0_211 br_0_211 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c211
+ bl_0_211 br_0_211 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c211
+ bl_0_211 br_0_211 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c211
+ bl_0_211 br_0_211 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c212
+ bl_0_212 br_0_212 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c212
+ bl_0_212 br_0_212 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c212
+ bl_0_212 br_0_212 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c212
+ bl_0_212 br_0_212 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c212
+ bl_0_212 br_0_212 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c212
+ bl_0_212 br_0_212 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c212
+ bl_0_212 br_0_212 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c212
+ bl_0_212 br_0_212 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c212
+ bl_0_212 br_0_212 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c212
+ bl_0_212 br_0_212 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c212
+ bl_0_212 br_0_212 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c212
+ bl_0_212 br_0_212 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c212
+ bl_0_212 br_0_212 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c212
+ bl_0_212 br_0_212 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c212
+ bl_0_212 br_0_212 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c212
+ bl_0_212 br_0_212 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c212
+ bl_0_212 br_0_212 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c212
+ bl_0_212 br_0_212 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c212
+ bl_0_212 br_0_212 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c212
+ bl_0_212 br_0_212 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c212
+ bl_0_212 br_0_212 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c212
+ bl_0_212 br_0_212 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c212
+ bl_0_212 br_0_212 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c212
+ bl_0_212 br_0_212 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c212
+ bl_0_212 br_0_212 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c212
+ bl_0_212 br_0_212 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c212
+ bl_0_212 br_0_212 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c212
+ bl_0_212 br_0_212 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c212
+ bl_0_212 br_0_212 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c212
+ bl_0_212 br_0_212 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c212
+ bl_0_212 br_0_212 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c212
+ bl_0_212 br_0_212 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c212
+ bl_0_212 br_0_212 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c212
+ bl_0_212 br_0_212 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c212
+ bl_0_212 br_0_212 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c212
+ bl_0_212 br_0_212 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c212
+ bl_0_212 br_0_212 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c212
+ bl_0_212 br_0_212 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c212
+ bl_0_212 br_0_212 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c212
+ bl_0_212 br_0_212 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c212
+ bl_0_212 br_0_212 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c212
+ bl_0_212 br_0_212 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c212
+ bl_0_212 br_0_212 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c212
+ bl_0_212 br_0_212 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c213
+ bl_0_213 br_0_213 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c213
+ bl_0_213 br_0_213 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c213
+ bl_0_213 br_0_213 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c213
+ bl_0_213 br_0_213 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c213
+ bl_0_213 br_0_213 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c213
+ bl_0_213 br_0_213 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c213
+ bl_0_213 br_0_213 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c213
+ bl_0_213 br_0_213 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c213
+ bl_0_213 br_0_213 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c213
+ bl_0_213 br_0_213 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c213
+ bl_0_213 br_0_213 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c213
+ bl_0_213 br_0_213 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c213
+ bl_0_213 br_0_213 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c213
+ bl_0_213 br_0_213 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c213
+ bl_0_213 br_0_213 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c213
+ bl_0_213 br_0_213 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c213
+ bl_0_213 br_0_213 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c213
+ bl_0_213 br_0_213 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c213
+ bl_0_213 br_0_213 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c213
+ bl_0_213 br_0_213 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c213
+ bl_0_213 br_0_213 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c213
+ bl_0_213 br_0_213 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c213
+ bl_0_213 br_0_213 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c213
+ bl_0_213 br_0_213 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c213
+ bl_0_213 br_0_213 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c213
+ bl_0_213 br_0_213 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c213
+ bl_0_213 br_0_213 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c213
+ bl_0_213 br_0_213 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c213
+ bl_0_213 br_0_213 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c213
+ bl_0_213 br_0_213 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c213
+ bl_0_213 br_0_213 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c213
+ bl_0_213 br_0_213 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c213
+ bl_0_213 br_0_213 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c213
+ bl_0_213 br_0_213 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c213
+ bl_0_213 br_0_213 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c213
+ bl_0_213 br_0_213 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c213
+ bl_0_213 br_0_213 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c213
+ bl_0_213 br_0_213 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c213
+ bl_0_213 br_0_213 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c213
+ bl_0_213 br_0_213 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c213
+ bl_0_213 br_0_213 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c213
+ bl_0_213 br_0_213 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c213
+ bl_0_213 br_0_213 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c213
+ bl_0_213 br_0_213 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c214
+ bl_0_214 br_0_214 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c214
+ bl_0_214 br_0_214 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c214
+ bl_0_214 br_0_214 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c214
+ bl_0_214 br_0_214 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c214
+ bl_0_214 br_0_214 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c214
+ bl_0_214 br_0_214 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c214
+ bl_0_214 br_0_214 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c214
+ bl_0_214 br_0_214 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c214
+ bl_0_214 br_0_214 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c214
+ bl_0_214 br_0_214 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c214
+ bl_0_214 br_0_214 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c214
+ bl_0_214 br_0_214 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c214
+ bl_0_214 br_0_214 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c214
+ bl_0_214 br_0_214 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c214
+ bl_0_214 br_0_214 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c214
+ bl_0_214 br_0_214 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c214
+ bl_0_214 br_0_214 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c214
+ bl_0_214 br_0_214 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c214
+ bl_0_214 br_0_214 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c214
+ bl_0_214 br_0_214 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c214
+ bl_0_214 br_0_214 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c214
+ bl_0_214 br_0_214 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c214
+ bl_0_214 br_0_214 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c214
+ bl_0_214 br_0_214 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c214
+ bl_0_214 br_0_214 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c214
+ bl_0_214 br_0_214 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c214
+ bl_0_214 br_0_214 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c214
+ bl_0_214 br_0_214 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c214
+ bl_0_214 br_0_214 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c214
+ bl_0_214 br_0_214 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c214
+ bl_0_214 br_0_214 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c214
+ bl_0_214 br_0_214 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c214
+ bl_0_214 br_0_214 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c214
+ bl_0_214 br_0_214 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c214
+ bl_0_214 br_0_214 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c214
+ bl_0_214 br_0_214 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c214
+ bl_0_214 br_0_214 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c214
+ bl_0_214 br_0_214 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c214
+ bl_0_214 br_0_214 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c214
+ bl_0_214 br_0_214 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c214
+ bl_0_214 br_0_214 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c214
+ bl_0_214 br_0_214 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c214
+ bl_0_214 br_0_214 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c214
+ bl_0_214 br_0_214 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c215
+ bl_0_215 br_0_215 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c215
+ bl_0_215 br_0_215 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c215
+ bl_0_215 br_0_215 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c215
+ bl_0_215 br_0_215 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c215
+ bl_0_215 br_0_215 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c215
+ bl_0_215 br_0_215 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c215
+ bl_0_215 br_0_215 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c215
+ bl_0_215 br_0_215 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c215
+ bl_0_215 br_0_215 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c215
+ bl_0_215 br_0_215 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c215
+ bl_0_215 br_0_215 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c215
+ bl_0_215 br_0_215 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c215
+ bl_0_215 br_0_215 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c215
+ bl_0_215 br_0_215 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c215
+ bl_0_215 br_0_215 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c215
+ bl_0_215 br_0_215 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c215
+ bl_0_215 br_0_215 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c215
+ bl_0_215 br_0_215 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c215
+ bl_0_215 br_0_215 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c215
+ bl_0_215 br_0_215 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c215
+ bl_0_215 br_0_215 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c215
+ bl_0_215 br_0_215 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c215
+ bl_0_215 br_0_215 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c215
+ bl_0_215 br_0_215 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c215
+ bl_0_215 br_0_215 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c215
+ bl_0_215 br_0_215 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c215
+ bl_0_215 br_0_215 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c215
+ bl_0_215 br_0_215 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c215
+ bl_0_215 br_0_215 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c215
+ bl_0_215 br_0_215 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c215
+ bl_0_215 br_0_215 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c215
+ bl_0_215 br_0_215 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c215
+ bl_0_215 br_0_215 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c215
+ bl_0_215 br_0_215 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c215
+ bl_0_215 br_0_215 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c215
+ bl_0_215 br_0_215 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c215
+ bl_0_215 br_0_215 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c215
+ bl_0_215 br_0_215 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c215
+ bl_0_215 br_0_215 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c215
+ bl_0_215 br_0_215 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c215
+ bl_0_215 br_0_215 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c215
+ bl_0_215 br_0_215 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c215
+ bl_0_215 br_0_215 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c215
+ bl_0_215 br_0_215 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c216
+ bl_0_216 br_0_216 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c216
+ bl_0_216 br_0_216 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c216
+ bl_0_216 br_0_216 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c216
+ bl_0_216 br_0_216 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c216
+ bl_0_216 br_0_216 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c216
+ bl_0_216 br_0_216 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c216
+ bl_0_216 br_0_216 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c216
+ bl_0_216 br_0_216 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c216
+ bl_0_216 br_0_216 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c216
+ bl_0_216 br_0_216 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c216
+ bl_0_216 br_0_216 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c216
+ bl_0_216 br_0_216 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c216
+ bl_0_216 br_0_216 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c216
+ bl_0_216 br_0_216 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c216
+ bl_0_216 br_0_216 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c216
+ bl_0_216 br_0_216 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c216
+ bl_0_216 br_0_216 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c216
+ bl_0_216 br_0_216 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c216
+ bl_0_216 br_0_216 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c216
+ bl_0_216 br_0_216 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c216
+ bl_0_216 br_0_216 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c216
+ bl_0_216 br_0_216 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c216
+ bl_0_216 br_0_216 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c216
+ bl_0_216 br_0_216 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c216
+ bl_0_216 br_0_216 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c216
+ bl_0_216 br_0_216 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c216
+ bl_0_216 br_0_216 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c216
+ bl_0_216 br_0_216 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c216
+ bl_0_216 br_0_216 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c216
+ bl_0_216 br_0_216 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c216
+ bl_0_216 br_0_216 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c216
+ bl_0_216 br_0_216 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c216
+ bl_0_216 br_0_216 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c216
+ bl_0_216 br_0_216 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c216
+ bl_0_216 br_0_216 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c216
+ bl_0_216 br_0_216 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c216
+ bl_0_216 br_0_216 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c216
+ bl_0_216 br_0_216 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c216
+ bl_0_216 br_0_216 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c216
+ bl_0_216 br_0_216 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c216
+ bl_0_216 br_0_216 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c216
+ bl_0_216 br_0_216 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c216
+ bl_0_216 br_0_216 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c216
+ bl_0_216 br_0_216 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c217
+ bl_0_217 br_0_217 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c217
+ bl_0_217 br_0_217 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c217
+ bl_0_217 br_0_217 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c217
+ bl_0_217 br_0_217 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c217
+ bl_0_217 br_0_217 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c217
+ bl_0_217 br_0_217 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c217
+ bl_0_217 br_0_217 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c217
+ bl_0_217 br_0_217 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c217
+ bl_0_217 br_0_217 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c217
+ bl_0_217 br_0_217 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c217
+ bl_0_217 br_0_217 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c217
+ bl_0_217 br_0_217 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c217
+ bl_0_217 br_0_217 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c217
+ bl_0_217 br_0_217 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c217
+ bl_0_217 br_0_217 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c217
+ bl_0_217 br_0_217 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c217
+ bl_0_217 br_0_217 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c217
+ bl_0_217 br_0_217 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c217
+ bl_0_217 br_0_217 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c217
+ bl_0_217 br_0_217 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c217
+ bl_0_217 br_0_217 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c217
+ bl_0_217 br_0_217 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c217
+ bl_0_217 br_0_217 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c217
+ bl_0_217 br_0_217 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c217
+ bl_0_217 br_0_217 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c217
+ bl_0_217 br_0_217 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c217
+ bl_0_217 br_0_217 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c217
+ bl_0_217 br_0_217 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c217
+ bl_0_217 br_0_217 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c217
+ bl_0_217 br_0_217 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c217
+ bl_0_217 br_0_217 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c217
+ bl_0_217 br_0_217 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c217
+ bl_0_217 br_0_217 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c217
+ bl_0_217 br_0_217 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c217
+ bl_0_217 br_0_217 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c217
+ bl_0_217 br_0_217 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c217
+ bl_0_217 br_0_217 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c217
+ bl_0_217 br_0_217 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c217
+ bl_0_217 br_0_217 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c217
+ bl_0_217 br_0_217 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c217
+ bl_0_217 br_0_217 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c217
+ bl_0_217 br_0_217 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c217
+ bl_0_217 br_0_217 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c217
+ bl_0_217 br_0_217 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c218
+ bl_0_218 br_0_218 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c218
+ bl_0_218 br_0_218 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c218
+ bl_0_218 br_0_218 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c218
+ bl_0_218 br_0_218 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c218
+ bl_0_218 br_0_218 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c218
+ bl_0_218 br_0_218 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c218
+ bl_0_218 br_0_218 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c218
+ bl_0_218 br_0_218 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c218
+ bl_0_218 br_0_218 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c218
+ bl_0_218 br_0_218 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c218
+ bl_0_218 br_0_218 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c218
+ bl_0_218 br_0_218 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c218
+ bl_0_218 br_0_218 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c218
+ bl_0_218 br_0_218 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c218
+ bl_0_218 br_0_218 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c218
+ bl_0_218 br_0_218 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c218
+ bl_0_218 br_0_218 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c218
+ bl_0_218 br_0_218 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c218
+ bl_0_218 br_0_218 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c218
+ bl_0_218 br_0_218 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c218
+ bl_0_218 br_0_218 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c218
+ bl_0_218 br_0_218 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c218
+ bl_0_218 br_0_218 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c218
+ bl_0_218 br_0_218 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c218
+ bl_0_218 br_0_218 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c218
+ bl_0_218 br_0_218 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c218
+ bl_0_218 br_0_218 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c218
+ bl_0_218 br_0_218 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c218
+ bl_0_218 br_0_218 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c218
+ bl_0_218 br_0_218 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c218
+ bl_0_218 br_0_218 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c218
+ bl_0_218 br_0_218 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c218
+ bl_0_218 br_0_218 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c218
+ bl_0_218 br_0_218 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c218
+ bl_0_218 br_0_218 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c218
+ bl_0_218 br_0_218 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c218
+ bl_0_218 br_0_218 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c218
+ bl_0_218 br_0_218 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c218
+ bl_0_218 br_0_218 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c218
+ bl_0_218 br_0_218 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c218
+ bl_0_218 br_0_218 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c218
+ bl_0_218 br_0_218 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c218
+ bl_0_218 br_0_218 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c218
+ bl_0_218 br_0_218 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c219
+ bl_0_219 br_0_219 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c219
+ bl_0_219 br_0_219 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c219
+ bl_0_219 br_0_219 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c219
+ bl_0_219 br_0_219 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c219
+ bl_0_219 br_0_219 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c219
+ bl_0_219 br_0_219 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c219
+ bl_0_219 br_0_219 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c219
+ bl_0_219 br_0_219 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c219
+ bl_0_219 br_0_219 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c219
+ bl_0_219 br_0_219 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c219
+ bl_0_219 br_0_219 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c219
+ bl_0_219 br_0_219 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c219
+ bl_0_219 br_0_219 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c219
+ bl_0_219 br_0_219 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c219
+ bl_0_219 br_0_219 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c219
+ bl_0_219 br_0_219 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c219
+ bl_0_219 br_0_219 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c219
+ bl_0_219 br_0_219 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c219
+ bl_0_219 br_0_219 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c219
+ bl_0_219 br_0_219 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c219
+ bl_0_219 br_0_219 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c219
+ bl_0_219 br_0_219 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c219
+ bl_0_219 br_0_219 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c219
+ bl_0_219 br_0_219 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c219
+ bl_0_219 br_0_219 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c219
+ bl_0_219 br_0_219 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c219
+ bl_0_219 br_0_219 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c219
+ bl_0_219 br_0_219 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c219
+ bl_0_219 br_0_219 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c219
+ bl_0_219 br_0_219 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c219
+ bl_0_219 br_0_219 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c219
+ bl_0_219 br_0_219 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c219
+ bl_0_219 br_0_219 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c219
+ bl_0_219 br_0_219 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c219
+ bl_0_219 br_0_219 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c219
+ bl_0_219 br_0_219 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c219
+ bl_0_219 br_0_219 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c219
+ bl_0_219 br_0_219 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c219
+ bl_0_219 br_0_219 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c219
+ bl_0_219 br_0_219 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c219
+ bl_0_219 br_0_219 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c219
+ bl_0_219 br_0_219 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c219
+ bl_0_219 br_0_219 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c219
+ bl_0_219 br_0_219 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c220
+ bl_0_220 br_0_220 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c220
+ bl_0_220 br_0_220 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c220
+ bl_0_220 br_0_220 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c220
+ bl_0_220 br_0_220 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c220
+ bl_0_220 br_0_220 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c220
+ bl_0_220 br_0_220 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c220
+ bl_0_220 br_0_220 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c220
+ bl_0_220 br_0_220 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c220
+ bl_0_220 br_0_220 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c220
+ bl_0_220 br_0_220 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c220
+ bl_0_220 br_0_220 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c220
+ bl_0_220 br_0_220 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c220
+ bl_0_220 br_0_220 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c220
+ bl_0_220 br_0_220 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c220
+ bl_0_220 br_0_220 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c220
+ bl_0_220 br_0_220 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c220
+ bl_0_220 br_0_220 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c220
+ bl_0_220 br_0_220 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c220
+ bl_0_220 br_0_220 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c220
+ bl_0_220 br_0_220 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c220
+ bl_0_220 br_0_220 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c220
+ bl_0_220 br_0_220 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c220
+ bl_0_220 br_0_220 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c220
+ bl_0_220 br_0_220 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c220
+ bl_0_220 br_0_220 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c220
+ bl_0_220 br_0_220 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c220
+ bl_0_220 br_0_220 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c220
+ bl_0_220 br_0_220 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c220
+ bl_0_220 br_0_220 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c220
+ bl_0_220 br_0_220 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c220
+ bl_0_220 br_0_220 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c220
+ bl_0_220 br_0_220 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c220
+ bl_0_220 br_0_220 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c220
+ bl_0_220 br_0_220 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c220
+ bl_0_220 br_0_220 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c220
+ bl_0_220 br_0_220 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c220
+ bl_0_220 br_0_220 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c220
+ bl_0_220 br_0_220 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c220
+ bl_0_220 br_0_220 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c220
+ bl_0_220 br_0_220 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c220
+ bl_0_220 br_0_220 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c220
+ bl_0_220 br_0_220 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c220
+ bl_0_220 br_0_220 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c220
+ bl_0_220 br_0_220 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c221
+ bl_0_221 br_0_221 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c221
+ bl_0_221 br_0_221 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c221
+ bl_0_221 br_0_221 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c221
+ bl_0_221 br_0_221 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c221
+ bl_0_221 br_0_221 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c221
+ bl_0_221 br_0_221 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c221
+ bl_0_221 br_0_221 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c221
+ bl_0_221 br_0_221 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c221
+ bl_0_221 br_0_221 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c221
+ bl_0_221 br_0_221 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c221
+ bl_0_221 br_0_221 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c221
+ bl_0_221 br_0_221 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c221
+ bl_0_221 br_0_221 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c221
+ bl_0_221 br_0_221 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c221
+ bl_0_221 br_0_221 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c221
+ bl_0_221 br_0_221 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c221
+ bl_0_221 br_0_221 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c221
+ bl_0_221 br_0_221 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c221
+ bl_0_221 br_0_221 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c221
+ bl_0_221 br_0_221 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c221
+ bl_0_221 br_0_221 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c221
+ bl_0_221 br_0_221 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c221
+ bl_0_221 br_0_221 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c221
+ bl_0_221 br_0_221 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c221
+ bl_0_221 br_0_221 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c221
+ bl_0_221 br_0_221 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c221
+ bl_0_221 br_0_221 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c221
+ bl_0_221 br_0_221 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c221
+ bl_0_221 br_0_221 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c221
+ bl_0_221 br_0_221 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c221
+ bl_0_221 br_0_221 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c221
+ bl_0_221 br_0_221 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c221
+ bl_0_221 br_0_221 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c221
+ bl_0_221 br_0_221 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c221
+ bl_0_221 br_0_221 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c221
+ bl_0_221 br_0_221 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c221
+ bl_0_221 br_0_221 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c221
+ bl_0_221 br_0_221 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c221
+ bl_0_221 br_0_221 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c221
+ bl_0_221 br_0_221 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c221
+ bl_0_221 br_0_221 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c221
+ bl_0_221 br_0_221 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c221
+ bl_0_221 br_0_221 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c221
+ bl_0_221 br_0_221 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c222
+ bl_0_222 br_0_222 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c222
+ bl_0_222 br_0_222 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c222
+ bl_0_222 br_0_222 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c222
+ bl_0_222 br_0_222 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c222
+ bl_0_222 br_0_222 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c222
+ bl_0_222 br_0_222 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c222
+ bl_0_222 br_0_222 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c222
+ bl_0_222 br_0_222 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c222
+ bl_0_222 br_0_222 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c222
+ bl_0_222 br_0_222 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c222
+ bl_0_222 br_0_222 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c222
+ bl_0_222 br_0_222 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c222
+ bl_0_222 br_0_222 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c222
+ bl_0_222 br_0_222 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c222
+ bl_0_222 br_0_222 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c222
+ bl_0_222 br_0_222 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c222
+ bl_0_222 br_0_222 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c222
+ bl_0_222 br_0_222 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c222
+ bl_0_222 br_0_222 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c222
+ bl_0_222 br_0_222 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c222
+ bl_0_222 br_0_222 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c222
+ bl_0_222 br_0_222 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c222
+ bl_0_222 br_0_222 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c222
+ bl_0_222 br_0_222 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c222
+ bl_0_222 br_0_222 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c222
+ bl_0_222 br_0_222 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c222
+ bl_0_222 br_0_222 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c222
+ bl_0_222 br_0_222 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c222
+ bl_0_222 br_0_222 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c222
+ bl_0_222 br_0_222 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c222
+ bl_0_222 br_0_222 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c222
+ bl_0_222 br_0_222 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c222
+ bl_0_222 br_0_222 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c222
+ bl_0_222 br_0_222 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c222
+ bl_0_222 br_0_222 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c222
+ bl_0_222 br_0_222 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c222
+ bl_0_222 br_0_222 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c222
+ bl_0_222 br_0_222 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c222
+ bl_0_222 br_0_222 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c222
+ bl_0_222 br_0_222 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c222
+ bl_0_222 br_0_222 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c222
+ bl_0_222 br_0_222 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c222
+ bl_0_222 br_0_222 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c222
+ bl_0_222 br_0_222 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c223
+ bl_0_223 br_0_223 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c223
+ bl_0_223 br_0_223 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c223
+ bl_0_223 br_0_223 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c223
+ bl_0_223 br_0_223 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c223
+ bl_0_223 br_0_223 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c223
+ bl_0_223 br_0_223 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c223
+ bl_0_223 br_0_223 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c223
+ bl_0_223 br_0_223 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c223
+ bl_0_223 br_0_223 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c223
+ bl_0_223 br_0_223 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c223
+ bl_0_223 br_0_223 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c223
+ bl_0_223 br_0_223 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c223
+ bl_0_223 br_0_223 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c223
+ bl_0_223 br_0_223 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c223
+ bl_0_223 br_0_223 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c223
+ bl_0_223 br_0_223 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c223
+ bl_0_223 br_0_223 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c223
+ bl_0_223 br_0_223 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c223
+ bl_0_223 br_0_223 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c223
+ bl_0_223 br_0_223 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c223
+ bl_0_223 br_0_223 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c223
+ bl_0_223 br_0_223 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c223
+ bl_0_223 br_0_223 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c223
+ bl_0_223 br_0_223 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c223
+ bl_0_223 br_0_223 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c223
+ bl_0_223 br_0_223 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c223
+ bl_0_223 br_0_223 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c223
+ bl_0_223 br_0_223 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c223
+ bl_0_223 br_0_223 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c223
+ bl_0_223 br_0_223 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c223
+ bl_0_223 br_0_223 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c223
+ bl_0_223 br_0_223 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c223
+ bl_0_223 br_0_223 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c223
+ bl_0_223 br_0_223 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c223
+ bl_0_223 br_0_223 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c223
+ bl_0_223 br_0_223 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c223
+ bl_0_223 br_0_223 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c223
+ bl_0_223 br_0_223 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c223
+ bl_0_223 br_0_223 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c223
+ bl_0_223 br_0_223 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c223
+ bl_0_223 br_0_223 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c223
+ bl_0_223 br_0_223 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c223
+ bl_0_223 br_0_223 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c223
+ bl_0_223 br_0_223 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c224
+ bl_0_224 br_0_224 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c224
+ bl_0_224 br_0_224 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c224
+ bl_0_224 br_0_224 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c224
+ bl_0_224 br_0_224 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c224
+ bl_0_224 br_0_224 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c224
+ bl_0_224 br_0_224 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c224
+ bl_0_224 br_0_224 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c224
+ bl_0_224 br_0_224 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c224
+ bl_0_224 br_0_224 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c224
+ bl_0_224 br_0_224 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c224
+ bl_0_224 br_0_224 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c224
+ bl_0_224 br_0_224 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c224
+ bl_0_224 br_0_224 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c224
+ bl_0_224 br_0_224 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c224
+ bl_0_224 br_0_224 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c224
+ bl_0_224 br_0_224 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c224
+ bl_0_224 br_0_224 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c224
+ bl_0_224 br_0_224 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c224
+ bl_0_224 br_0_224 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c224
+ bl_0_224 br_0_224 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c224
+ bl_0_224 br_0_224 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c224
+ bl_0_224 br_0_224 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c224
+ bl_0_224 br_0_224 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c224
+ bl_0_224 br_0_224 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c224
+ bl_0_224 br_0_224 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c224
+ bl_0_224 br_0_224 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c224
+ bl_0_224 br_0_224 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c224
+ bl_0_224 br_0_224 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c224
+ bl_0_224 br_0_224 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c224
+ bl_0_224 br_0_224 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c224
+ bl_0_224 br_0_224 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c224
+ bl_0_224 br_0_224 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c224
+ bl_0_224 br_0_224 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c224
+ bl_0_224 br_0_224 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c224
+ bl_0_224 br_0_224 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c224
+ bl_0_224 br_0_224 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c224
+ bl_0_224 br_0_224 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c224
+ bl_0_224 br_0_224 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c224
+ bl_0_224 br_0_224 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c224
+ bl_0_224 br_0_224 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c224
+ bl_0_224 br_0_224 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c224
+ bl_0_224 br_0_224 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c224
+ bl_0_224 br_0_224 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c224
+ bl_0_224 br_0_224 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c225
+ bl_0_225 br_0_225 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c225
+ bl_0_225 br_0_225 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c225
+ bl_0_225 br_0_225 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c225
+ bl_0_225 br_0_225 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c225
+ bl_0_225 br_0_225 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c225
+ bl_0_225 br_0_225 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c225
+ bl_0_225 br_0_225 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c225
+ bl_0_225 br_0_225 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c225
+ bl_0_225 br_0_225 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c225
+ bl_0_225 br_0_225 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c225
+ bl_0_225 br_0_225 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c225
+ bl_0_225 br_0_225 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c225
+ bl_0_225 br_0_225 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c225
+ bl_0_225 br_0_225 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c225
+ bl_0_225 br_0_225 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c225
+ bl_0_225 br_0_225 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c225
+ bl_0_225 br_0_225 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c225
+ bl_0_225 br_0_225 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c225
+ bl_0_225 br_0_225 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c225
+ bl_0_225 br_0_225 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c225
+ bl_0_225 br_0_225 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c225
+ bl_0_225 br_0_225 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c225
+ bl_0_225 br_0_225 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c225
+ bl_0_225 br_0_225 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c225
+ bl_0_225 br_0_225 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c225
+ bl_0_225 br_0_225 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c225
+ bl_0_225 br_0_225 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c225
+ bl_0_225 br_0_225 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c225
+ bl_0_225 br_0_225 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c225
+ bl_0_225 br_0_225 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c225
+ bl_0_225 br_0_225 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c225
+ bl_0_225 br_0_225 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c225
+ bl_0_225 br_0_225 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c225
+ bl_0_225 br_0_225 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c225
+ bl_0_225 br_0_225 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c225
+ bl_0_225 br_0_225 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c225
+ bl_0_225 br_0_225 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c225
+ bl_0_225 br_0_225 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c225
+ bl_0_225 br_0_225 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c225
+ bl_0_225 br_0_225 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c225
+ bl_0_225 br_0_225 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c225
+ bl_0_225 br_0_225 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c225
+ bl_0_225 br_0_225 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c225
+ bl_0_225 br_0_225 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c226
+ bl_0_226 br_0_226 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c226
+ bl_0_226 br_0_226 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c226
+ bl_0_226 br_0_226 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c226
+ bl_0_226 br_0_226 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c226
+ bl_0_226 br_0_226 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c226
+ bl_0_226 br_0_226 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c226
+ bl_0_226 br_0_226 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c226
+ bl_0_226 br_0_226 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c226
+ bl_0_226 br_0_226 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c226
+ bl_0_226 br_0_226 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c226
+ bl_0_226 br_0_226 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c226
+ bl_0_226 br_0_226 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c226
+ bl_0_226 br_0_226 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c226
+ bl_0_226 br_0_226 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c226
+ bl_0_226 br_0_226 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c226
+ bl_0_226 br_0_226 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c226
+ bl_0_226 br_0_226 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c226
+ bl_0_226 br_0_226 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c226
+ bl_0_226 br_0_226 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c226
+ bl_0_226 br_0_226 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c226
+ bl_0_226 br_0_226 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c226
+ bl_0_226 br_0_226 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c226
+ bl_0_226 br_0_226 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c226
+ bl_0_226 br_0_226 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c226
+ bl_0_226 br_0_226 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c226
+ bl_0_226 br_0_226 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c226
+ bl_0_226 br_0_226 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c226
+ bl_0_226 br_0_226 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c226
+ bl_0_226 br_0_226 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c226
+ bl_0_226 br_0_226 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c226
+ bl_0_226 br_0_226 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c226
+ bl_0_226 br_0_226 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c226
+ bl_0_226 br_0_226 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c226
+ bl_0_226 br_0_226 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c226
+ bl_0_226 br_0_226 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c226
+ bl_0_226 br_0_226 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c226
+ bl_0_226 br_0_226 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c226
+ bl_0_226 br_0_226 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c226
+ bl_0_226 br_0_226 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c226
+ bl_0_226 br_0_226 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c226
+ bl_0_226 br_0_226 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c226
+ bl_0_226 br_0_226 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c226
+ bl_0_226 br_0_226 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c226
+ bl_0_226 br_0_226 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c227
+ bl_0_227 br_0_227 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c227
+ bl_0_227 br_0_227 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c227
+ bl_0_227 br_0_227 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c227
+ bl_0_227 br_0_227 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c227
+ bl_0_227 br_0_227 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c227
+ bl_0_227 br_0_227 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c227
+ bl_0_227 br_0_227 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c227
+ bl_0_227 br_0_227 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c227
+ bl_0_227 br_0_227 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c227
+ bl_0_227 br_0_227 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c227
+ bl_0_227 br_0_227 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c227
+ bl_0_227 br_0_227 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c227
+ bl_0_227 br_0_227 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c227
+ bl_0_227 br_0_227 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c227
+ bl_0_227 br_0_227 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c227
+ bl_0_227 br_0_227 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c227
+ bl_0_227 br_0_227 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c227
+ bl_0_227 br_0_227 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c227
+ bl_0_227 br_0_227 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c227
+ bl_0_227 br_0_227 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c227
+ bl_0_227 br_0_227 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c227
+ bl_0_227 br_0_227 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c227
+ bl_0_227 br_0_227 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c227
+ bl_0_227 br_0_227 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c227
+ bl_0_227 br_0_227 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c227
+ bl_0_227 br_0_227 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c227
+ bl_0_227 br_0_227 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c227
+ bl_0_227 br_0_227 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c227
+ bl_0_227 br_0_227 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c227
+ bl_0_227 br_0_227 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c227
+ bl_0_227 br_0_227 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c227
+ bl_0_227 br_0_227 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c227
+ bl_0_227 br_0_227 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c227
+ bl_0_227 br_0_227 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c227
+ bl_0_227 br_0_227 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c227
+ bl_0_227 br_0_227 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c227
+ bl_0_227 br_0_227 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c227
+ bl_0_227 br_0_227 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c227
+ bl_0_227 br_0_227 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c227
+ bl_0_227 br_0_227 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c227
+ bl_0_227 br_0_227 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c227
+ bl_0_227 br_0_227 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c227
+ bl_0_227 br_0_227 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c227
+ bl_0_227 br_0_227 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c228
+ bl_0_228 br_0_228 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c228
+ bl_0_228 br_0_228 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c228
+ bl_0_228 br_0_228 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c228
+ bl_0_228 br_0_228 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c228
+ bl_0_228 br_0_228 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c228
+ bl_0_228 br_0_228 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c228
+ bl_0_228 br_0_228 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c228
+ bl_0_228 br_0_228 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c228
+ bl_0_228 br_0_228 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c228
+ bl_0_228 br_0_228 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c228
+ bl_0_228 br_0_228 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c228
+ bl_0_228 br_0_228 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c228
+ bl_0_228 br_0_228 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c228
+ bl_0_228 br_0_228 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c228
+ bl_0_228 br_0_228 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c228
+ bl_0_228 br_0_228 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c228
+ bl_0_228 br_0_228 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c228
+ bl_0_228 br_0_228 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c228
+ bl_0_228 br_0_228 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c228
+ bl_0_228 br_0_228 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c228
+ bl_0_228 br_0_228 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c228
+ bl_0_228 br_0_228 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c228
+ bl_0_228 br_0_228 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c228
+ bl_0_228 br_0_228 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c228
+ bl_0_228 br_0_228 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c228
+ bl_0_228 br_0_228 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c228
+ bl_0_228 br_0_228 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c228
+ bl_0_228 br_0_228 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c228
+ bl_0_228 br_0_228 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c228
+ bl_0_228 br_0_228 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c228
+ bl_0_228 br_0_228 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c228
+ bl_0_228 br_0_228 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c228
+ bl_0_228 br_0_228 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c228
+ bl_0_228 br_0_228 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c228
+ bl_0_228 br_0_228 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c228
+ bl_0_228 br_0_228 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c228
+ bl_0_228 br_0_228 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c228
+ bl_0_228 br_0_228 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c228
+ bl_0_228 br_0_228 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c228
+ bl_0_228 br_0_228 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c228
+ bl_0_228 br_0_228 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c228
+ bl_0_228 br_0_228 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c228
+ bl_0_228 br_0_228 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c228
+ bl_0_228 br_0_228 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c229
+ bl_0_229 br_0_229 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c229
+ bl_0_229 br_0_229 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c229
+ bl_0_229 br_0_229 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c229
+ bl_0_229 br_0_229 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c229
+ bl_0_229 br_0_229 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c229
+ bl_0_229 br_0_229 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c229
+ bl_0_229 br_0_229 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c229
+ bl_0_229 br_0_229 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c229
+ bl_0_229 br_0_229 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c229
+ bl_0_229 br_0_229 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c229
+ bl_0_229 br_0_229 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c229
+ bl_0_229 br_0_229 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c229
+ bl_0_229 br_0_229 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c229
+ bl_0_229 br_0_229 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c229
+ bl_0_229 br_0_229 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c229
+ bl_0_229 br_0_229 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c229
+ bl_0_229 br_0_229 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c229
+ bl_0_229 br_0_229 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c229
+ bl_0_229 br_0_229 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c229
+ bl_0_229 br_0_229 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c229
+ bl_0_229 br_0_229 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c229
+ bl_0_229 br_0_229 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c229
+ bl_0_229 br_0_229 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c229
+ bl_0_229 br_0_229 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c229
+ bl_0_229 br_0_229 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c229
+ bl_0_229 br_0_229 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c229
+ bl_0_229 br_0_229 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c229
+ bl_0_229 br_0_229 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c229
+ bl_0_229 br_0_229 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c229
+ bl_0_229 br_0_229 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c229
+ bl_0_229 br_0_229 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c229
+ bl_0_229 br_0_229 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c229
+ bl_0_229 br_0_229 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c229
+ bl_0_229 br_0_229 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c229
+ bl_0_229 br_0_229 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c229
+ bl_0_229 br_0_229 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c229
+ bl_0_229 br_0_229 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c229
+ bl_0_229 br_0_229 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c229
+ bl_0_229 br_0_229 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c229
+ bl_0_229 br_0_229 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c229
+ bl_0_229 br_0_229 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c229
+ bl_0_229 br_0_229 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c229
+ bl_0_229 br_0_229 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c229
+ bl_0_229 br_0_229 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c230
+ bl_0_230 br_0_230 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c230
+ bl_0_230 br_0_230 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c230
+ bl_0_230 br_0_230 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c230
+ bl_0_230 br_0_230 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c230
+ bl_0_230 br_0_230 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c230
+ bl_0_230 br_0_230 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c230
+ bl_0_230 br_0_230 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c230
+ bl_0_230 br_0_230 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c230
+ bl_0_230 br_0_230 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c230
+ bl_0_230 br_0_230 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c230
+ bl_0_230 br_0_230 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c230
+ bl_0_230 br_0_230 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c230
+ bl_0_230 br_0_230 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c230
+ bl_0_230 br_0_230 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c230
+ bl_0_230 br_0_230 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c230
+ bl_0_230 br_0_230 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c230
+ bl_0_230 br_0_230 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c230
+ bl_0_230 br_0_230 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c230
+ bl_0_230 br_0_230 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c230
+ bl_0_230 br_0_230 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c230
+ bl_0_230 br_0_230 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c230
+ bl_0_230 br_0_230 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c230
+ bl_0_230 br_0_230 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c230
+ bl_0_230 br_0_230 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c230
+ bl_0_230 br_0_230 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c230
+ bl_0_230 br_0_230 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c230
+ bl_0_230 br_0_230 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c230
+ bl_0_230 br_0_230 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c230
+ bl_0_230 br_0_230 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c230
+ bl_0_230 br_0_230 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c230
+ bl_0_230 br_0_230 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c230
+ bl_0_230 br_0_230 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c230
+ bl_0_230 br_0_230 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c230
+ bl_0_230 br_0_230 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c230
+ bl_0_230 br_0_230 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c230
+ bl_0_230 br_0_230 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c230
+ bl_0_230 br_0_230 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c230
+ bl_0_230 br_0_230 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c230
+ bl_0_230 br_0_230 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c230
+ bl_0_230 br_0_230 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c230
+ bl_0_230 br_0_230 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c230
+ bl_0_230 br_0_230 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c230
+ bl_0_230 br_0_230 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c230
+ bl_0_230 br_0_230 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c231
+ bl_0_231 br_0_231 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c231
+ bl_0_231 br_0_231 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c231
+ bl_0_231 br_0_231 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c231
+ bl_0_231 br_0_231 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c231
+ bl_0_231 br_0_231 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c231
+ bl_0_231 br_0_231 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c231
+ bl_0_231 br_0_231 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c231
+ bl_0_231 br_0_231 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c231
+ bl_0_231 br_0_231 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c231
+ bl_0_231 br_0_231 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c231
+ bl_0_231 br_0_231 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c231
+ bl_0_231 br_0_231 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c231
+ bl_0_231 br_0_231 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c231
+ bl_0_231 br_0_231 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c231
+ bl_0_231 br_0_231 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c231
+ bl_0_231 br_0_231 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c231
+ bl_0_231 br_0_231 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c231
+ bl_0_231 br_0_231 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c231
+ bl_0_231 br_0_231 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c231
+ bl_0_231 br_0_231 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c231
+ bl_0_231 br_0_231 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c231
+ bl_0_231 br_0_231 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c231
+ bl_0_231 br_0_231 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c231
+ bl_0_231 br_0_231 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c231
+ bl_0_231 br_0_231 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c231
+ bl_0_231 br_0_231 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c231
+ bl_0_231 br_0_231 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c231
+ bl_0_231 br_0_231 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c231
+ bl_0_231 br_0_231 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c231
+ bl_0_231 br_0_231 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c231
+ bl_0_231 br_0_231 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c231
+ bl_0_231 br_0_231 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c231
+ bl_0_231 br_0_231 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c231
+ bl_0_231 br_0_231 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c231
+ bl_0_231 br_0_231 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c231
+ bl_0_231 br_0_231 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c231
+ bl_0_231 br_0_231 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c231
+ bl_0_231 br_0_231 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c231
+ bl_0_231 br_0_231 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c231
+ bl_0_231 br_0_231 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c231
+ bl_0_231 br_0_231 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c231
+ bl_0_231 br_0_231 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c231
+ bl_0_231 br_0_231 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c231
+ bl_0_231 br_0_231 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c232
+ bl_0_232 br_0_232 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c232
+ bl_0_232 br_0_232 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c232
+ bl_0_232 br_0_232 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c232
+ bl_0_232 br_0_232 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c232
+ bl_0_232 br_0_232 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c232
+ bl_0_232 br_0_232 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c232
+ bl_0_232 br_0_232 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c232
+ bl_0_232 br_0_232 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c232
+ bl_0_232 br_0_232 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c232
+ bl_0_232 br_0_232 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c232
+ bl_0_232 br_0_232 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c232
+ bl_0_232 br_0_232 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c232
+ bl_0_232 br_0_232 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c232
+ bl_0_232 br_0_232 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c232
+ bl_0_232 br_0_232 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c232
+ bl_0_232 br_0_232 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c232
+ bl_0_232 br_0_232 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c232
+ bl_0_232 br_0_232 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c232
+ bl_0_232 br_0_232 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c232
+ bl_0_232 br_0_232 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c232
+ bl_0_232 br_0_232 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c232
+ bl_0_232 br_0_232 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c232
+ bl_0_232 br_0_232 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c232
+ bl_0_232 br_0_232 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c232
+ bl_0_232 br_0_232 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c232
+ bl_0_232 br_0_232 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c232
+ bl_0_232 br_0_232 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c232
+ bl_0_232 br_0_232 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c232
+ bl_0_232 br_0_232 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c232
+ bl_0_232 br_0_232 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c232
+ bl_0_232 br_0_232 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c232
+ bl_0_232 br_0_232 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c232
+ bl_0_232 br_0_232 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c232
+ bl_0_232 br_0_232 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c232
+ bl_0_232 br_0_232 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c232
+ bl_0_232 br_0_232 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c232
+ bl_0_232 br_0_232 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c232
+ bl_0_232 br_0_232 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c232
+ bl_0_232 br_0_232 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c232
+ bl_0_232 br_0_232 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c232
+ bl_0_232 br_0_232 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c232
+ bl_0_232 br_0_232 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c232
+ bl_0_232 br_0_232 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c232
+ bl_0_232 br_0_232 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c233
+ bl_0_233 br_0_233 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c233
+ bl_0_233 br_0_233 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c233
+ bl_0_233 br_0_233 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c233
+ bl_0_233 br_0_233 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c233
+ bl_0_233 br_0_233 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c233
+ bl_0_233 br_0_233 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c233
+ bl_0_233 br_0_233 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c233
+ bl_0_233 br_0_233 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c233
+ bl_0_233 br_0_233 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c233
+ bl_0_233 br_0_233 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c233
+ bl_0_233 br_0_233 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c233
+ bl_0_233 br_0_233 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c233
+ bl_0_233 br_0_233 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c233
+ bl_0_233 br_0_233 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c233
+ bl_0_233 br_0_233 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c233
+ bl_0_233 br_0_233 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c233
+ bl_0_233 br_0_233 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c233
+ bl_0_233 br_0_233 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c233
+ bl_0_233 br_0_233 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c233
+ bl_0_233 br_0_233 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c233
+ bl_0_233 br_0_233 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c233
+ bl_0_233 br_0_233 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c233
+ bl_0_233 br_0_233 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c233
+ bl_0_233 br_0_233 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c233
+ bl_0_233 br_0_233 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c233
+ bl_0_233 br_0_233 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c233
+ bl_0_233 br_0_233 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c233
+ bl_0_233 br_0_233 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c233
+ bl_0_233 br_0_233 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c233
+ bl_0_233 br_0_233 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c233
+ bl_0_233 br_0_233 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c233
+ bl_0_233 br_0_233 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c233
+ bl_0_233 br_0_233 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c233
+ bl_0_233 br_0_233 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c233
+ bl_0_233 br_0_233 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c233
+ bl_0_233 br_0_233 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c233
+ bl_0_233 br_0_233 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c233
+ bl_0_233 br_0_233 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c233
+ bl_0_233 br_0_233 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c233
+ bl_0_233 br_0_233 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c233
+ bl_0_233 br_0_233 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c233
+ bl_0_233 br_0_233 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c233
+ bl_0_233 br_0_233 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c233
+ bl_0_233 br_0_233 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c234
+ bl_0_234 br_0_234 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c234
+ bl_0_234 br_0_234 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c234
+ bl_0_234 br_0_234 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c234
+ bl_0_234 br_0_234 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c234
+ bl_0_234 br_0_234 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c234
+ bl_0_234 br_0_234 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c234
+ bl_0_234 br_0_234 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c234
+ bl_0_234 br_0_234 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c234
+ bl_0_234 br_0_234 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c234
+ bl_0_234 br_0_234 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c234
+ bl_0_234 br_0_234 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c234
+ bl_0_234 br_0_234 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c234
+ bl_0_234 br_0_234 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c234
+ bl_0_234 br_0_234 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c234
+ bl_0_234 br_0_234 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c234
+ bl_0_234 br_0_234 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c234
+ bl_0_234 br_0_234 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c234
+ bl_0_234 br_0_234 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c234
+ bl_0_234 br_0_234 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c234
+ bl_0_234 br_0_234 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c234
+ bl_0_234 br_0_234 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c234
+ bl_0_234 br_0_234 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c234
+ bl_0_234 br_0_234 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c234
+ bl_0_234 br_0_234 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c234
+ bl_0_234 br_0_234 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c234
+ bl_0_234 br_0_234 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c234
+ bl_0_234 br_0_234 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c234
+ bl_0_234 br_0_234 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c234
+ bl_0_234 br_0_234 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c234
+ bl_0_234 br_0_234 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c234
+ bl_0_234 br_0_234 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c234
+ bl_0_234 br_0_234 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c234
+ bl_0_234 br_0_234 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c234
+ bl_0_234 br_0_234 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c234
+ bl_0_234 br_0_234 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c234
+ bl_0_234 br_0_234 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c234
+ bl_0_234 br_0_234 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c234
+ bl_0_234 br_0_234 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c234
+ bl_0_234 br_0_234 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c234
+ bl_0_234 br_0_234 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c234
+ bl_0_234 br_0_234 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c234
+ bl_0_234 br_0_234 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c234
+ bl_0_234 br_0_234 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c234
+ bl_0_234 br_0_234 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c235
+ bl_0_235 br_0_235 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c235
+ bl_0_235 br_0_235 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c235
+ bl_0_235 br_0_235 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c235
+ bl_0_235 br_0_235 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c235
+ bl_0_235 br_0_235 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c235
+ bl_0_235 br_0_235 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c235
+ bl_0_235 br_0_235 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c235
+ bl_0_235 br_0_235 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c235
+ bl_0_235 br_0_235 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c235
+ bl_0_235 br_0_235 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c235
+ bl_0_235 br_0_235 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c235
+ bl_0_235 br_0_235 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c235
+ bl_0_235 br_0_235 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c235
+ bl_0_235 br_0_235 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c235
+ bl_0_235 br_0_235 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c235
+ bl_0_235 br_0_235 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c235
+ bl_0_235 br_0_235 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c235
+ bl_0_235 br_0_235 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c235
+ bl_0_235 br_0_235 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c235
+ bl_0_235 br_0_235 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c235
+ bl_0_235 br_0_235 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c235
+ bl_0_235 br_0_235 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c235
+ bl_0_235 br_0_235 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c235
+ bl_0_235 br_0_235 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c235
+ bl_0_235 br_0_235 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c235
+ bl_0_235 br_0_235 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c235
+ bl_0_235 br_0_235 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c235
+ bl_0_235 br_0_235 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c235
+ bl_0_235 br_0_235 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c235
+ bl_0_235 br_0_235 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c235
+ bl_0_235 br_0_235 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c235
+ bl_0_235 br_0_235 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c235
+ bl_0_235 br_0_235 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c235
+ bl_0_235 br_0_235 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c235
+ bl_0_235 br_0_235 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c235
+ bl_0_235 br_0_235 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c235
+ bl_0_235 br_0_235 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c235
+ bl_0_235 br_0_235 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c235
+ bl_0_235 br_0_235 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c235
+ bl_0_235 br_0_235 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c235
+ bl_0_235 br_0_235 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c235
+ bl_0_235 br_0_235 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c235
+ bl_0_235 br_0_235 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c235
+ bl_0_235 br_0_235 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c236
+ bl_0_236 br_0_236 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c236
+ bl_0_236 br_0_236 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c236
+ bl_0_236 br_0_236 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c236
+ bl_0_236 br_0_236 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c236
+ bl_0_236 br_0_236 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c236
+ bl_0_236 br_0_236 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c236
+ bl_0_236 br_0_236 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c236
+ bl_0_236 br_0_236 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c236
+ bl_0_236 br_0_236 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c236
+ bl_0_236 br_0_236 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c236
+ bl_0_236 br_0_236 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c236
+ bl_0_236 br_0_236 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c236
+ bl_0_236 br_0_236 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c236
+ bl_0_236 br_0_236 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c236
+ bl_0_236 br_0_236 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c236
+ bl_0_236 br_0_236 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c236
+ bl_0_236 br_0_236 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c236
+ bl_0_236 br_0_236 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c236
+ bl_0_236 br_0_236 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c236
+ bl_0_236 br_0_236 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c236
+ bl_0_236 br_0_236 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c236
+ bl_0_236 br_0_236 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c236
+ bl_0_236 br_0_236 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c236
+ bl_0_236 br_0_236 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c236
+ bl_0_236 br_0_236 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c236
+ bl_0_236 br_0_236 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c236
+ bl_0_236 br_0_236 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c236
+ bl_0_236 br_0_236 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c236
+ bl_0_236 br_0_236 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c236
+ bl_0_236 br_0_236 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c236
+ bl_0_236 br_0_236 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c236
+ bl_0_236 br_0_236 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c236
+ bl_0_236 br_0_236 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c236
+ bl_0_236 br_0_236 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c236
+ bl_0_236 br_0_236 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c236
+ bl_0_236 br_0_236 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c236
+ bl_0_236 br_0_236 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c236
+ bl_0_236 br_0_236 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c236
+ bl_0_236 br_0_236 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c236
+ bl_0_236 br_0_236 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c236
+ bl_0_236 br_0_236 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c236
+ bl_0_236 br_0_236 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c236
+ bl_0_236 br_0_236 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c236
+ bl_0_236 br_0_236 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c237
+ bl_0_237 br_0_237 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c237
+ bl_0_237 br_0_237 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c237
+ bl_0_237 br_0_237 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c237
+ bl_0_237 br_0_237 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c237
+ bl_0_237 br_0_237 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c237
+ bl_0_237 br_0_237 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c237
+ bl_0_237 br_0_237 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c237
+ bl_0_237 br_0_237 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c237
+ bl_0_237 br_0_237 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c237
+ bl_0_237 br_0_237 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c237
+ bl_0_237 br_0_237 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c237
+ bl_0_237 br_0_237 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c237
+ bl_0_237 br_0_237 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c237
+ bl_0_237 br_0_237 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c237
+ bl_0_237 br_0_237 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c237
+ bl_0_237 br_0_237 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c237
+ bl_0_237 br_0_237 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c237
+ bl_0_237 br_0_237 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c237
+ bl_0_237 br_0_237 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c237
+ bl_0_237 br_0_237 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c237
+ bl_0_237 br_0_237 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c237
+ bl_0_237 br_0_237 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c237
+ bl_0_237 br_0_237 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c237
+ bl_0_237 br_0_237 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c237
+ bl_0_237 br_0_237 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c237
+ bl_0_237 br_0_237 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c237
+ bl_0_237 br_0_237 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c237
+ bl_0_237 br_0_237 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c237
+ bl_0_237 br_0_237 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c237
+ bl_0_237 br_0_237 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c237
+ bl_0_237 br_0_237 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c237
+ bl_0_237 br_0_237 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c237
+ bl_0_237 br_0_237 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c237
+ bl_0_237 br_0_237 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c237
+ bl_0_237 br_0_237 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c237
+ bl_0_237 br_0_237 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c237
+ bl_0_237 br_0_237 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c237
+ bl_0_237 br_0_237 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c237
+ bl_0_237 br_0_237 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c237
+ bl_0_237 br_0_237 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c237
+ bl_0_237 br_0_237 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c237
+ bl_0_237 br_0_237 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c237
+ bl_0_237 br_0_237 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c237
+ bl_0_237 br_0_237 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c238
+ bl_0_238 br_0_238 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c238
+ bl_0_238 br_0_238 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c238
+ bl_0_238 br_0_238 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c238
+ bl_0_238 br_0_238 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c238
+ bl_0_238 br_0_238 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c238
+ bl_0_238 br_0_238 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c238
+ bl_0_238 br_0_238 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c238
+ bl_0_238 br_0_238 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c238
+ bl_0_238 br_0_238 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c238
+ bl_0_238 br_0_238 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c238
+ bl_0_238 br_0_238 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c238
+ bl_0_238 br_0_238 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c238
+ bl_0_238 br_0_238 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c238
+ bl_0_238 br_0_238 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c238
+ bl_0_238 br_0_238 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c238
+ bl_0_238 br_0_238 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c238
+ bl_0_238 br_0_238 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c238
+ bl_0_238 br_0_238 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c238
+ bl_0_238 br_0_238 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c238
+ bl_0_238 br_0_238 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c238
+ bl_0_238 br_0_238 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c238
+ bl_0_238 br_0_238 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c238
+ bl_0_238 br_0_238 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c238
+ bl_0_238 br_0_238 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c238
+ bl_0_238 br_0_238 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c238
+ bl_0_238 br_0_238 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c238
+ bl_0_238 br_0_238 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c238
+ bl_0_238 br_0_238 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c238
+ bl_0_238 br_0_238 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c238
+ bl_0_238 br_0_238 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c238
+ bl_0_238 br_0_238 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c238
+ bl_0_238 br_0_238 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c238
+ bl_0_238 br_0_238 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c238
+ bl_0_238 br_0_238 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c238
+ bl_0_238 br_0_238 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c238
+ bl_0_238 br_0_238 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c238
+ bl_0_238 br_0_238 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c238
+ bl_0_238 br_0_238 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c238
+ bl_0_238 br_0_238 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c238
+ bl_0_238 br_0_238 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c238
+ bl_0_238 br_0_238 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c238
+ bl_0_238 br_0_238 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c238
+ bl_0_238 br_0_238 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c238
+ bl_0_238 br_0_238 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c239
+ bl_0_239 br_0_239 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c239
+ bl_0_239 br_0_239 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c239
+ bl_0_239 br_0_239 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c239
+ bl_0_239 br_0_239 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c239
+ bl_0_239 br_0_239 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c239
+ bl_0_239 br_0_239 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c239
+ bl_0_239 br_0_239 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c239
+ bl_0_239 br_0_239 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c239
+ bl_0_239 br_0_239 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c239
+ bl_0_239 br_0_239 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c239
+ bl_0_239 br_0_239 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c239
+ bl_0_239 br_0_239 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c239
+ bl_0_239 br_0_239 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c239
+ bl_0_239 br_0_239 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c239
+ bl_0_239 br_0_239 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c239
+ bl_0_239 br_0_239 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c239
+ bl_0_239 br_0_239 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c239
+ bl_0_239 br_0_239 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c239
+ bl_0_239 br_0_239 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c239
+ bl_0_239 br_0_239 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c239
+ bl_0_239 br_0_239 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c239
+ bl_0_239 br_0_239 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c239
+ bl_0_239 br_0_239 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c239
+ bl_0_239 br_0_239 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c239
+ bl_0_239 br_0_239 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c239
+ bl_0_239 br_0_239 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c239
+ bl_0_239 br_0_239 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c239
+ bl_0_239 br_0_239 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c239
+ bl_0_239 br_0_239 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c239
+ bl_0_239 br_0_239 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c239
+ bl_0_239 br_0_239 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c239
+ bl_0_239 br_0_239 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c239
+ bl_0_239 br_0_239 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c239
+ bl_0_239 br_0_239 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c239
+ bl_0_239 br_0_239 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c239
+ bl_0_239 br_0_239 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c239
+ bl_0_239 br_0_239 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c239
+ bl_0_239 br_0_239 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c239
+ bl_0_239 br_0_239 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c239
+ bl_0_239 br_0_239 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c239
+ bl_0_239 br_0_239 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c239
+ bl_0_239 br_0_239 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c239
+ bl_0_239 br_0_239 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c239
+ bl_0_239 br_0_239 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c240
+ bl_0_240 br_0_240 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c240
+ bl_0_240 br_0_240 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c240
+ bl_0_240 br_0_240 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c240
+ bl_0_240 br_0_240 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c240
+ bl_0_240 br_0_240 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c240
+ bl_0_240 br_0_240 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c240
+ bl_0_240 br_0_240 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c240
+ bl_0_240 br_0_240 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c240
+ bl_0_240 br_0_240 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c240
+ bl_0_240 br_0_240 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c240
+ bl_0_240 br_0_240 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c240
+ bl_0_240 br_0_240 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c240
+ bl_0_240 br_0_240 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c240
+ bl_0_240 br_0_240 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c240
+ bl_0_240 br_0_240 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c240
+ bl_0_240 br_0_240 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c240
+ bl_0_240 br_0_240 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c240
+ bl_0_240 br_0_240 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c240
+ bl_0_240 br_0_240 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c240
+ bl_0_240 br_0_240 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c240
+ bl_0_240 br_0_240 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c240
+ bl_0_240 br_0_240 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c240
+ bl_0_240 br_0_240 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c240
+ bl_0_240 br_0_240 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c240
+ bl_0_240 br_0_240 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c240
+ bl_0_240 br_0_240 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c240
+ bl_0_240 br_0_240 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c240
+ bl_0_240 br_0_240 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c240
+ bl_0_240 br_0_240 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c240
+ bl_0_240 br_0_240 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c240
+ bl_0_240 br_0_240 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c240
+ bl_0_240 br_0_240 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c240
+ bl_0_240 br_0_240 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c240
+ bl_0_240 br_0_240 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c240
+ bl_0_240 br_0_240 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c240
+ bl_0_240 br_0_240 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c240
+ bl_0_240 br_0_240 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c240
+ bl_0_240 br_0_240 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c240
+ bl_0_240 br_0_240 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c240
+ bl_0_240 br_0_240 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c240
+ bl_0_240 br_0_240 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c240
+ bl_0_240 br_0_240 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c240
+ bl_0_240 br_0_240 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c240
+ bl_0_240 br_0_240 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c241
+ bl_0_241 br_0_241 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c241
+ bl_0_241 br_0_241 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c241
+ bl_0_241 br_0_241 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c241
+ bl_0_241 br_0_241 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c241
+ bl_0_241 br_0_241 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c241
+ bl_0_241 br_0_241 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c241
+ bl_0_241 br_0_241 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c241
+ bl_0_241 br_0_241 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c241
+ bl_0_241 br_0_241 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c241
+ bl_0_241 br_0_241 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c241
+ bl_0_241 br_0_241 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c241
+ bl_0_241 br_0_241 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c241
+ bl_0_241 br_0_241 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c241
+ bl_0_241 br_0_241 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c241
+ bl_0_241 br_0_241 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c241
+ bl_0_241 br_0_241 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c241
+ bl_0_241 br_0_241 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c241
+ bl_0_241 br_0_241 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c241
+ bl_0_241 br_0_241 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c241
+ bl_0_241 br_0_241 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c241
+ bl_0_241 br_0_241 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c241
+ bl_0_241 br_0_241 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c241
+ bl_0_241 br_0_241 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c241
+ bl_0_241 br_0_241 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c241
+ bl_0_241 br_0_241 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c241
+ bl_0_241 br_0_241 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c241
+ bl_0_241 br_0_241 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c241
+ bl_0_241 br_0_241 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c241
+ bl_0_241 br_0_241 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c241
+ bl_0_241 br_0_241 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c241
+ bl_0_241 br_0_241 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c241
+ bl_0_241 br_0_241 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c241
+ bl_0_241 br_0_241 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c241
+ bl_0_241 br_0_241 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c241
+ bl_0_241 br_0_241 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c241
+ bl_0_241 br_0_241 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c241
+ bl_0_241 br_0_241 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c241
+ bl_0_241 br_0_241 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c241
+ bl_0_241 br_0_241 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c241
+ bl_0_241 br_0_241 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c241
+ bl_0_241 br_0_241 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c241
+ bl_0_241 br_0_241 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c241
+ bl_0_241 br_0_241 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c241
+ bl_0_241 br_0_241 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c242
+ bl_0_242 br_0_242 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c242
+ bl_0_242 br_0_242 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c242
+ bl_0_242 br_0_242 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c242
+ bl_0_242 br_0_242 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c242
+ bl_0_242 br_0_242 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c242
+ bl_0_242 br_0_242 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c242
+ bl_0_242 br_0_242 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c242
+ bl_0_242 br_0_242 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c242
+ bl_0_242 br_0_242 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c242
+ bl_0_242 br_0_242 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c242
+ bl_0_242 br_0_242 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c242
+ bl_0_242 br_0_242 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c242
+ bl_0_242 br_0_242 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c242
+ bl_0_242 br_0_242 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c242
+ bl_0_242 br_0_242 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c242
+ bl_0_242 br_0_242 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c242
+ bl_0_242 br_0_242 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c242
+ bl_0_242 br_0_242 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c242
+ bl_0_242 br_0_242 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c242
+ bl_0_242 br_0_242 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c242
+ bl_0_242 br_0_242 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c242
+ bl_0_242 br_0_242 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c242
+ bl_0_242 br_0_242 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c242
+ bl_0_242 br_0_242 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c242
+ bl_0_242 br_0_242 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c242
+ bl_0_242 br_0_242 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c242
+ bl_0_242 br_0_242 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c242
+ bl_0_242 br_0_242 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c242
+ bl_0_242 br_0_242 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c242
+ bl_0_242 br_0_242 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c242
+ bl_0_242 br_0_242 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c242
+ bl_0_242 br_0_242 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c242
+ bl_0_242 br_0_242 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c242
+ bl_0_242 br_0_242 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c242
+ bl_0_242 br_0_242 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c242
+ bl_0_242 br_0_242 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c242
+ bl_0_242 br_0_242 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c242
+ bl_0_242 br_0_242 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c242
+ bl_0_242 br_0_242 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c242
+ bl_0_242 br_0_242 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c242
+ bl_0_242 br_0_242 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c242
+ bl_0_242 br_0_242 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c242
+ bl_0_242 br_0_242 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c242
+ bl_0_242 br_0_242 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c243
+ bl_0_243 br_0_243 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c243
+ bl_0_243 br_0_243 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c243
+ bl_0_243 br_0_243 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c243
+ bl_0_243 br_0_243 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c243
+ bl_0_243 br_0_243 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c243
+ bl_0_243 br_0_243 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c243
+ bl_0_243 br_0_243 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c243
+ bl_0_243 br_0_243 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c243
+ bl_0_243 br_0_243 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c243
+ bl_0_243 br_0_243 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c243
+ bl_0_243 br_0_243 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c243
+ bl_0_243 br_0_243 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c243
+ bl_0_243 br_0_243 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c243
+ bl_0_243 br_0_243 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c243
+ bl_0_243 br_0_243 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c243
+ bl_0_243 br_0_243 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c243
+ bl_0_243 br_0_243 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c243
+ bl_0_243 br_0_243 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c243
+ bl_0_243 br_0_243 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c243
+ bl_0_243 br_0_243 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c243
+ bl_0_243 br_0_243 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c243
+ bl_0_243 br_0_243 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c243
+ bl_0_243 br_0_243 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c243
+ bl_0_243 br_0_243 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c243
+ bl_0_243 br_0_243 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c243
+ bl_0_243 br_0_243 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c243
+ bl_0_243 br_0_243 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c243
+ bl_0_243 br_0_243 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c243
+ bl_0_243 br_0_243 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c243
+ bl_0_243 br_0_243 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c243
+ bl_0_243 br_0_243 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c243
+ bl_0_243 br_0_243 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c243
+ bl_0_243 br_0_243 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c243
+ bl_0_243 br_0_243 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c243
+ bl_0_243 br_0_243 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c243
+ bl_0_243 br_0_243 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c243
+ bl_0_243 br_0_243 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c243
+ bl_0_243 br_0_243 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c243
+ bl_0_243 br_0_243 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c243
+ bl_0_243 br_0_243 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c243
+ bl_0_243 br_0_243 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c243
+ bl_0_243 br_0_243 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c243
+ bl_0_243 br_0_243 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c243
+ bl_0_243 br_0_243 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c244
+ bl_0_244 br_0_244 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c244
+ bl_0_244 br_0_244 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c244
+ bl_0_244 br_0_244 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c244
+ bl_0_244 br_0_244 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c244
+ bl_0_244 br_0_244 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c244
+ bl_0_244 br_0_244 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c244
+ bl_0_244 br_0_244 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c244
+ bl_0_244 br_0_244 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c244
+ bl_0_244 br_0_244 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c244
+ bl_0_244 br_0_244 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c244
+ bl_0_244 br_0_244 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c244
+ bl_0_244 br_0_244 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c244
+ bl_0_244 br_0_244 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c244
+ bl_0_244 br_0_244 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c244
+ bl_0_244 br_0_244 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c244
+ bl_0_244 br_0_244 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c244
+ bl_0_244 br_0_244 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c244
+ bl_0_244 br_0_244 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c244
+ bl_0_244 br_0_244 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c244
+ bl_0_244 br_0_244 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c244
+ bl_0_244 br_0_244 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c244
+ bl_0_244 br_0_244 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c244
+ bl_0_244 br_0_244 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c244
+ bl_0_244 br_0_244 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c244
+ bl_0_244 br_0_244 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c244
+ bl_0_244 br_0_244 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c244
+ bl_0_244 br_0_244 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c244
+ bl_0_244 br_0_244 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c244
+ bl_0_244 br_0_244 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c244
+ bl_0_244 br_0_244 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c244
+ bl_0_244 br_0_244 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c244
+ bl_0_244 br_0_244 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c244
+ bl_0_244 br_0_244 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c244
+ bl_0_244 br_0_244 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c244
+ bl_0_244 br_0_244 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c244
+ bl_0_244 br_0_244 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c244
+ bl_0_244 br_0_244 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c244
+ bl_0_244 br_0_244 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c244
+ bl_0_244 br_0_244 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c244
+ bl_0_244 br_0_244 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c244
+ bl_0_244 br_0_244 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c244
+ bl_0_244 br_0_244 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c244
+ bl_0_244 br_0_244 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c244
+ bl_0_244 br_0_244 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c245
+ bl_0_245 br_0_245 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c245
+ bl_0_245 br_0_245 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c245
+ bl_0_245 br_0_245 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c245
+ bl_0_245 br_0_245 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c245
+ bl_0_245 br_0_245 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c245
+ bl_0_245 br_0_245 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c245
+ bl_0_245 br_0_245 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c245
+ bl_0_245 br_0_245 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c245
+ bl_0_245 br_0_245 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c245
+ bl_0_245 br_0_245 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c245
+ bl_0_245 br_0_245 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c245
+ bl_0_245 br_0_245 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c245
+ bl_0_245 br_0_245 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c245
+ bl_0_245 br_0_245 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c245
+ bl_0_245 br_0_245 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c245
+ bl_0_245 br_0_245 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c245
+ bl_0_245 br_0_245 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c245
+ bl_0_245 br_0_245 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c245
+ bl_0_245 br_0_245 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c245
+ bl_0_245 br_0_245 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c245
+ bl_0_245 br_0_245 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c245
+ bl_0_245 br_0_245 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c245
+ bl_0_245 br_0_245 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c245
+ bl_0_245 br_0_245 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c245
+ bl_0_245 br_0_245 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c245
+ bl_0_245 br_0_245 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c245
+ bl_0_245 br_0_245 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c245
+ bl_0_245 br_0_245 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c245
+ bl_0_245 br_0_245 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c245
+ bl_0_245 br_0_245 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c245
+ bl_0_245 br_0_245 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c245
+ bl_0_245 br_0_245 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c245
+ bl_0_245 br_0_245 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c245
+ bl_0_245 br_0_245 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c245
+ bl_0_245 br_0_245 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c245
+ bl_0_245 br_0_245 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c245
+ bl_0_245 br_0_245 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c245
+ bl_0_245 br_0_245 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c245
+ bl_0_245 br_0_245 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c245
+ bl_0_245 br_0_245 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c245
+ bl_0_245 br_0_245 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c245
+ bl_0_245 br_0_245 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c245
+ bl_0_245 br_0_245 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c245
+ bl_0_245 br_0_245 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c246
+ bl_0_246 br_0_246 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c246
+ bl_0_246 br_0_246 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c246
+ bl_0_246 br_0_246 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c246
+ bl_0_246 br_0_246 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c246
+ bl_0_246 br_0_246 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c246
+ bl_0_246 br_0_246 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c246
+ bl_0_246 br_0_246 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c246
+ bl_0_246 br_0_246 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c246
+ bl_0_246 br_0_246 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c246
+ bl_0_246 br_0_246 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c246
+ bl_0_246 br_0_246 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c246
+ bl_0_246 br_0_246 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c246
+ bl_0_246 br_0_246 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c246
+ bl_0_246 br_0_246 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c246
+ bl_0_246 br_0_246 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c246
+ bl_0_246 br_0_246 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c246
+ bl_0_246 br_0_246 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c246
+ bl_0_246 br_0_246 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c246
+ bl_0_246 br_0_246 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c246
+ bl_0_246 br_0_246 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c246
+ bl_0_246 br_0_246 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c246
+ bl_0_246 br_0_246 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c246
+ bl_0_246 br_0_246 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c246
+ bl_0_246 br_0_246 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c246
+ bl_0_246 br_0_246 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c246
+ bl_0_246 br_0_246 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c246
+ bl_0_246 br_0_246 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c246
+ bl_0_246 br_0_246 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c246
+ bl_0_246 br_0_246 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c246
+ bl_0_246 br_0_246 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c246
+ bl_0_246 br_0_246 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c246
+ bl_0_246 br_0_246 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c246
+ bl_0_246 br_0_246 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c246
+ bl_0_246 br_0_246 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c246
+ bl_0_246 br_0_246 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c246
+ bl_0_246 br_0_246 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c246
+ bl_0_246 br_0_246 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c246
+ bl_0_246 br_0_246 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c246
+ bl_0_246 br_0_246 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c246
+ bl_0_246 br_0_246 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c246
+ bl_0_246 br_0_246 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c246
+ bl_0_246 br_0_246 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c246
+ bl_0_246 br_0_246 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c246
+ bl_0_246 br_0_246 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c247
+ bl_0_247 br_0_247 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c247
+ bl_0_247 br_0_247 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c247
+ bl_0_247 br_0_247 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c247
+ bl_0_247 br_0_247 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c247
+ bl_0_247 br_0_247 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c247
+ bl_0_247 br_0_247 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c247
+ bl_0_247 br_0_247 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c247
+ bl_0_247 br_0_247 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c247
+ bl_0_247 br_0_247 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c247
+ bl_0_247 br_0_247 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c247
+ bl_0_247 br_0_247 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c247
+ bl_0_247 br_0_247 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c247
+ bl_0_247 br_0_247 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c247
+ bl_0_247 br_0_247 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c247
+ bl_0_247 br_0_247 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c247
+ bl_0_247 br_0_247 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c247
+ bl_0_247 br_0_247 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c247
+ bl_0_247 br_0_247 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c247
+ bl_0_247 br_0_247 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c247
+ bl_0_247 br_0_247 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c247
+ bl_0_247 br_0_247 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c247
+ bl_0_247 br_0_247 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c247
+ bl_0_247 br_0_247 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c247
+ bl_0_247 br_0_247 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c247
+ bl_0_247 br_0_247 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c247
+ bl_0_247 br_0_247 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c247
+ bl_0_247 br_0_247 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c247
+ bl_0_247 br_0_247 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c247
+ bl_0_247 br_0_247 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c247
+ bl_0_247 br_0_247 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c247
+ bl_0_247 br_0_247 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c247
+ bl_0_247 br_0_247 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c247
+ bl_0_247 br_0_247 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c247
+ bl_0_247 br_0_247 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c247
+ bl_0_247 br_0_247 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c247
+ bl_0_247 br_0_247 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c247
+ bl_0_247 br_0_247 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c247
+ bl_0_247 br_0_247 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c247
+ bl_0_247 br_0_247 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c247
+ bl_0_247 br_0_247 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c247
+ bl_0_247 br_0_247 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c247
+ bl_0_247 br_0_247 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c247
+ bl_0_247 br_0_247 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c247
+ bl_0_247 br_0_247 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c248
+ bl_0_248 br_0_248 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c248
+ bl_0_248 br_0_248 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c248
+ bl_0_248 br_0_248 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c248
+ bl_0_248 br_0_248 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c248
+ bl_0_248 br_0_248 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c248
+ bl_0_248 br_0_248 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c248
+ bl_0_248 br_0_248 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c248
+ bl_0_248 br_0_248 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c248
+ bl_0_248 br_0_248 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c248
+ bl_0_248 br_0_248 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c248
+ bl_0_248 br_0_248 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c248
+ bl_0_248 br_0_248 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c248
+ bl_0_248 br_0_248 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c248
+ bl_0_248 br_0_248 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c248
+ bl_0_248 br_0_248 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c248
+ bl_0_248 br_0_248 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c248
+ bl_0_248 br_0_248 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c248
+ bl_0_248 br_0_248 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c248
+ bl_0_248 br_0_248 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c248
+ bl_0_248 br_0_248 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c248
+ bl_0_248 br_0_248 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c248
+ bl_0_248 br_0_248 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c248
+ bl_0_248 br_0_248 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c248
+ bl_0_248 br_0_248 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c248
+ bl_0_248 br_0_248 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c248
+ bl_0_248 br_0_248 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c248
+ bl_0_248 br_0_248 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c248
+ bl_0_248 br_0_248 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c248
+ bl_0_248 br_0_248 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c248
+ bl_0_248 br_0_248 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c248
+ bl_0_248 br_0_248 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c248
+ bl_0_248 br_0_248 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c248
+ bl_0_248 br_0_248 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c248
+ bl_0_248 br_0_248 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c248
+ bl_0_248 br_0_248 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c248
+ bl_0_248 br_0_248 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c248
+ bl_0_248 br_0_248 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c248
+ bl_0_248 br_0_248 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c248
+ bl_0_248 br_0_248 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c248
+ bl_0_248 br_0_248 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c248
+ bl_0_248 br_0_248 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c248
+ bl_0_248 br_0_248 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c248
+ bl_0_248 br_0_248 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c248
+ bl_0_248 br_0_248 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c249
+ bl_0_249 br_0_249 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c249
+ bl_0_249 br_0_249 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c249
+ bl_0_249 br_0_249 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c249
+ bl_0_249 br_0_249 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c249
+ bl_0_249 br_0_249 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c249
+ bl_0_249 br_0_249 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c249
+ bl_0_249 br_0_249 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c249
+ bl_0_249 br_0_249 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c249
+ bl_0_249 br_0_249 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c249
+ bl_0_249 br_0_249 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c249
+ bl_0_249 br_0_249 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c249
+ bl_0_249 br_0_249 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c249
+ bl_0_249 br_0_249 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c249
+ bl_0_249 br_0_249 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c249
+ bl_0_249 br_0_249 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c249
+ bl_0_249 br_0_249 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c249
+ bl_0_249 br_0_249 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c249
+ bl_0_249 br_0_249 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c249
+ bl_0_249 br_0_249 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c249
+ bl_0_249 br_0_249 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c249
+ bl_0_249 br_0_249 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c249
+ bl_0_249 br_0_249 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c249
+ bl_0_249 br_0_249 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c249
+ bl_0_249 br_0_249 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c249
+ bl_0_249 br_0_249 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c249
+ bl_0_249 br_0_249 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c249
+ bl_0_249 br_0_249 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c249
+ bl_0_249 br_0_249 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c249
+ bl_0_249 br_0_249 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c249
+ bl_0_249 br_0_249 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c249
+ bl_0_249 br_0_249 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c249
+ bl_0_249 br_0_249 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c249
+ bl_0_249 br_0_249 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c249
+ bl_0_249 br_0_249 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c249
+ bl_0_249 br_0_249 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c249
+ bl_0_249 br_0_249 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c249
+ bl_0_249 br_0_249 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c249
+ bl_0_249 br_0_249 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c249
+ bl_0_249 br_0_249 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c249
+ bl_0_249 br_0_249 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c249
+ bl_0_249 br_0_249 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c249
+ bl_0_249 br_0_249 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c249
+ bl_0_249 br_0_249 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c249
+ bl_0_249 br_0_249 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c250
+ bl_0_250 br_0_250 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c250
+ bl_0_250 br_0_250 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c250
+ bl_0_250 br_0_250 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c250
+ bl_0_250 br_0_250 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c250
+ bl_0_250 br_0_250 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c250
+ bl_0_250 br_0_250 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c250
+ bl_0_250 br_0_250 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c250
+ bl_0_250 br_0_250 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c250
+ bl_0_250 br_0_250 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c250
+ bl_0_250 br_0_250 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c250
+ bl_0_250 br_0_250 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c250
+ bl_0_250 br_0_250 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c250
+ bl_0_250 br_0_250 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c250
+ bl_0_250 br_0_250 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c250
+ bl_0_250 br_0_250 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c250
+ bl_0_250 br_0_250 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c250
+ bl_0_250 br_0_250 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c250
+ bl_0_250 br_0_250 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c250
+ bl_0_250 br_0_250 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c250
+ bl_0_250 br_0_250 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c250
+ bl_0_250 br_0_250 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c250
+ bl_0_250 br_0_250 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c250
+ bl_0_250 br_0_250 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c250
+ bl_0_250 br_0_250 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c250
+ bl_0_250 br_0_250 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c250
+ bl_0_250 br_0_250 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c250
+ bl_0_250 br_0_250 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c250
+ bl_0_250 br_0_250 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c250
+ bl_0_250 br_0_250 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c250
+ bl_0_250 br_0_250 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c250
+ bl_0_250 br_0_250 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c250
+ bl_0_250 br_0_250 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c250
+ bl_0_250 br_0_250 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c250
+ bl_0_250 br_0_250 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c250
+ bl_0_250 br_0_250 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c250
+ bl_0_250 br_0_250 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c250
+ bl_0_250 br_0_250 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c250
+ bl_0_250 br_0_250 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c250
+ bl_0_250 br_0_250 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c250
+ bl_0_250 br_0_250 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c250
+ bl_0_250 br_0_250 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c250
+ bl_0_250 br_0_250 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c250
+ bl_0_250 br_0_250 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c250
+ bl_0_250 br_0_250 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c251
+ bl_0_251 br_0_251 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c251
+ bl_0_251 br_0_251 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c251
+ bl_0_251 br_0_251 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c251
+ bl_0_251 br_0_251 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c251
+ bl_0_251 br_0_251 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c251
+ bl_0_251 br_0_251 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c251
+ bl_0_251 br_0_251 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c251
+ bl_0_251 br_0_251 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c251
+ bl_0_251 br_0_251 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c251
+ bl_0_251 br_0_251 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c251
+ bl_0_251 br_0_251 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c251
+ bl_0_251 br_0_251 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c251
+ bl_0_251 br_0_251 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c251
+ bl_0_251 br_0_251 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c251
+ bl_0_251 br_0_251 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c251
+ bl_0_251 br_0_251 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c251
+ bl_0_251 br_0_251 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c251
+ bl_0_251 br_0_251 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c251
+ bl_0_251 br_0_251 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c251
+ bl_0_251 br_0_251 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c251
+ bl_0_251 br_0_251 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c251
+ bl_0_251 br_0_251 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c251
+ bl_0_251 br_0_251 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c251
+ bl_0_251 br_0_251 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c251
+ bl_0_251 br_0_251 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c251
+ bl_0_251 br_0_251 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c251
+ bl_0_251 br_0_251 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c251
+ bl_0_251 br_0_251 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c251
+ bl_0_251 br_0_251 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c251
+ bl_0_251 br_0_251 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c251
+ bl_0_251 br_0_251 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c251
+ bl_0_251 br_0_251 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c251
+ bl_0_251 br_0_251 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c251
+ bl_0_251 br_0_251 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c251
+ bl_0_251 br_0_251 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c251
+ bl_0_251 br_0_251 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c251
+ bl_0_251 br_0_251 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c251
+ bl_0_251 br_0_251 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c251
+ bl_0_251 br_0_251 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c251
+ bl_0_251 br_0_251 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c251
+ bl_0_251 br_0_251 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c251
+ bl_0_251 br_0_251 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c251
+ bl_0_251 br_0_251 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c251
+ bl_0_251 br_0_251 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c252
+ bl_0_252 br_0_252 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c252
+ bl_0_252 br_0_252 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c252
+ bl_0_252 br_0_252 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c252
+ bl_0_252 br_0_252 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c252
+ bl_0_252 br_0_252 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c252
+ bl_0_252 br_0_252 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c252
+ bl_0_252 br_0_252 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c252
+ bl_0_252 br_0_252 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c252
+ bl_0_252 br_0_252 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c252
+ bl_0_252 br_0_252 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c252
+ bl_0_252 br_0_252 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c252
+ bl_0_252 br_0_252 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c252
+ bl_0_252 br_0_252 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c252
+ bl_0_252 br_0_252 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c252
+ bl_0_252 br_0_252 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c252
+ bl_0_252 br_0_252 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c252
+ bl_0_252 br_0_252 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c252
+ bl_0_252 br_0_252 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c252
+ bl_0_252 br_0_252 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c252
+ bl_0_252 br_0_252 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c252
+ bl_0_252 br_0_252 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c252
+ bl_0_252 br_0_252 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c252
+ bl_0_252 br_0_252 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c252
+ bl_0_252 br_0_252 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c252
+ bl_0_252 br_0_252 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c252
+ bl_0_252 br_0_252 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c252
+ bl_0_252 br_0_252 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c252
+ bl_0_252 br_0_252 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c252
+ bl_0_252 br_0_252 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c252
+ bl_0_252 br_0_252 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c252
+ bl_0_252 br_0_252 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c252
+ bl_0_252 br_0_252 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c252
+ bl_0_252 br_0_252 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c252
+ bl_0_252 br_0_252 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c252
+ bl_0_252 br_0_252 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c252
+ bl_0_252 br_0_252 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c252
+ bl_0_252 br_0_252 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c252
+ bl_0_252 br_0_252 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c252
+ bl_0_252 br_0_252 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c252
+ bl_0_252 br_0_252 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c252
+ bl_0_252 br_0_252 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c252
+ bl_0_252 br_0_252 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c252
+ bl_0_252 br_0_252 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c252
+ bl_0_252 br_0_252 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c253
+ bl_0_253 br_0_253 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c253
+ bl_0_253 br_0_253 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c253
+ bl_0_253 br_0_253 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c253
+ bl_0_253 br_0_253 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c253
+ bl_0_253 br_0_253 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c253
+ bl_0_253 br_0_253 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c253
+ bl_0_253 br_0_253 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c253
+ bl_0_253 br_0_253 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c253
+ bl_0_253 br_0_253 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c253
+ bl_0_253 br_0_253 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c253
+ bl_0_253 br_0_253 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c253
+ bl_0_253 br_0_253 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c253
+ bl_0_253 br_0_253 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c253
+ bl_0_253 br_0_253 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c253
+ bl_0_253 br_0_253 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c253
+ bl_0_253 br_0_253 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c253
+ bl_0_253 br_0_253 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c253
+ bl_0_253 br_0_253 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c253
+ bl_0_253 br_0_253 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c253
+ bl_0_253 br_0_253 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c253
+ bl_0_253 br_0_253 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c253
+ bl_0_253 br_0_253 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c253
+ bl_0_253 br_0_253 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c253
+ bl_0_253 br_0_253 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c253
+ bl_0_253 br_0_253 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c253
+ bl_0_253 br_0_253 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c253
+ bl_0_253 br_0_253 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c253
+ bl_0_253 br_0_253 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c253
+ bl_0_253 br_0_253 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c253
+ bl_0_253 br_0_253 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c253
+ bl_0_253 br_0_253 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c253
+ bl_0_253 br_0_253 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c253
+ bl_0_253 br_0_253 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c253
+ bl_0_253 br_0_253 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c253
+ bl_0_253 br_0_253 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c253
+ bl_0_253 br_0_253 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c253
+ bl_0_253 br_0_253 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c253
+ bl_0_253 br_0_253 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c253
+ bl_0_253 br_0_253 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c253
+ bl_0_253 br_0_253 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c253
+ bl_0_253 br_0_253 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c253
+ bl_0_253 br_0_253 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c253
+ bl_0_253 br_0_253 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c253
+ bl_0_253 br_0_253 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c254
+ bl_0_254 br_0_254 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c254
+ bl_0_254 br_0_254 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c254
+ bl_0_254 br_0_254 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c254
+ bl_0_254 br_0_254 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c254
+ bl_0_254 br_0_254 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c254
+ bl_0_254 br_0_254 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c254
+ bl_0_254 br_0_254 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c254
+ bl_0_254 br_0_254 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c254
+ bl_0_254 br_0_254 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c254
+ bl_0_254 br_0_254 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c254
+ bl_0_254 br_0_254 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c254
+ bl_0_254 br_0_254 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c254
+ bl_0_254 br_0_254 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c254
+ bl_0_254 br_0_254 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c254
+ bl_0_254 br_0_254 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c254
+ bl_0_254 br_0_254 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c254
+ bl_0_254 br_0_254 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c254
+ bl_0_254 br_0_254 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c254
+ bl_0_254 br_0_254 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c254
+ bl_0_254 br_0_254 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c254
+ bl_0_254 br_0_254 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c254
+ bl_0_254 br_0_254 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c254
+ bl_0_254 br_0_254 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c254
+ bl_0_254 br_0_254 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c254
+ bl_0_254 br_0_254 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c254
+ bl_0_254 br_0_254 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c254
+ bl_0_254 br_0_254 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c254
+ bl_0_254 br_0_254 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c254
+ bl_0_254 br_0_254 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c254
+ bl_0_254 br_0_254 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c254
+ bl_0_254 br_0_254 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c254
+ bl_0_254 br_0_254 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c254
+ bl_0_254 br_0_254 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c254
+ bl_0_254 br_0_254 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c254
+ bl_0_254 br_0_254 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c254
+ bl_0_254 br_0_254 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c254
+ bl_0_254 br_0_254 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c254
+ bl_0_254 br_0_254 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c254
+ bl_0_254 br_0_254 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c254
+ bl_0_254 br_0_254 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c254
+ bl_0_254 br_0_254 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c254
+ bl_0_254 br_0_254 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c254
+ bl_0_254 br_0_254 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c254
+ bl_0_254 br_0_254 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c255
+ bl_0_255 br_0_255 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c255
+ bl_0_255 br_0_255 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c255
+ bl_0_255 br_0_255 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c255
+ bl_0_255 br_0_255 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c255
+ bl_0_255 br_0_255 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c255
+ bl_0_255 br_0_255 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c255
+ bl_0_255 br_0_255 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c255
+ bl_0_255 br_0_255 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c255
+ bl_0_255 br_0_255 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c255
+ bl_0_255 br_0_255 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c255
+ bl_0_255 br_0_255 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c255
+ bl_0_255 br_0_255 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c255
+ bl_0_255 br_0_255 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c255
+ bl_0_255 br_0_255 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c255
+ bl_0_255 br_0_255 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c255
+ bl_0_255 br_0_255 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c255
+ bl_0_255 br_0_255 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c255
+ bl_0_255 br_0_255 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c255
+ bl_0_255 br_0_255 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c255
+ bl_0_255 br_0_255 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c255
+ bl_0_255 br_0_255 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c255
+ bl_0_255 br_0_255 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c255
+ bl_0_255 br_0_255 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c255
+ bl_0_255 br_0_255 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c255
+ bl_0_255 br_0_255 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c255
+ bl_0_255 br_0_255 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c255
+ bl_0_255 br_0_255 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c255
+ bl_0_255 br_0_255 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c255
+ bl_0_255 br_0_255 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c255
+ bl_0_255 br_0_255 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c255
+ bl_0_255 br_0_255 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c255
+ bl_0_255 br_0_255 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c255
+ bl_0_255 br_0_255 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c255
+ bl_0_255 br_0_255 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c255
+ bl_0_255 br_0_255 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c255
+ bl_0_255 br_0_255 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c255
+ bl_0_255 br_0_255 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c255
+ bl_0_255 br_0_255 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c255
+ bl_0_255 br_0_255 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c255
+ bl_0_255 br_0_255 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c255
+ bl_0_255 br_0_255 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c255
+ bl_0_255 br_0_255 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c255
+ bl_0_255 br_0_255 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c255
+ bl_0_255 br_0_255 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c256
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c256
+ bl_0_256 br_0_256 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c256
+ bl_0_256 br_0_256 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c256
+ bl_0_256 br_0_256 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c256
+ bl_0_256 br_0_256 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c256
+ bl_0_256 br_0_256 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c256
+ bl_0_256 br_0_256 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c256
+ bl_0_256 br_0_256 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c256
+ bl_0_256 br_0_256 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c256
+ bl_0_256 br_0_256 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c256
+ bl_0_256 br_0_256 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c256
+ bl_0_256 br_0_256 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c256
+ bl_0_256 br_0_256 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c256
+ bl_0_256 br_0_256 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c256
+ bl_0_256 br_0_256 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c256
+ bl_0_256 br_0_256 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c256
+ bl_0_256 br_0_256 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c256
+ bl_0_256 br_0_256 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c256
+ bl_0_256 br_0_256 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c256
+ bl_0_256 br_0_256 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c256
+ bl_0_256 br_0_256 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c256
+ bl_0_256 br_0_256 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c256
+ bl_0_256 br_0_256 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c256
+ bl_0_256 br_0_256 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c256
+ bl_0_256 br_0_256 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c256
+ bl_0_256 br_0_256 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c256
+ bl_0_256 br_0_256 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c256
+ bl_0_256 br_0_256 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c256
+ bl_0_256 br_0_256 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c256
+ bl_0_256 br_0_256 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c256
+ bl_0_256 br_0_256 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c256
+ bl_0_256 br_0_256 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c256
+ bl_0_256 br_0_256 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c256
+ bl_0_256 br_0_256 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c256
+ bl_0_256 br_0_256 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c256
+ bl_0_256 br_0_256 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c256
+ bl_0_256 br_0_256 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c256
+ bl_0_256 br_0_256 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c256
+ bl_0_256 br_0_256 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c256
+ bl_0_256 br_0_256 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c256
+ bl_0_256 br_0_256 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c256
+ bl_0_256 br_0_256 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c256
+ bl_0_256 br_0_256 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c256
+ bl_0_256 br_0_256 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c256
+ bl_0_256 br_0_256 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c257
+ bl_0_257 br_0_257 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c257
+ bl_0_257 br_0_257 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c257
+ bl_0_257 br_0_257 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c257
+ bl_0_257 br_0_257 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c257
+ bl_0_257 br_0_257 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c257
+ bl_0_257 br_0_257 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c257
+ bl_0_257 br_0_257 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c257
+ bl_0_257 br_0_257 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c257
+ bl_0_257 br_0_257 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c257
+ bl_0_257 br_0_257 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c257
+ bl_0_257 br_0_257 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c257
+ bl_0_257 br_0_257 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c257
+ bl_0_257 br_0_257 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c257
+ bl_0_257 br_0_257 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c257
+ bl_0_257 br_0_257 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c257
+ bl_0_257 br_0_257 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c257
+ bl_0_257 br_0_257 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c257
+ bl_0_257 br_0_257 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c257
+ bl_0_257 br_0_257 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c257
+ bl_0_257 br_0_257 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c257
+ bl_0_257 br_0_257 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c257
+ bl_0_257 br_0_257 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c257
+ bl_0_257 br_0_257 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c257
+ bl_0_257 br_0_257 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c257
+ bl_0_257 br_0_257 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c257
+ bl_0_257 br_0_257 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c257
+ bl_0_257 br_0_257 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c257
+ bl_0_257 br_0_257 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c257
+ bl_0_257 br_0_257 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c257
+ bl_0_257 br_0_257 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c257
+ bl_0_257 br_0_257 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c257
+ bl_0_257 br_0_257 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c257
+ bl_0_257 br_0_257 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c257
+ bl_0_257 br_0_257 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c257
+ bl_0_257 br_0_257 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c257
+ bl_0_257 br_0_257 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c257
+ bl_0_257 br_0_257 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c257
+ bl_0_257 br_0_257 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c257
+ bl_0_257 br_0_257 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c257
+ bl_0_257 br_0_257 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c257
+ bl_0_257 br_0_257 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c257
+ bl_0_257 br_0_257 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c257
+ bl_0_257 br_0_257 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c257
+ bl_0_257 br_0_257 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c257
+ bl_0_257 br_0_257 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c258
+ bl_0_258 br_0_258 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c258
+ bl_0_258 br_0_258 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c258
+ bl_0_258 br_0_258 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c258
+ bl_0_258 br_0_258 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c258
+ bl_0_258 br_0_258 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c258
+ bl_0_258 br_0_258 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c258
+ bl_0_258 br_0_258 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c258
+ bl_0_258 br_0_258 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c258
+ bl_0_258 br_0_258 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c258
+ bl_0_258 br_0_258 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c258
+ bl_0_258 br_0_258 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c258
+ bl_0_258 br_0_258 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c258
+ bl_0_258 br_0_258 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c258
+ bl_0_258 br_0_258 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c258
+ bl_0_258 br_0_258 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c258
+ bl_0_258 br_0_258 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c258
+ bl_0_258 br_0_258 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c258
+ bl_0_258 br_0_258 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c258
+ bl_0_258 br_0_258 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c258
+ bl_0_258 br_0_258 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c258
+ bl_0_258 br_0_258 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c258
+ bl_0_258 br_0_258 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c258
+ bl_0_258 br_0_258 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c258
+ bl_0_258 br_0_258 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c258
+ bl_0_258 br_0_258 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c258
+ bl_0_258 br_0_258 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c258
+ bl_0_258 br_0_258 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c258
+ bl_0_258 br_0_258 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c258
+ bl_0_258 br_0_258 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c258
+ bl_0_258 br_0_258 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c258
+ bl_0_258 br_0_258 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c258
+ bl_0_258 br_0_258 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c258
+ bl_0_258 br_0_258 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c258
+ bl_0_258 br_0_258 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c258
+ bl_0_258 br_0_258 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c258
+ bl_0_258 br_0_258 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c258
+ bl_0_258 br_0_258 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c258
+ bl_0_258 br_0_258 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c258
+ bl_0_258 br_0_258 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c258
+ bl_0_258 br_0_258 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c258
+ bl_0_258 br_0_258 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c258
+ bl_0_258 br_0_258 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c258
+ bl_0_258 br_0_258 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c258
+ bl_0_258 br_0_258 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c258
+ bl_0_258 br_0_258 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c259
+ bl_0_259 br_0_259 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c259
+ bl_0_259 br_0_259 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c259
+ bl_0_259 br_0_259 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c259
+ bl_0_259 br_0_259 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c259
+ bl_0_259 br_0_259 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c259
+ bl_0_259 br_0_259 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c259
+ bl_0_259 br_0_259 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c259
+ bl_0_259 br_0_259 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c259
+ bl_0_259 br_0_259 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c259
+ bl_0_259 br_0_259 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c259
+ bl_0_259 br_0_259 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c259
+ bl_0_259 br_0_259 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c259
+ bl_0_259 br_0_259 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c259
+ bl_0_259 br_0_259 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c259
+ bl_0_259 br_0_259 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c259
+ bl_0_259 br_0_259 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c259
+ bl_0_259 br_0_259 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c259
+ bl_0_259 br_0_259 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c259
+ bl_0_259 br_0_259 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c259
+ bl_0_259 br_0_259 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c259
+ bl_0_259 br_0_259 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c259
+ bl_0_259 br_0_259 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c259
+ bl_0_259 br_0_259 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c259
+ bl_0_259 br_0_259 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c259
+ bl_0_259 br_0_259 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c259
+ bl_0_259 br_0_259 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c259
+ bl_0_259 br_0_259 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c259
+ bl_0_259 br_0_259 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c259
+ bl_0_259 br_0_259 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c259
+ bl_0_259 br_0_259 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c259
+ bl_0_259 br_0_259 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c259
+ bl_0_259 br_0_259 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c259
+ bl_0_259 br_0_259 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c259
+ bl_0_259 br_0_259 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c259
+ bl_0_259 br_0_259 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c259
+ bl_0_259 br_0_259 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c259
+ bl_0_259 br_0_259 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c259
+ bl_0_259 br_0_259 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c259
+ bl_0_259 br_0_259 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c259
+ bl_0_259 br_0_259 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c259
+ bl_0_259 br_0_259 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c259
+ bl_0_259 br_0_259 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c259
+ bl_0_259 br_0_259 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c259
+ bl_0_259 br_0_259 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c259
+ bl_0_259 br_0_259 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c260
+ bl_0_260 br_0_260 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c260
+ bl_0_260 br_0_260 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c260
+ bl_0_260 br_0_260 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c260
+ bl_0_260 br_0_260 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c260
+ bl_0_260 br_0_260 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c260
+ bl_0_260 br_0_260 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c260
+ bl_0_260 br_0_260 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c260
+ bl_0_260 br_0_260 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c260
+ bl_0_260 br_0_260 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c260
+ bl_0_260 br_0_260 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c260
+ bl_0_260 br_0_260 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c260
+ bl_0_260 br_0_260 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c260
+ bl_0_260 br_0_260 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c260
+ bl_0_260 br_0_260 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c260
+ bl_0_260 br_0_260 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c260
+ bl_0_260 br_0_260 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c260
+ bl_0_260 br_0_260 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c260
+ bl_0_260 br_0_260 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c260
+ bl_0_260 br_0_260 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c260
+ bl_0_260 br_0_260 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c260
+ bl_0_260 br_0_260 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c260
+ bl_0_260 br_0_260 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c260
+ bl_0_260 br_0_260 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c260
+ bl_0_260 br_0_260 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c260
+ bl_0_260 br_0_260 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c260
+ bl_0_260 br_0_260 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c260
+ bl_0_260 br_0_260 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c260
+ bl_0_260 br_0_260 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c260
+ bl_0_260 br_0_260 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c260
+ bl_0_260 br_0_260 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c260
+ bl_0_260 br_0_260 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c260
+ bl_0_260 br_0_260 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c260
+ bl_0_260 br_0_260 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c260
+ bl_0_260 br_0_260 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c260
+ bl_0_260 br_0_260 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c260
+ bl_0_260 br_0_260 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c260
+ bl_0_260 br_0_260 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c260
+ bl_0_260 br_0_260 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c260
+ bl_0_260 br_0_260 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c260
+ bl_0_260 br_0_260 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c260
+ bl_0_260 br_0_260 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c260
+ bl_0_260 br_0_260 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c260
+ bl_0_260 br_0_260 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c260
+ bl_0_260 br_0_260 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c260
+ bl_0_260 br_0_260 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c261
+ bl_0_261 br_0_261 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c261
+ bl_0_261 br_0_261 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c261
+ bl_0_261 br_0_261 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c261
+ bl_0_261 br_0_261 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c261
+ bl_0_261 br_0_261 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c261
+ bl_0_261 br_0_261 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c261
+ bl_0_261 br_0_261 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c261
+ bl_0_261 br_0_261 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c261
+ bl_0_261 br_0_261 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c261
+ bl_0_261 br_0_261 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c261
+ bl_0_261 br_0_261 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c261
+ bl_0_261 br_0_261 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c261
+ bl_0_261 br_0_261 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c261
+ bl_0_261 br_0_261 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c261
+ bl_0_261 br_0_261 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c261
+ bl_0_261 br_0_261 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c261
+ bl_0_261 br_0_261 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c261
+ bl_0_261 br_0_261 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c261
+ bl_0_261 br_0_261 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c261
+ bl_0_261 br_0_261 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c261
+ bl_0_261 br_0_261 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c261
+ bl_0_261 br_0_261 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c261
+ bl_0_261 br_0_261 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c261
+ bl_0_261 br_0_261 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c261
+ bl_0_261 br_0_261 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c261
+ bl_0_261 br_0_261 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c261
+ bl_0_261 br_0_261 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c261
+ bl_0_261 br_0_261 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c261
+ bl_0_261 br_0_261 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c261
+ bl_0_261 br_0_261 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c261
+ bl_0_261 br_0_261 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c261
+ bl_0_261 br_0_261 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c261
+ bl_0_261 br_0_261 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c261
+ bl_0_261 br_0_261 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c261
+ bl_0_261 br_0_261 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c261
+ bl_0_261 br_0_261 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c261
+ bl_0_261 br_0_261 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c261
+ bl_0_261 br_0_261 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c261
+ bl_0_261 br_0_261 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c261
+ bl_0_261 br_0_261 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c261
+ bl_0_261 br_0_261 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c261
+ bl_0_261 br_0_261 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c261
+ bl_0_261 br_0_261 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c261
+ bl_0_261 br_0_261 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c261
+ bl_0_261 br_0_261 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c262
+ bl_0_262 br_0_262 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c262
+ bl_0_262 br_0_262 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c262
+ bl_0_262 br_0_262 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c262
+ bl_0_262 br_0_262 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c262
+ bl_0_262 br_0_262 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c262
+ bl_0_262 br_0_262 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c262
+ bl_0_262 br_0_262 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c262
+ bl_0_262 br_0_262 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c262
+ bl_0_262 br_0_262 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c262
+ bl_0_262 br_0_262 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c262
+ bl_0_262 br_0_262 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c262
+ bl_0_262 br_0_262 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c262
+ bl_0_262 br_0_262 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c262
+ bl_0_262 br_0_262 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c262
+ bl_0_262 br_0_262 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c262
+ bl_0_262 br_0_262 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c262
+ bl_0_262 br_0_262 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c262
+ bl_0_262 br_0_262 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c262
+ bl_0_262 br_0_262 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c262
+ bl_0_262 br_0_262 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c262
+ bl_0_262 br_0_262 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c262
+ bl_0_262 br_0_262 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c262
+ bl_0_262 br_0_262 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c262
+ bl_0_262 br_0_262 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c262
+ bl_0_262 br_0_262 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c262
+ bl_0_262 br_0_262 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c262
+ bl_0_262 br_0_262 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c262
+ bl_0_262 br_0_262 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c262
+ bl_0_262 br_0_262 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c262
+ bl_0_262 br_0_262 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c262
+ bl_0_262 br_0_262 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c262
+ bl_0_262 br_0_262 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c262
+ bl_0_262 br_0_262 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c262
+ bl_0_262 br_0_262 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c262
+ bl_0_262 br_0_262 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c262
+ bl_0_262 br_0_262 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c262
+ bl_0_262 br_0_262 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c262
+ bl_0_262 br_0_262 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c262
+ bl_0_262 br_0_262 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c262
+ bl_0_262 br_0_262 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c262
+ bl_0_262 br_0_262 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c262
+ bl_0_262 br_0_262 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c262
+ bl_0_262 br_0_262 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c262
+ bl_0_262 br_0_262 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c262
+ bl_0_262 br_0_262 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c263
+ bl_0_263 br_0_263 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c263
+ bl_0_263 br_0_263 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c263
+ bl_0_263 br_0_263 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c263
+ bl_0_263 br_0_263 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c263
+ bl_0_263 br_0_263 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c263
+ bl_0_263 br_0_263 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c263
+ bl_0_263 br_0_263 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c263
+ bl_0_263 br_0_263 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c263
+ bl_0_263 br_0_263 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c263
+ bl_0_263 br_0_263 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c263
+ bl_0_263 br_0_263 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c263
+ bl_0_263 br_0_263 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c263
+ bl_0_263 br_0_263 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c263
+ bl_0_263 br_0_263 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c263
+ bl_0_263 br_0_263 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c263
+ bl_0_263 br_0_263 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c263
+ bl_0_263 br_0_263 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c263
+ bl_0_263 br_0_263 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c263
+ bl_0_263 br_0_263 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c263
+ bl_0_263 br_0_263 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c263
+ bl_0_263 br_0_263 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c263
+ bl_0_263 br_0_263 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c263
+ bl_0_263 br_0_263 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c263
+ bl_0_263 br_0_263 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c263
+ bl_0_263 br_0_263 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c263
+ bl_0_263 br_0_263 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c263
+ bl_0_263 br_0_263 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c263
+ bl_0_263 br_0_263 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c263
+ bl_0_263 br_0_263 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c263
+ bl_0_263 br_0_263 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c263
+ bl_0_263 br_0_263 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c263
+ bl_0_263 br_0_263 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c263
+ bl_0_263 br_0_263 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c263
+ bl_0_263 br_0_263 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c263
+ bl_0_263 br_0_263 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c263
+ bl_0_263 br_0_263 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c263
+ bl_0_263 br_0_263 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c263
+ bl_0_263 br_0_263 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c263
+ bl_0_263 br_0_263 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c263
+ bl_0_263 br_0_263 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c263
+ bl_0_263 br_0_263 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c263
+ bl_0_263 br_0_263 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c263
+ bl_0_263 br_0_263 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c263
+ bl_0_263 br_0_263 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c263
+ bl_0_263 br_0_263 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c264
+ bl_0_264 br_0_264 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c264
+ bl_0_264 br_0_264 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c264
+ bl_0_264 br_0_264 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c264
+ bl_0_264 br_0_264 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c264
+ bl_0_264 br_0_264 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c264
+ bl_0_264 br_0_264 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c264
+ bl_0_264 br_0_264 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c264
+ bl_0_264 br_0_264 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c264
+ bl_0_264 br_0_264 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c264
+ bl_0_264 br_0_264 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c264
+ bl_0_264 br_0_264 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c264
+ bl_0_264 br_0_264 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c264
+ bl_0_264 br_0_264 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c264
+ bl_0_264 br_0_264 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c264
+ bl_0_264 br_0_264 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c264
+ bl_0_264 br_0_264 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c264
+ bl_0_264 br_0_264 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c264
+ bl_0_264 br_0_264 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c264
+ bl_0_264 br_0_264 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c264
+ bl_0_264 br_0_264 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c264
+ bl_0_264 br_0_264 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c264
+ bl_0_264 br_0_264 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c264
+ bl_0_264 br_0_264 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c264
+ bl_0_264 br_0_264 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c264
+ bl_0_264 br_0_264 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c264
+ bl_0_264 br_0_264 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c264
+ bl_0_264 br_0_264 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c264
+ bl_0_264 br_0_264 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c264
+ bl_0_264 br_0_264 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c264
+ bl_0_264 br_0_264 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c264
+ bl_0_264 br_0_264 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c264
+ bl_0_264 br_0_264 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c264
+ bl_0_264 br_0_264 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c264
+ bl_0_264 br_0_264 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c264
+ bl_0_264 br_0_264 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c264
+ bl_0_264 br_0_264 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c264
+ bl_0_264 br_0_264 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c264
+ bl_0_264 br_0_264 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c264
+ bl_0_264 br_0_264 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c264
+ bl_0_264 br_0_264 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c264
+ bl_0_264 br_0_264 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c264
+ bl_0_264 br_0_264 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c264
+ bl_0_264 br_0_264 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c264
+ bl_0_264 br_0_264 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c264
+ bl_0_264 br_0_264 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c265
+ bl_0_265 br_0_265 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c265
+ bl_0_265 br_0_265 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c265
+ bl_0_265 br_0_265 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c265
+ bl_0_265 br_0_265 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c265
+ bl_0_265 br_0_265 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c265
+ bl_0_265 br_0_265 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c265
+ bl_0_265 br_0_265 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c265
+ bl_0_265 br_0_265 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c265
+ bl_0_265 br_0_265 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c265
+ bl_0_265 br_0_265 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c265
+ bl_0_265 br_0_265 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c265
+ bl_0_265 br_0_265 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c265
+ bl_0_265 br_0_265 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c265
+ bl_0_265 br_0_265 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c265
+ bl_0_265 br_0_265 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c265
+ bl_0_265 br_0_265 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c265
+ bl_0_265 br_0_265 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c265
+ bl_0_265 br_0_265 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c265
+ bl_0_265 br_0_265 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c265
+ bl_0_265 br_0_265 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c265
+ bl_0_265 br_0_265 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c265
+ bl_0_265 br_0_265 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c265
+ bl_0_265 br_0_265 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c265
+ bl_0_265 br_0_265 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c265
+ bl_0_265 br_0_265 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c265
+ bl_0_265 br_0_265 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c265
+ bl_0_265 br_0_265 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c265
+ bl_0_265 br_0_265 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c265
+ bl_0_265 br_0_265 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c265
+ bl_0_265 br_0_265 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c265
+ bl_0_265 br_0_265 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c265
+ bl_0_265 br_0_265 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c265
+ bl_0_265 br_0_265 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c265
+ bl_0_265 br_0_265 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c265
+ bl_0_265 br_0_265 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c265
+ bl_0_265 br_0_265 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c265
+ bl_0_265 br_0_265 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c265
+ bl_0_265 br_0_265 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c265
+ bl_0_265 br_0_265 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c265
+ bl_0_265 br_0_265 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c265
+ bl_0_265 br_0_265 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c265
+ bl_0_265 br_0_265 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c265
+ bl_0_265 br_0_265 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c265
+ bl_0_265 br_0_265 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c265
+ bl_0_265 br_0_265 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c266
+ bl_0_266 br_0_266 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c266
+ bl_0_266 br_0_266 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c266
+ bl_0_266 br_0_266 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c266
+ bl_0_266 br_0_266 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c266
+ bl_0_266 br_0_266 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c266
+ bl_0_266 br_0_266 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c266
+ bl_0_266 br_0_266 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c266
+ bl_0_266 br_0_266 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c266
+ bl_0_266 br_0_266 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c266
+ bl_0_266 br_0_266 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c266
+ bl_0_266 br_0_266 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c266
+ bl_0_266 br_0_266 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c266
+ bl_0_266 br_0_266 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c266
+ bl_0_266 br_0_266 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c266
+ bl_0_266 br_0_266 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c266
+ bl_0_266 br_0_266 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c266
+ bl_0_266 br_0_266 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c266
+ bl_0_266 br_0_266 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c266
+ bl_0_266 br_0_266 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c266
+ bl_0_266 br_0_266 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c266
+ bl_0_266 br_0_266 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c266
+ bl_0_266 br_0_266 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c266
+ bl_0_266 br_0_266 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c266
+ bl_0_266 br_0_266 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c266
+ bl_0_266 br_0_266 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c266
+ bl_0_266 br_0_266 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c266
+ bl_0_266 br_0_266 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c266
+ bl_0_266 br_0_266 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c266
+ bl_0_266 br_0_266 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c266
+ bl_0_266 br_0_266 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c266
+ bl_0_266 br_0_266 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c266
+ bl_0_266 br_0_266 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c266
+ bl_0_266 br_0_266 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c266
+ bl_0_266 br_0_266 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c266
+ bl_0_266 br_0_266 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c266
+ bl_0_266 br_0_266 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c266
+ bl_0_266 br_0_266 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c266
+ bl_0_266 br_0_266 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c266
+ bl_0_266 br_0_266 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c266
+ bl_0_266 br_0_266 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c266
+ bl_0_266 br_0_266 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c266
+ bl_0_266 br_0_266 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c266
+ bl_0_266 br_0_266 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c266
+ bl_0_266 br_0_266 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c266
+ bl_0_266 br_0_266 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c267
+ bl_0_267 br_0_267 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c267
+ bl_0_267 br_0_267 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c267
+ bl_0_267 br_0_267 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c267
+ bl_0_267 br_0_267 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c267
+ bl_0_267 br_0_267 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c267
+ bl_0_267 br_0_267 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c267
+ bl_0_267 br_0_267 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c267
+ bl_0_267 br_0_267 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c267
+ bl_0_267 br_0_267 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c267
+ bl_0_267 br_0_267 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c267
+ bl_0_267 br_0_267 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c267
+ bl_0_267 br_0_267 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c267
+ bl_0_267 br_0_267 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c267
+ bl_0_267 br_0_267 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c267
+ bl_0_267 br_0_267 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c267
+ bl_0_267 br_0_267 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c267
+ bl_0_267 br_0_267 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c267
+ bl_0_267 br_0_267 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c267
+ bl_0_267 br_0_267 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c267
+ bl_0_267 br_0_267 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c267
+ bl_0_267 br_0_267 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c267
+ bl_0_267 br_0_267 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c267
+ bl_0_267 br_0_267 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c267
+ bl_0_267 br_0_267 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c267
+ bl_0_267 br_0_267 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c267
+ bl_0_267 br_0_267 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c267
+ bl_0_267 br_0_267 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c267
+ bl_0_267 br_0_267 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c267
+ bl_0_267 br_0_267 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c267
+ bl_0_267 br_0_267 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c267
+ bl_0_267 br_0_267 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c267
+ bl_0_267 br_0_267 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c267
+ bl_0_267 br_0_267 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c267
+ bl_0_267 br_0_267 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c267
+ bl_0_267 br_0_267 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c267
+ bl_0_267 br_0_267 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c267
+ bl_0_267 br_0_267 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c267
+ bl_0_267 br_0_267 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c267
+ bl_0_267 br_0_267 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c267
+ bl_0_267 br_0_267 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c267
+ bl_0_267 br_0_267 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c267
+ bl_0_267 br_0_267 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c267
+ bl_0_267 br_0_267 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c267
+ bl_0_267 br_0_267 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c267
+ bl_0_267 br_0_267 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c268
+ bl_0_268 br_0_268 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c268
+ bl_0_268 br_0_268 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c268
+ bl_0_268 br_0_268 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c268
+ bl_0_268 br_0_268 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c268
+ bl_0_268 br_0_268 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c268
+ bl_0_268 br_0_268 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c268
+ bl_0_268 br_0_268 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c268
+ bl_0_268 br_0_268 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c268
+ bl_0_268 br_0_268 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c268
+ bl_0_268 br_0_268 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c268
+ bl_0_268 br_0_268 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c268
+ bl_0_268 br_0_268 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c268
+ bl_0_268 br_0_268 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c268
+ bl_0_268 br_0_268 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c268
+ bl_0_268 br_0_268 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c268
+ bl_0_268 br_0_268 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c268
+ bl_0_268 br_0_268 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c268
+ bl_0_268 br_0_268 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c268
+ bl_0_268 br_0_268 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c268
+ bl_0_268 br_0_268 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c268
+ bl_0_268 br_0_268 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c268
+ bl_0_268 br_0_268 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c268
+ bl_0_268 br_0_268 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c268
+ bl_0_268 br_0_268 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c268
+ bl_0_268 br_0_268 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c268
+ bl_0_268 br_0_268 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c268
+ bl_0_268 br_0_268 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c268
+ bl_0_268 br_0_268 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c268
+ bl_0_268 br_0_268 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c268
+ bl_0_268 br_0_268 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c268
+ bl_0_268 br_0_268 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c268
+ bl_0_268 br_0_268 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c268
+ bl_0_268 br_0_268 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c268
+ bl_0_268 br_0_268 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c268
+ bl_0_268 br_0_268 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c268
+ bl_0_268 br_0_268 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c268
+ bl_0_268 br_0_268 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c268
+ bl_0_268 br_0_268 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c268
+ bl_0_268 br_0_268 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c268
+ bl_0_268 br_0_268 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c268
+ bl_0_268 br_0_268 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c268
+ bl_0_268 br_0_268 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c268
+ bl_0_268 br_0_268 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c268
+ bl_0_268 br_0_268 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c268
+ bl_0_268 br_0_268 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c269
+ bl_0_269 br_0_269 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c269
+ bl_0_269 br_0_269 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c269
+ bl_0_269 br_0_269 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c269
+ bl_0_269 br_0_269 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c269
+ bl_0_269 br_0_269 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c269
+ bl_0_269 br_0_269 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c269
+ bl_0_269 br_0_269 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c269
+ bl_0_269 br_0_269 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c269
+ bl_0_269 br_0_269 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c269
+ bl_0_269 br_0_269 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c269
+ bl_0_269 br_0_269 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c269
+ bl_0_269 br_0_269 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c269
+ bl_0_269 br_0_269 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c269
+ bl_0_269 br_0_269 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c269
+ bl_0_269 br_0_269 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c269
+ bl_0_269 br_0_269 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c269
+ bl_0_269 br_0_269 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c269
+ bl_0_269 br_0_269 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c269
+ bl_0_269 br_0_269 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c269
+ bl_0_269 br_0_269 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c269
+ bl_0_269 br_0_269 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c269
+ bl_0_269 br_0_269 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c269
+ bl_0_269 br_0_269 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c269
+ bl_0_269 br_0_269 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c269
+ bl_0_269 br_0_269 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c269
+ bl_0_269 br_0_269 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c269
+ bl_0_269 br_0_269 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c269
+ bl_0_269 br_0_269 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c269
+ bl_0_269 br_0_269 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c269
+ bl_0_269 br_0_269 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c269
+ bl_0_269 br_0_269 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c269
+ bl_0_269 br_0_269 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c269
+ bl_0_269 br_0_269 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c269
+ bl_0_269 br_0_269 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c269
+ bl_0_269 br_0_269 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c269
+ bl_0_269 br_0_269 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c269
+ bl_0_269 br_0_269 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c269
+ bl_0_269 br_0_269 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c269
+ bl_0_269 br_0_269 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c269
+ bl_0_269 br_0_269 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c269
+ bl_0_269 br_0_269 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c269
+ bl_0_269 br_0_269 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c269
+ bl_0_269 br_0_269 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c269
+ bl_0_269 br_0_269 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c269
+ bl_0_269 br_0_269 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c270
+ bl_0_270 br_0_270 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c270
+ bl_0_270 br_0_270 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c270
+ bl_0_270 br_0_270 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c270
+ bl_0_270 br_0_270 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c270
+ bl_0_270 br_0_270 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c270
+ bl_0_270 br_0_270 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c270
+ bl_0_270 br_0_270 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c270
+ bl_0_270 br_0_270 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c270
+ bl_0_270 br_0_270 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c270
+ bl_0_270 br_0_270 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c270
+ bl_0_270 br_0_270 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c270
+ bl_0_270 br_0_270 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c270
+ bl_0_270 br_0_270 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c270
+ bl_0_270 br_0_270 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c270
+ bl_0_270 br_0_270 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c270
+ bl_0_270 br_0_270 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c270
+ bl_0_270 br_0_270 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c270
+ bl_0_270 br_0_270 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c270
+ bl_0_270 br_0_270 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c270
+ bl_0_270 br_0_270 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c270
+ bl_0_270 br_0_270 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c270
+ bl_0_270 br_0_270 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c270
+ bl_0_270 br_0_270 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c270
+ bl_0_270 br_0_270 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c270
+ bl_0_270 br_0_270 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c270
+ bl_0_270 br_0_270 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c270
+ bl_0_270 br_0_270 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c270
+ bl_0_270 br_0_270 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c270
+ bl_0_270 br_0_270 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c270
+ bl_0_270 br_0_270 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c270
+ bl_0_270 br_0_270 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c270
+ bl_0_270 br_0_270 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c270
+ bl_0_270 br_0_270 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c270
+ bl_0_270 br_0_270 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c270
+ bl_0_270 br_0_270 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c270
+ bl_0_270 br_0_270 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c270
+ bl_0_270 br_0_270 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c270
+ bl_0_270 br_0_270 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c270
+ bl_0_270 br_0_270 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c270
+ bl_0_270 br_0_270 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c270
+ bl_0_270 br_0_270 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c270
+ bl_0_270 br_0_270 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c270
+ bl_0_270 br_0_270 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c270
+ bl_0_270 br_0_270 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c270
+ bl_0_270 br_0_270 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c271
+ bl_0_271 br_0_271 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c271
+ bl_0_271 br_0_271 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c271
+ bl_0_271 br_0_271 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c271
+ bl_0_271 br_0_271 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c271
+ bl_0_271 br_0_271 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c271
+ bl_0_271 br_0_271 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c271
+ bl_0_271 br_0_271 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c271
+ bl_0_271 br_0_271 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c271
+ bl_0_271 br_0_271 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c271
+ bl_0_271 br_0_271 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c271
+ bl_0_271 br_0_271 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c271
+ bl_0_271 br_0_271 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c271
+ bl_0_271 br_0_271 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c271
+ bl_0_271 br_0_271 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c271
+ bl_0_271 br_0_271 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c271
+ bl_0_271 br_0_271 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c271
+ bl_0_271 br_0_271 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c271
+ bl_0_271 br_0_271 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c271
+ bl_0_271 br_0_271 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c271
+ bl_0_271 br_0_271 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c271
+ bl_0_271 br_0_271 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c271
+ bl_0_271 br_0_271 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c271
+ bl_0_271 br_0_271 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c271
+ bl_0_271 br_0_271 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c271
+ bl_0_271 br_0_271 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c271
+ bl_0_271 br_0_271 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c271
+ bl_0_271 br_0_271 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c271
+ bl_0_271 br_0_271 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c271
+ bl_0_271 br_0_271 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c271
+ bl_0_271 br_0_271 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c271
+ bl_0_271 br_0_271 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c271
+ bl_0_271 br_0_271 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c271
+ bl_0_271 br_0_271 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c271
+ bl_0_271 br_0_271 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c271
+ bl_0_271 br_0_271 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c271
+ bl_0_271 br_0_271 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c271
+ bl_0_271 br_0_271 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c271
+ bl_0_271 br_0_271 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c271
+ bl_0_271 br_0_271 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c271
+ bl_0_271 br_0_271 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c271
+ bl_0_271 br_0_271 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c271
+ bl_0_271 br_0_271 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c271
+ bl_0_271 br_0_271 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c271
+ bl_0_271 br_0_271 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c271
+ bl_0_271 br_0_271 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c272
+ bl_0_272 br_0_272 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c272
+ bl_0_272 br_0_272 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c272
+ bl_0_272 br_0_272 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c272
+ bl_0_272 br_0_272 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c272
+ bl_0_272 br_0_272 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c272
+ bl_0_272 br_0_272 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c272
+ bl_0_272 br_0_272 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c272
+ bl_0_272 br_0_272 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c272
+ bl_0_272 br_0_272 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c272
+ bl_0_272 br_0_272 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c272
+ bl_0_272 br_0_272 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c272
+ bl_0_272 br_0_272 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c272
+ bl_0_272 br_0_272 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c272
+ bl_0_272 br_0_272 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c272
+ bl_0_272 br_0_272 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c272
+ bl_0_272 br_0_272 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c272
+ bl_0_272 br_0_272 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c272
+ bl_0_272 br_0_272 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c272
+ bl_0_272 br_0_272 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c272
+ bl_0_272 br_0_272 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c272
+ bl_0_272 br_0_272 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c272
+ bl_0_272 br_0_272 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c272
+ bl_0_272 br_0_272 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c272
+ bl_0_272 br_0_272 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c272
+ bl_0_272 br_0_272 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c272
+ bl_0_272 br_0_272 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c272
+ bl_0_272 br_0_272 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c272
+ bl_0_272 br_0_272 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c272
+ bl_0_272 br_0_272 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c272
+ bl_0_272 br_0_272 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c272
+ bl_0_272 br_0_272 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c272
+ bl_0_272 br_0_272 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c272
+ bl_0_272 br_0_272 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c272
+ bl_0_272 br_0_272 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c272
+ bl_0_272 br_0_272 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c272
+ bl_0_272 br_0_272 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c272
+ bl_0_272 br_0_272 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c272
+ bl_0_272 br_0_272 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c272
+ bl_0_272 br_0_272 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c272
+ bl_0_272 br_0_272 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c272
+ bl_0_272 br_0_272 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c272
+ bl_0_272 br_0_272 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c272
+ bl_0_272 br_0_272 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c272
+ bl_0_272 br_0_272 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c272
+ bl_0_272 br_0_272 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c273
+ bl_0_273 br_0_273 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c273
+ bl_0_273 br_0_273 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c273
+ bl_0_273 br_0_273 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c273
+ bl_0_273 br_0_273 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c273
+ bl_0_273 br_0_273 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c273
+ bl_0_273 br_0_273 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c273
+ bl_0_273 br_0_273 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c273
+ bl_0_273 br_0_273 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c273
+ bl_0_273 br_0_273 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c273
+ bl_0_273 br_0_273 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c273
+ bl_0_273 br_0_273 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c273
+ bl_0_273 br_0_273 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c273
+ bl_0_273 br_0_273 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c273
+ bl_0_273 br_0_273 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c273
+ bl_0_273 br_0_273 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c273
+ bl_0_273 br_0_273 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c273
+ bl_0_273 br_0_273 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c273
+ bl_0_273 br_0_273 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c273
+ bl_0_273 br_0_273 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c273
+ bl_0_273 br_0_273 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c273
+ bl_0_273 br_0_273 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c273
+ bl_0_273 br_0_273 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c273
+ bl_0_273 br_0_273 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c273
+ bl_0_273 br_0_273 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c273
+ bl_0_273 br_0_273 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c273
+ bl_0_273 br_0_273 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c273
+ bl_0_273 br_0_273 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c273
+ bl_0_273 br_0_273 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c273
+ bl_0_273 br_0_273 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c273
+ bl_0_273 br_0_273 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c273
+ bl_0_273 br_0_273 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c273
+ bl_0_273 br_0_273 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c273
+ bl_0_273 br_0_273 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c273
+ bl_0_273 br_0_273 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c273
+ bl_0_273 br_0_273 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c273
+ bl_0_273 br_0_273 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c273
+ bl_0_273 br_0_273 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c273
+ bl_0_273 br_0_273 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c273
+ bl_0_273 br_0_273 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c273
+ bl_0_273 br_0_273 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c273
+ bl_0_273 br_0_273 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c273
+ bl_0_273 br_0_273 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c273
+ bl_0_273 br_0_273 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c273
+ bl_0_273 br_0_273 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c273
+ bl_0_273 br_0_273 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c274
+ bl_0_274 br_0_274 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c274
+ bl_0_274 br_0_274 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c274
+ bl_0_274 br_0_274 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c274
+ bl_0_274 br_0_274 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c274
+ bl_0_274 br_0_274 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c274
+ bl_0_274 br_0_274 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c274
+ bl_0_274 br_0_274 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c274
+ bl_0_274 br_0_274 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c274
+ bl_0_274 br_0_274 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c274
+ bl_0_274 br_0_274 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c274
+ bl_0_274 br_0_274 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c274
+ bl_0_274 br_0_274 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c274
+ bl_0_274 br_0_274 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c274
+ bl_0_274 br_0_274 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c274
+ bl_0_274 br_0_274 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c274
+ bl_0_274 br_0_274 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c274
+ bl_0_274 br_0_274 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c274
+ bl_0_274 br_0_274 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c274
+ bl_0_274 br_0_274 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c274
+ bl_0_274 br_0_274 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c274
+ bl_0_274 br_0_274 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c274
+ bl_0_274 br_0_274 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c274
+ bl_0_274 br_0_274 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c274
+ bl_0_274 br_0_274 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c274
+ bl_0_274 br_0_274 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c274
+ bl_0_274 br_0_274 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c274
+ bl_0_274 br_0_274 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c274
+ bl_0_274 br_0_274 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c274
+ bl_0_274 br_0_274 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c274
+ bl_0_274 br_0_274 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c274
+ bl_0_274 br_0_274 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c274
+ bl_0_274 br_0_274 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c274
+ bl_0_274 br_0_274 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c274
+ bl_0_274 br_0_274 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c274
+ bl_0_274 br_0_274 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c274
+ bl_0_274 br_0_274 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c274
+ bl_0_274 br_0_274 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c274
+ bl_0_274 br_0_274 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c274
+ bl_0_274 br_0_274 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c274
+ bl_0_274 br_0_274 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c274
+ bl_0_274 br_0_274 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c274
+ bl_0_274 br_0_274 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c274
+ bl_0_274 br_0_274 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c274
+ bl_0_274 br_0_274 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c274
+ bl_0_274 br_0_274 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c275
+ bl_0_275 br_0_275 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c275
+ bl_0_275 br_0_275 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c275
+ bl_0_275 br_0_275 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c275
+ bl_0_275 br_0_275 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c275
+ bl_0_275 br_0_275 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c275
+ bl_0_275 br_0_275 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c275
+ bl_0_275 br_0_275 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c275
+ bl_0_275 br_0_275 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c275
+ bl_0_275 br_0_275 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c275
+ bl_0_275 br_0_275 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c275
+ bl_0_275 br_0_275 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c275
+ bl_0_275 br_0_275 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c275
+ bl_0_275 br_0_275 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c275
+ bl_0_275 br_0_275 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c275
+ bl_0_275 br_0_275 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c275
+ bl_0_275 br_0_275 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c275
+ bl_0_275 br_0_275 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c275
+ bl_0_275 br_0_275 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c275
+ bl_0_275 br_0_275 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c275
+ bl_0_275 br_0_275 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c275
+ bl_0_275 br_0_275 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c275
+ bl_0_275 br_0_275 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c275
+ bl_0_275 br_0_275 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c275
+ bl_0_275 br_0_275 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c275
+ bl_0_275 br_0_275 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c275
+ bl_0_275 br_0_275 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c275
+ bl_0_275 br_0_275 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c275
+ bl_0_275 br_0_275 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c275
+ bl_0_275 br_0_275 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c275
+ bl_0_275 br_0_275 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c275
+ bl_0_275 br_0_275 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c275
+ bl_0_275 br_0_275 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c275
+ bl_0_275 br_0_275 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c275
+ bl_0_275 br_0_275 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c275
+ bl_0_275 br_0_275 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c275
+ bl_0_275 br_0_275 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c275
+ bl_0_275 br_0_275 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c275
+ bl_0_275 br_0_275 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c275
+ bl_0_275 br_0_275 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c275
+ bl_0_275 br_0_275 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c275
+ bl_0_275 br_0_275 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c275
+ bl_0_275 br_0_275 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c275
+ bl_0_275 br_0_275 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c275
+ bl_0_275 br_0_275 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c275
+ bl_0_275 br_0_275 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c276
+ bl_0_276 br_0_276 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c276
+ bl_0_276 br_0_276 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c276
+ bl_0_276 br_0_276 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c276
+ bl_0_276 br_0_276 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c276
+ bl_0_276 br_0_276 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c276
+ bl_0_276 br_0_276 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c276
+ bl_0_276 br_0_276 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c276
+ bl_0_276 br_0_276 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c276
+ bl_0_276 br_0_276 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c276
+ bl_0_276 br_0_276 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c276
+ bl_0_276 br_0_276 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c276
+ bl_0_276 br_0_276 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c276
+ bl_0_276 br_0_276 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c276
+ bl_0_276 br_0_276 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c276
+ bl_0_276 br_0_276 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c276
+ bl_0_276 br_0_276 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c276
+ bl_0_276 br_0_276 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c276
+ bl_0_276 br_0_276 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c276
+ bl_0_276 br_0_276 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c276
+ bl_0_276 br_0_276 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c276
+ bl_0_276 br_0_276 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c276
+ bl_0_276 br_0_276 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c276
+ bl_0_276 br_0_276 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c276
+ bl_0_276 br_0_276 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c276
+ bl_0_276 br_0_276 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c276
+ bl_0_276 br_0_276 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c276
+ bl_0_276 br_0_276 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c276
+ bl_0_276 br_0_276 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c276
+ bl_0_276 br_0_276 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c276
+ bl_0_276 br_0_276 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c276
+ bl_0_276 br_0_276 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c276
+ bl_0_276 br_0_276 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c276
+ bl_0_276 br_0_276 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c276
+ bl_0_276 br_0_276 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c276
+ bl_0_276 br_0_276 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c276
+ bl_0_276 br_0_276 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c276
+ bl_0_276 br_0_276 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c276
+ bl_0_276 br_0_276 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c276
+ bl_0_276 br_0_276 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c276
+ bl_0_276 br_0_276 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c276
+ bl_0_276 br_0_276 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c276
+ bl_0_276 br_0_276 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c276
+ bl_0_276 br_0_276 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c276
+ bl_0_276 br_0_276 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c276
+ bl_0_276 br_0_276 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c277
+ bl_0_277 br_0_277 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c277
+ bl_0_277 br_0_277 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c277
+ bl_0_277 br_0_277 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c277
+ bl_0_277 br_0_277 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c277
+ bl_0_277 br_0_277 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c277
+ bl_0_277 br_0_277 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c277
+ bl_0_277 br_0_277 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c277
+ bl_0_277 br_0_277 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c277
+ bl_0_277 br_0_277 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c277
+ bl_0_277 br_0_277 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c277
+ bl_0_277 br_0_277 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c277
+ bl_0_277 br_0_277 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c277
+ bl_0_277 br_0_277 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c277
+ bl_0_277 br_0_277 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c277
+ bl_0_277 br_0_277 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c277
+ bl_0_277 br_0_277 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c277
+ bl_0_277 br_0_277 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c277
+ bl_0_277 br_0_277 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c277
+ bl_0_277 br_0_277 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c277
+ bl_0_277 br_0_277 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c277
+ bl_0_277 br_0_277 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c277
+ bl_0_277 br_0_277 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c277
+ bl_0_277 br_0_277 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c277
+ bl_0_277 br_0_277 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c277
+ bl_0_277 br_0_277 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c277
+ bl_0_277 br_0_277 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c277
+ bl_0_277 br_0_277 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c277
+ bl_0_277 br_0_277 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c277
+ bl_0_277 br_0_277 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c277
+ bl_0_277 br_0_277 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c277
+ bl_0_277 br_0_277 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c277
+ bl_0_277 br_0_277 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c277
+ bl_0_277 br_0_277 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c277
+ bl_0_277 br_0_277 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c277
+ bl_0_277 br_0_277 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c277
+ bl_0_277 br_0_277 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c277
+ bl_0_277 br_0_277 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c277
+ bl_0_277 br_0_277 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c277
+ bl_0_277 br_0_277 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c277
+ bl_0_277 br_0_277 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c277
+ bl_0_277 br_0_277 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c277
+ bl_0_277 br_0_277 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c277
+ bl_0_277 br_0_277 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c277
+ bl_0_277 br_0_277 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c277
+ bl_0_277 br_0_277 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c278
+ bl_0_278 br_0_278 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c278
+ bl_0_278 br_0_278 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c278
+ bl_0_278 br_0_278 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c278
+ bl_0_278 br_0_278 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c278
+ bl_0_278 br_0_278 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c278
+ bl_0_278 br_0_278 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c278
+ bl_0_278 br_0_278 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c278
+ bl_0_278 br_0_278 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c278
+ bl_0_278 br_0_278 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c278
+ bl_0_278 br_0_278 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c278
+ bl_0_278 br_0_278 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c278
+ bl_0_278 br_0_278 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c278
+ bl_0_278 br_0_278 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c278
+ bl_0_278 br_0_278 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c278
+ bl_0_278 br_0_278 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c278
+ bl_0_278 br_0_278 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c278
+ bl_0_278 br_0_278 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c278
+ bl_0_278 br_0_278 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c278
+ bl_0_278 br_0_278 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c278
+ bl_0_278 br_0_278 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c278
+ bl_0_278 br_0_278 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c278
+ bl_0_278 br_0_278 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c278
+ bl_0_278 br_0_278 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c278
+ bl_0_278 br_0_278 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c278
+ bl_0_278 br_0_278 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c278
+ bl_0_278 br_0_278 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c278
+ bl_0_278 br_0_278 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c278
+ bl_0_278 br_0_278 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c278
+ bl_0_278 br_0_278 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c278
+ bl_0_278 br_0_278 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c278
+ bl_0_278 br_0_278 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c278
+ bl_0_278 br_0_278 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c278
+ bl_0_278 br_0_278 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c278
+ bl_0_278 br_0_278 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c278
+ bl_0_278 br_0_278 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c278
+ bl_0_278 br_0_278 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c278
+ bl_0_278 br_0_278 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c278
+ bl_0_278 br_0_278 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c278
+ bl_0_278 br_0_278 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c278
+ bl_0_278 br_0_278 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c278
+ bl_0_278 br_0_278 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c278
+ bl_0_278 br_0_278 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c278
+ bl_0_278 br_0_278 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c278
+ bl_0_278 br_0_278 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c278
+ bl_0_278 br_0_278 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c279
+ bl_0_279 br_0_279 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c279
+ bl_0_279 br_0_279 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c279
+ bl_0_279 br_0_279 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c279
+ bl_0_279 br_0_279 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c279
+ bl_0_279 br_0_279 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c279
+ bl_0_279 br_0_279 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c279
+ bl_0_279 br_0_279 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c279
+ bl_0_279 br_0_279 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c279
+ bl_0_279 br_0_279 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c279
+ bl_0_279 br_0_279 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c279
+ bl_0_279 br_0_279 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c279
+ bl_0_279 br_0_279 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c279
+ bl_0_279 br_0_279 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c279
+ bl_0_279 br_0_279 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c279
+ bl_0_279 br_0_279 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c279
+ bl_0_279 br_0_279 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c279
+ bl_0_279 br_0_279 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c279
+ bl_0_279 br_0_279 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c279
+ bl_0_279 br_0_279 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c279
+ bl_0_279 br_0_279 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c279
+ bl_0_279 br_0_279 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c279
+ bl_0_279 br_0_279 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c279
+ bl_0_279 br_0_279 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c279
+ bl_0_279 br_0_279 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c279
+ bl_0_279 br_0_279 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c279
+ bl_0_279 br_0_279 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c279
+ bl_0_279 br_0_279 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c279
+ bl_0_279 br_0_279 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c279
+ bl_0_279 br_0_279 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c279
+ bl_0_279 br_0_279 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c279
+ bl_0_279 br_0_279 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c279
+ bl_0_279 br_0_279 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c279
+ bl_0_279 br_0_279 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c279
+ bl_0_279 br_0_279 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c279
+ bl_0_279 br_0_279 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c279
+ bl_0_279 br_0_279 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c279
+ bl_0_279 br_0_279 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c279
+ bl_0_279 br_0_279 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c279
+ bl_0_279 br_0_279 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c279
+ bl_0_279 br_0_279 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c279
+ bl_0_279 br_0_279 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c279
+ bl_0_279 br_0_279 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c279
+ bl_0_279 br_0_279 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c279
+ bl_0_279 br_0_279 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c279
+ bl_0_279 br_0_279 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c280
+ bl_0_280 br_0_280 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c280
+ bl_0_280 br_0_280 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c280
+ bl_0_280 br_0_280 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c280
+ bl_0_280 br_0_280 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c280
+ bl_0_280 br_0_280 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c280
+ bl_0_280 br_0_280 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c280
+ bl_0_280 br_0_280 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c280
+ bl_0_280 br_0_280 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c280
+ bl_0_280 br_0_280 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c280
+ bl_0_280 br_0_280 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c280
+ bl_0_280 br_0_280 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c280
+ bl_0_280 br_0_280 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c280
+ bl_0_280 br_0_280 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c280
+ bl_0_280 br_0_280 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c280
+ bl_0_280 br_0_280 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c280
+ bl_0_280 br_0_280 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c280
+ bl_0_280 br_0_280 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c280
+ bl_0_280 br_0_280 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c280
+ bl_0_280 br_0_280 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c280
+ bl_0_280 br_0_280 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c280
+ bl_0_280 br_0_280 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c280
+ bl_0_280 br_0_280 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c280
+ bl_0_280 br_0_280 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c280
+ bl_0_280 br_0_280 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c280
+ bl_0_280 br_0_280 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c280
+ bl_0_280 br_0_280 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c280
+ bl_0_280 br_0_280 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c280
+ bl_0_280 br_0_280 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c280
+ bl_0_280 br_0_280 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c280
+ bl_0_280 br_0_280 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c280
+ bl_0_280 br_0_280 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c280
+ bl_0_280 br_0_280 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c280
+ bl_0_280 br_0_280 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c280
+ bl_0_280 br_0_280 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c280
+ bl_0_280 br_0_280 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c280
+ bl_0_280 br_0_280 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c280
+ bl_0_280 br_0_280 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c280
+ bl_0_280 br_0_280 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c280
+ bl_0_280 br_0_280 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c280
+ bl_0_280 br_0_280 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c280
+ bl_0_280 br_0_280 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c280
+ bl_0_280 br_0_280 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c280
+ bl_0_280 br_0_280 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c280
+ bl_0_280 br_0_280 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c280
+ bl_0_280 br_0_280 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c281
+ bl_0_281 br_0_281 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c281
+ bl_0_281 br_0_281 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c281
+ bl_0_281 br_0_281 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c281
+ bl_0_281 br_0_281 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c281
+ bl_0_281 br_0_281 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c281
+ bl_0_281 br_0_281 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c281
+ bl_0_281 br_0_281 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c281
+ bl_0_281 br_0_281 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c281
+ bl_0_281 br_0_281 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c281
+ bl_0_281 br_0_281 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c281
+ bl_0_281 br_0_281 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c281
+ bl_0_281 br_0_281 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c281
+ bl_0_281 br_0_281 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c281
+ bl_0_281 br_0_281 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c281
+ bl_0_281 br_0_281 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c281
+ bl_0_281 br_0_281 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c281
+ bl_0_281 br_0_281 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c281
+ bl_0_281 br_0_281 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c281
+ bl_0_281 br_0_281 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c281
+ bl_0_281 br_0_281 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c281
+ bl_0_281 br_0_281 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c281
+ bl_0_281 br_0_281 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c281
+ bl_0_281 br_0_281 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c281
+ bl_0_281 br_0_281 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c281
+ bl_0_281 br_0_281 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c281
+ bl_0_281 br_0_281 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c281
+ bl_0_281 br_0_281 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c281
+ bl_0_281 br_0_281 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c281
+ bl_0_281 br_0_281 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c281
+ bl_0_281 br_0_281 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c281
+ bl_0_281 br_0_281 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c281
+ bl_0_281 br_0_281 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c281
+ bl_0_281 br_0_281 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c281
+ bl_0_281 br_0_281 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c281
+ bl_0_281 br_0_281 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c281
+ bl_0_281 br_0_281 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c281
+ bl_0_281 br_0_281 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c281
+ bl_0_281 br_0_281 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c281
+ bl_0_281 br_0_281 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c281
+ bl_0_281 br_0_281 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c281
+ bl_0_281 br_0_281 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c281
+ bl_0_281 br_0_281 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c281
+ bl_0_281 br_0_281 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c281
+ bl_0_281 br_0_281 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c281
+ bl_0_281 br_0_281 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c282
+ bl_0_282 br_0_282 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c282
+ bl_0_282 br_0_282 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c282
+ bl_0_282 br_0_282 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c282
+ bl_0_282 br_0_282 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c282
+ bl_0_282 br_0_282 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c282
+ bl_0_282 br_0_282 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c282
+ bl_0_282 br_0_282 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c282
+ bl_0_282 br_0_282 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c282
+ bl_0_282 br_0_282 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c282
+ bl_0_282 br_0_282 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c282
+ bl_0_282 br_0_282 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c282
+ bl_0_282 br_0_282 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c282
+ bl_0_282 br_0_282 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c282
+ bl_0_282 br_0_282 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c282
+ bl_0_282 br_0_282 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c282
+ bl_0_282 br_0_282 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c282
+ bl_0_282 br_0_282 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c282
+ bl_0_282 br_0_282 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c282
+ bl_0_282 br_0_282 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c282
+ bl_0_282 br_0_282 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c282
+ bl_0_282 br_0_282 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c282
+ bl_0_282 br_0_282 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c282
+ bl_0_282 br_0_282 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c282
+ bl_0_282 br_0_282 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c282
+ bl_0_282 br_0_282 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c282
+ bl_0_282 br_0_282 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c282
+ bl_0_282 br_0_282 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c282
+ bl_0_282 br_0_282 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c282
+ bl_0_282 br_0_282 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c282
+ bl_0_282 br_0_282 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c282
+ bl_0_282 br_0_282 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c282
+ bl_0_282 br_0_282 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c282
+ bl_0_282 br_0_282 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c282
+ bl_0_282 br_0_282 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c282
+ bl_0_282 br_0_282 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c282
+ bl_0_282 br_0_282 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c282
+ bl_0_282 br_0_282 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c282
+ bl_0_282 br_0_282 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c282
+ bl_0_282 br_0_282 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c282
+ bl_0_282 br_0_282 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c282
+ bl_0_282 br_0_282 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c282
+ bl_0_282 br_0_282 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c282
+ bl_0_282 br_0_282 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c282
+ bl_0_282 br_0_282 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c282
+ bl_0_282 br_0_282 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c283
+ bl_0_283 br_0_283 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c283
+ bl_0_283 br_0_283 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c283
+ bl_0_283 br_0_283 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c283
+ bl_0_283 br_0_283 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c283
+ bl_0_283 br_0_283 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c283
+ bl_0_283 br_0_283 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c283
+ bl_0_283 br_0_283 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c283
+ bl_0_283 br_0_283 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c283
+ bl_0_283 br_0_283 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c283
+ bl_0_283 br_0_283 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c283
+ bl_0_283 br_0_283 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c283
+ bl_0_283 br_0_283 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c283
+ bl_0_283 br_0_283 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c283
+ bl_0_283 br_0_283 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c283
+ bl_0_283 br_0_283 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c283
+ bl_0_283 br_0_283 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c283
+ bl_0_283 br_0_283 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c283
+ bl_0_283 br_0_283 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c283
+ bl_0_283 br_0_283 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c283
+ bl_0_283 br_0_283 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c283
+ bl_0_283 br_0_283 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c283
+ bl_0_283 br_0_283 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c283
+ bl_0_283 br_0_283 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c283
+ bl_0_283 br_0_283 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c283
+ bl_0_283 br_0_283 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c283
+ bl_0_283 br_0_283 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c283
+ bl_0_283 br_0_283 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c283
+ bl_0_283 br_0_283 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c283
+ bl_0_283 br_0_283 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c283
+ bl_0_283 br_0_283 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c283
+ bl_0_283 br_0_283 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c283
+ bl_0_283 br_0_283 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c283
+ bl_0_283 br_0_283 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c283
+ bl_0_283 br_0_283 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c283
+ bl_0_283 br_0_283 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c283
+ bl_0_283 br_0_283 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c283
+ bl_0_283 br_0_283 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c283
+ bl_0_283 br_0_283 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c283
+ bl_0_283 br_0_283 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c283
+ bl_0_283 br_0_283 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c283
+ bl_0_283 br_0_283 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c283
+ bl_0_283 br_0_283 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c283
+ bl_0_283 br_0_283 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c283
+ bl_0_283 br_0_283 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c283
+ bl_0_283 br_0_283 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c284
+ bl_0_284 br_0_284 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c284
+ bl_0_284 br_0_284 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c284
+ bl_0_284 br_0_284 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c284
+ bl_0_284 br_0_284 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c284
+ bl_0_284 br_0_284 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c284
+ bl_0_284 br_0_284 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c284
+ bl_0_284 br_0_284 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c284
+ bl_0_284 br_0_284 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c284
+ bl_0_284 br_0_284 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c284
+ bl_0_284 br_0_284 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c284
+ bl_0_284 br_0_284 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c284
+ bl_0_284 br_0_284 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c284
+ bl_0_284 br_0_284 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c284
+ bl_0_284 br_0_284 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c284
+ bl_0_284 br_0_284 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c284
+ bl_0_284 br_0_284 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c284
+ bl_0_284 br_0_284 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c284
+ bl_0_284 br_0_284 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c284
+ bl_0_284 br_0_284 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c284
+ bl_0_284 br_0_284 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c284
+ bl_0_284 br_0_284 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c284
+ bl_0_284 br_0_284 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c284
+ bl_0_284 br_0_284 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c284
+ bl_0_284 br_0_284 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c284
+ bl_0_284 br_0_284 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c284
+ bl_0_284 br_0_284 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c284
+ bl_0_284 br_0_284 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c284
+ bl_0_284 br_0_284 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c284
+ bl_0_284 br_0_284 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c284
+ bl_0_284 br_0_284 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c284
+ bl_0_284 br_0_284 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c284
+ bl_0_284 br_0_284 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c284
+ bl_0_284 br_0_284 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c284
+ bl_0_284 br_0_284 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c284
+ bl_0_284 br_0_284 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c284
+ bl_0_284 br_0_284 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c284
+ bl_0_284 br_0_284 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c284
+ bl_0_284 br_0_284 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c284
+ bl_0_284 br_0_284 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c284
+ bl_0_284 br_0_284 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c284
+ bl_0_284 br_0_284 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c284
+ bl_0_284 br_0_284 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c284
+ bl_0_284 br_0_284 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c284
+ bl_0_284 br_0_284 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c284
+ bl_0_284 br_0_284 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c285
+ bl_0_285 br_0_285 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c285
+ bl_0_285 br_0_285 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c285
+ bl_0_285 br_0_285 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c285
+ bl_0_285 br_0_285 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c285
+ bl_0_285 br_0_285 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c285
+ bl_0_285 br_0_285 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c285
+ bl_0_285 br_0_285 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c285
+ bl_0_285 br_0_285 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c285
+ bl_0_285 br_0_285 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c285
+ bl_0_285 br_0_285 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c285
+ bl_0_285 br_0_285 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c285
+ bl_0_285 br_0_285 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c285
+ bl_0_285 br_0_285 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c285
+ bl_0_285 br_0_285 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c285
+ bl_0_285 br_0_285 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c285
+ bl_0_285 br_0_285 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c285
+ bl_0_285 br_0_285 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c285
+ bl_0_285 br_0_285 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c285
+ bl_0_285 br_0_285 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c285
+ bl_0_285 br_0_285 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c285
+ bl_0_285 br_0_285 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c285
+ bl_0_285 br_0_285 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c285
+ bl_0_285 br_0_285 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c285
+ bl_0_285 br_0_285 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c285
+ bl_0_285 br_0_285 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c285
+ bl_0_285 br_0_285 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c285
+ bl_0_285 br_0_285 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c285
+ bl_0_285 br_0_285 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c285
+ bl_0_285 br_0_285 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c285
+ bl_0_285 br_0_285 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c285
+ bl_0_285 br_0_285 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c285
+ bl_0_285 br_0_285 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c285
+ bl_0_285 br_0_285 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c285
+ bl_0_285 br_0_285 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c285
+ bl_0_285 br_0_285 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c285
+ bl_0_285 br_0_285 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c285
+ bl_0_285 br_0_285 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c285
+ bl_0_285 br_0_285 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c285
+ bl_0_285 br_0_285 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c285
+ bl_0_285 br_0_285 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c285
+ bl_0_285 br_0_285 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c285
+ bl_0_285 br_0_285 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c285
+ bl_0_285 br_0_285 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c285
+ bl_0_285 br_0_285 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c285
+ bl_0_285 br_0_285 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c286
+ bl_0_286 br_0_286 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c286
+ bl_0_286 br_0_286 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c286
+ bl_0_286 br_0_286 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c286
+ bl_0_286 br_0_286 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c286
+ bl_0_286 br_0_286 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c286
+ bl_0_286 br_0_286 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c286
+ bl_0_286 br_0_286 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c286
+ bl_0_286 br_0_286 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c286
+ bl_0_286 br_0_286 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c286
+ bl_0_286 br_0_286 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c286
+ bl_0_286 br_0_286 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c286
+ bl_0_286 br_0_286 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c286
+ bl_0_286 br_0_286 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c286
+ bl_0_286 br_0_286 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c286
+ bl_0_286 br_0_286 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c286
+ bl_0_286 br_0_286 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c286
+ bl_0_286 br_0_286 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c286
+ bl_0_286 br_0_286 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c286
+ bl_0_286 br_0_286 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c286
+ bl_0_286 br_0_286 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c286
+ bl_0_286 br_0_286 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c286
+ bl_0_286 br_0_286 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c286
+ bl_0_286 br_0_286 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c286
+ bl_0_286 br_0_286 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c286
+ bl_0_286 br_0_286 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c286
+ bl_0_286 br_0_286 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c286
+ bl_0_286 br_0_286 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c286
+ bl_0_286 br_0_286 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c286
+ bl_0_286 br_0_286 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c286
+ bl_0_286 br_0_286 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c286
+ bl_0_286 br_0_286 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c286
+ bl_0_286 br_0_286 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c286
+ bl_0_286 br_0_286 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c286
+ bl_0_286 br_0_286 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c286
+ bl_0_286 br_0_286 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c286
+ bl_0_286 br_0_286 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c286
+ bl_0_286 br_0_286 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c286
+ bl_0_286 br_0_286 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c286
+ bl_0_286 br_0_286 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c286
+ bl_0_286 br_0_286 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c286
+ bl_0_286 br_0_286 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c286
+ bl_0_286 br_0_286 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c286
+ bl_0_286 br_0_286 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c286
+ bl_0_286 br_0_286 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c286
+ bl_0_286 br_0_286 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c287
+ bl_0_287 br_0_287 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c287
+ bl_0_287 br_0_287 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c287
+ bl_0_287 br_0_287 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c287
+ bl_0_287 br_0_287 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c287
+ bl_0_287 br_0_287 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c287
+ bl_0_287 br_0_287 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c287
+ bl_0_287 br_0_287 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c287
+ bl_0_287 br_0_287 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c287
+ bl_0_287 br_0_287 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c287
+ bl_0_287 br_0_287 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c287
+ bl_0_287 br_0_287 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c287
+ bl_0_287 br_0_287 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c287
+ bl_0_287 br_0_287 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c287
+ bl_0_287 br_0_287 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c287
+ bl_0_287 br_0_287 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c287
+ bl_0_287 br_0_287 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c287
+ bl_0_287 br_0_287 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c287
+ bl_0_287 br_0_287 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c287
+ bl_0_287 br_0_287 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c287
+ bl_0_287 br_0_287 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c287
+ bl_0_287 br_0_287 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c287
+ bl_0_287 br_0_287 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c287
+ bl_0_287 br_0_287 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c287
+ bl_0_287 br_0_287 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c287
+ bl_0_287 br_0_287 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c287
+ bl_0_287 br_0_287 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c287
+ bl_0_287 br_0_287 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c287
+ bl_0_287 br_0_287 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c287
+ bl_0_287 br_0_287 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c287
+ bl_0_287 br_0_287 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c287
+ bl_0_287 br_0_287 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c287
+ bl_0_287 br_0_287 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c287
+ bl_0_287 br_0_287 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c287
+ bl_0_287 br_0_287 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c287
+ bl_0_287 br_0_287 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c287
+ bl_0_287 br_0_287 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c287
+ bl_0_287 br_0_287 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c287
+ bl_0_287 br_0_287 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c287
+ bl_0_287 br_0_287 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c287
+ bl_0_287 br_0_287 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c287
+ bl_0_287 br_0_287 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c287
+ bl_0_287 br_0_287 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c287
+ bl_0_287 br_0_287 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c287
+ bl_0_287 br_0_287 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c287
+ bl_0_287 br_0_287 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c288
+ bl_0_288 br_0_288 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c288
+ bl_0_288 br_0_288 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c288
+ bl_0_288 br_0_288 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c288
+ bl_0_288 br_0_288 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c288
+ bl_0_288 br_0_288 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c288
+ bl_0_288 br_0_288 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c288
+ bl_0_288 br_0_288 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c288
+ bl_0_288 br_0_288 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c288
+ bl_0_288 br_0_288 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c288
+ bl_0_288 br_0_288 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c288
+ bl_0_288 br_0_288 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c288
+ bl_0_288 br_0_288 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c288
+ bl_0_288 br_0_288 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c288
+ bl_0_288 br_0_288 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c288
+ bl_0_288 br_0_288 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c288
+ bl_0_288 br_0_288 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c288
+ bl_0_288 br_0_288 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c288
+ bl_0_288 br_0_288 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c288
+ bl_0_288 br_0_288 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c288
+ bl_0_288 br_0_288 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c288
+ bl_0_288 br_0_288 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c288
+ bl_0_288 br_0_288 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c288
+ bl_0_288 br_0_288 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c288
+ bl_0_288 br_0_288 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c288
+ bl_0_288 br_0_288 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c288
+ bl_0_288 br_0_288 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c288
+ bl_0_288 br_0_288 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c288
+ bl_0_288 br_0_288 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c288
+ bl_0_288 br_0_288 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c288
+ bl_0_288 br_0_288 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c288
+ bl_0_288 br_0_288 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c288
+ bl_0_288 br_0_288 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c288
+ bl_0_288 br_0_288 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c288
+ bl_0_288 br_0_288 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c288
+ bl_0_288 br_0_288 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c288
+ bl_0_288 br_0_288 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c288
+ bl_0_288 br_0_288 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c288
+ bl_0_288 br_0_288 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c288
+ bl_0_288 br_0_288 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c288
+ bl_0_288 br_0_288 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c288
+ bl_0_288 br_0_288 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c288
+ bl_0_288 br_0_288 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c288
+ bl_0_288 br_0_288 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c288
+ bl_0_288 br_0_288 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c288
+ bl_0_288 br_0_288 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c289
+ bl_0_289 br_0_289 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c289
+ bl_0_289 br_0_289 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c289
+ bl_0_289 br_0_289 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c289
+ bl_0_289 br_0_289 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c289
+ bl_0_289 br_0_289 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c289
+ bl_0_289 br_0_289 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c289
+ bl_0_289 br_0_289 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c289
+ bl_0_289 br_0_289 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c289
+ bl_0_289 br_0_289 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c289
+ bl_0_289 br_0_289 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c289
+ bl_0_289 br_0_289 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c289
+ bl_0_289 br_0_289 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c289
+ bl_0_289 br_0_289 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c289
+ bl_0_289 br_0_289 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c289
+ bl_0_289 br_0_289 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c289
+ bl_0_289 br_0_289 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c289
+ bl_0_289 br_0_289 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c289
+ bl_0_289 br_0_289 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c289
+ bl_0_289 br_0_289 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c289
+ bl_0_289 br_0_289 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c289
+ bl_0_289 br_0_289 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c289
+ bl_0_289 br_0_289 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c289
+ bl_0_289 br_0_289 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c289
+ bl_0_289 br_0_289 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c289
+ bl_0_289 br_0_289 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c289
+ bl_0_289 br_0_289 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c289
+ bl_0_289 br_0_289 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c289
+ bl_0_289 br_0_289 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c289
+ bl_0_289 br_0_289 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c289
+ bl_0_289 br_0_289 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c289
+ bl_0_289 br_0_289 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c289
+ bl_0_289 br_0_289 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c289
+ bl_0_289 br_0_289 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c289
+ bl_0_289 br_0_289 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c289
+ bl_0_289 br_0_289 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c289
+ bl_0_289 br_0_289 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c289
+ bl_0_289 br_0_289 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c289
+ bl_0_289 br_0_289 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c289
+ bl_0_289 br_0_289 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c289
+ bl_0_289 br_0_289 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c289
+ bl_0_289 br_0_289 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c289
+ bl_0_289 br_0_289 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c289
+ bl_0_289 br_0_289 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c289
+ bl_0_289 br_0_289 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c289
+ bl_0_289 br_0_289 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c290
+ bl_0_290 br_0_290 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c290
+ bl_0_290 br_0_290 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c290
+ bl_0_290 br_0_290 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c290
+ bl_0_290 br_0_290 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c290
+ bl_0_290 br_0_290 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c290
+ bl_0_290 br_0_290 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c290
+ bl_0_290 br_0_290 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c290
+ bl_0_290 br_0_290 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c290
+ bl_0_290 br_0_290 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c290
+ bl_0_290 br_0_290 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c290
+ bl_0_290 br_0_290 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c290
+ bl_0_290 br_0_290 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c290
+ bl_0_290 br_0_290 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c290
+ bl_0_290 br_0_290 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c290
+ bl_0_290 br_0_290 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c290
+ bl_0_290 br_0_290 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c290
+ bl_0_290 br_0_290 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c290
+ bl_0_290 br_0_290 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c290
+ bl_0_290 br_0_290 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c290
+ bl_0_290 br_0_290 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c290
+ bl_0_290 br_0_290 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c290
+ bl_0_290 br_0_290 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c290
+ bl_0_290 br_0_290 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c290
+ bl_0_290 br_0_290 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c290
+ bl_0_290 br_0_290 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c290
+ bl_0_290 br_0_290 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c290
+ bl_0_290 br_0_290 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c290
+ bl_0_290 br_0_290 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c290
+ bl_0_290 br_0_290 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c290
+ bl_0_290 br_0_290 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c290
+ bl_0_290 br_0_290 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c290
+ bl_0_290 br_0_290 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c290
+ bl_0_290 br_0_290 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c290
+ bl_0_290 br_0_290 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c290
+ bl_0_290 br_0_290 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c290
+ bl_0_290 br_0_290 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c290
+ bl_0_290 br_0_290 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c290
+ bl_0_290 br_0_290 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c290
+ bl_0_290 br_0_290 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c290
+ bl_0_290 br_0_290 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c290
+ bl_0_290 br_0_290 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c290
+ bl_0_290 br_0_290 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c290
+ bl_0_290 br_0_290 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c290
+ bl_0_290 br_0_290 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c290
+ bl_0_290 br_0_290 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c291
+ bl_0_291 br_0_291 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c291
+ bl_0_291 br_0_291 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c291
+ bl_0_291 br_0_291 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c291
+ bl_0_291 br_0_291 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c291
+ bl_0_291 br_0_291 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c291
+ bl_0_291 br_0_291 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c291
+ bl_0_291 br_0_291 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c291
+ bl_0_291 br_0_291 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c291
+ bl_0_291 br_0_291 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c291
+ bl_0_291 br_0_291 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c291
+ bl_0_291 br_0_291 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c291
+ bl_0_291 br_0_291 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c291
+ bl_0_291 br_0_291 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c291
+ bl_0_291 br_0_291 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c291
+ bl_0_291 br_0_291 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c291
+ bl_0_291 br_0_291 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c291
+ bl_0_291 br_0_291 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c291
+ bl_0_291 br_0_291 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c291
+ bl_0_291 br_0_291 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c291
+ bl_0_291 br_0_291 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c291
+ bl_0_291 br_0_291 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c291
+ bl_0_291 br_0_291 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c291
+ bl_0_291 br_0_291 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c291
+ bl_0_291 br_0_291 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c291
+ bl_0_291 br_0_291 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c291
+ bl_0_291 br_0_291 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c291
+ bl_0_291 br_0_291 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c291
+ bl_0_291 br_0_291 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c291
+ bl_0_291 br_0_291 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c291
+ bl_0_291 br_0_291 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c291
+ bl_0_291 br_0_291 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c291
+ bl_0_291 br_0_291 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c291
+ bl_0_291 br_0_291 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c291
+ bl_0_291 br_0_291 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c291
+ bl_0_291 br_0_291 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c291
+ bl_0_291 br_0_291 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c291
+ bl_0_291 br_0_291 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c291
+ bl_0_291 br_0_291 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c291
+ bl_0_291 br_0_291 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c291
+ bl_0_291 br_0_291 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c291
+ bl_0_291 br_0_291 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c291
+ bl_0_291 br_0_291 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c291
+ bl_0_291 br_0_291 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c291
+ bl_0_291 br_0_291 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c291
+ bl_0_291 br_0_291 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c292
+ bl_0_292 br_0_292 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c292
+ bl_0_292 br_0_292 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c292
+ bl_0_292 br_0_292 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c292
+ bl_0_292 br_0_292 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c292
+ bl_0_292 br_0_292 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c292
+ bl_0_292 br_0_292 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c292
+ bl_0_292 br_0_292 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c292
+ bl_0_292 br_0_292 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c292
+ bl_0_292 br_0_292 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c292
+ bl_0_292 br_0_292 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c292
+ bl_0_292 br_0_292 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c292
+ bl_0_292 br_0_292 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c292
+ bl_0_292 br_0_292 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c292
+ bl_0_292 br_0_292 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c292
+ bl_0_292 br_0_292 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c292
+ bl_0_292 br_0_292 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c292
+ bl_0_292 br_0_292 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c292
+ bl_0_292 br_0_292 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c292
+ bl_0_292 br_0_292 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c292
+ bl_0_292 br_0_292 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c292
+ bl_0_292 br_0_292 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c292
+ bl_0_292 br_0_292 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c292
+ bl_0_292 br_0_292 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c292
+ bl_0_292 br_0_292 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c292
+ bl_0_292 br_0_292 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c292
+ bl_0_292 br_0_292 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c292
+ bl_0_292 br_0_292 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c292
+ bl_0_292 br_0_292 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c292
+ bl_0_292 br_0_292 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c292
+ bl_0_292 br_0_292 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c292
+ bl_0_292 br_0_292 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c292
+ bl_0_292 br_0_292 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c292
+ bl_0_292 br_0_292 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c292
+ bl_0_292 br_0_292 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c292
+ bl_0_292 br_0_292 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c292
+ bl_0_292 br_0_292 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c292
+ bl_0_292 br_0_292 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c292
+ bl_0_292 br_0_292 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c292
+ bl_0_292 br_0_292 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c292
+ bl_0_292 br_0_292 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c292
+ bl_0_292 br_0_292 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c292
+ bl_0_292 br_0_292 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c292
+ bl_0_292 br_0_292 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c292
+ bl_0_292 br_0_292 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c292
+ bl_0_292 br_0_292 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c293
+ bl_0_293 br_0_293 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c293
+ bl_0_293 br_0_293 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c293
+ bl_0_293 br_0_293 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c293
+ bl_0_293 br_0_293 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c293
+ bl_0_293 br_0_293 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c293
+ bl_0_293 br_0_293 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c293
+ bl_0_293 br_0_293 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c293
+ bl_0_293 br_0_293 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c293
+ bl_0_293 br_0_293 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c293
+ bl_0_293 br_0_293 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c293
+ bl_0_293 br_0_293 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c293
+ bl_0_293 br_0_293 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c293
+ bl_0_293 br_0_293 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c293
+ bl_0_293 br_0_293 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c293
+ bl_0_293 br_0_293 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c293
+ bl_0_293 br_0_293 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c293
+ bl_0_293 br_0_293 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c293
+ bl_0_293 br_0_293 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c293
+ bl_0_293 br_0_293 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c293
+ bl_0_293 br_0_293 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c293
+ bl_0_293 br_0_293 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c293
+ bl_0_293 br_0_293 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c293
+ bl_0_293 br_0_293 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c293
+ bl_0_293 br_0_293 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c293
+ bl_0_293 br_0_293 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c293
+ bl_0_293 br_0_293 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c293
+ bl_0_293 br_0_293 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c293
+ bl_0_293 br_0_293 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c293
+ bl_0_293 br_0_293 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c293
+ bl_0_293 br_0_293 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c293
+ bl_0_293 br_0_293 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c293
+ bl_0_293 br_0_293 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c293
+ bl_0_293 br_0_293 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c293
+ bl_0_293 br_0_293 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c293
+ bl_0_293 br_0_293 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c293
+ bl_0_293 br_0_293 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c293
+ bl_0_293 br_0_293 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c293
+ bl_0_293 br_0_293 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c293
+ bl_0_293 br_0_293 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c293
+ bl_0_293 br_0_293 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c293
+ bl_0_293 br_0_293 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c293
+ bl_0_293 br_0_293 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c293
+ bl_0_293 br_0_293 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c293
+ bl_0_293 br_0_293 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c293
+ bl_0_293 br_0_293 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c294
+ bl_0_294 br_0_294 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c294
+ bl_0_294 br_0_294 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c294
+ bl_0_294 br_0_294 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c294
+ bl_0_294 br_0_294 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c294
+ bl_0_294 br_0_294 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c294
+ bl_0_294 br_0_294 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c294
+ bl_0_294 br_0_294 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c294
+ bl_0_294 br_0_294 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c294
+ bl_0_294 br_0_294 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c294
+ bl_0_294 br_0_294 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c294
+ bl_0_294 br_0_294 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c294
+ bl_0_294 br_0_294 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c294
+ bl_0_294 br_0_294 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c294
+ bl_0_294 br_0_294 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c294
+ bl_0_294 br_0_294 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c294
+ bl_0_294 br_0_294 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c294
+ bl_0_294 br_0_294 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c294
+ bl_0_294 br_0_294 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c294
+ bl_0_294 br_0_294 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c294
+ bl_0_294 br_0_294 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c294
+ bl_0_294 br_0_294 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c294
+ bl_0_294 br_0_294 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c294
+ bl_0_294 br_0_294 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c294
+ bl_0_294 br_0_294 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c294
+ bl_0_294 br_0_294 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c294
+ bl_0_294 br_0_294 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c294
+ bl_0_294 br_0_294 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c294
+ bl_0_294 br_0_294 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c294
+ bl_0_294 br_0_294 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c294
+ bl_0_294 br_0_294 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c294
+ bl_0_294 br_0_294 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c294
+ bl_0_294 br_0_294 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c294
+ bl_0_294 br_0_294 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c294
+ bl_0_294 br_0_294 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c294
+ bl_0_294 br_0_294 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c294
+ bl_0_294 br_0_294 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c294
+ bl_0_294 br_0_294 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c294
+ bl_0_294 br_0_294 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c294
+ bl_0_294 br_0_294 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c294
+ bl_0_294 br_0_294 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c294
+ bl_0_294 br_0_294 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c294
+ bl_0_294 br_0_294 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c294
+ bl_0_294 br_0_294 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c294
+ bl_0_294 br_0_294 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c294
+ bl_0_294 br_0_294 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c295
+ bl_0_295 br_0_295 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c295
+ bl_0_295 br_0_295 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c295
+ bl_0_295 br_0_295 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c295
+ bl_0_295 br_0_295 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c295
+ bl_0_295 br_0_295 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c295
+ bl_0_295 br_0_295 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c295
+ bl_0_295 br_0_295 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c295
+ bl_0_295 br_0_295 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c295
+ bl_0_295 br_0_295 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c295
+ bl_0_295 br_0_295 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c295
+ bl_0_295 br_0_295 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c295
+ bl_0_295 br_0_295 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c295
+ bl_0_295 br_0_295 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c295
+ bl_0_295 br_0_295 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c295
+ bl_0_295 br_0_295 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c295
+ bl_0_295 br_0_295 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c295
+ bl_0_295 br_0_295 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c295
+ bl_0_295 br_0_295 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c295
+ bl_0_295 br_0_295 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c295
+ bl_0_295 br_0_295 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c295
+ bl_0_295 br_0_295 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c295
+ bl_0_295 br_0_295 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c295
+ bl_0_295 br_0_295 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c295
+ bl_0_295 br_0_295 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c295
+ bl_0_295 br_0_295 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c295
+ bl_0_295 br_0_295 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c295
+ bl_0_295 br_0_295 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c295
+ bl_0_295 br_0_295 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c295
+ bl_0_295 br_0_295 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c295
+ bl_0_295 br_0_295 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c295
+ bl_0_295 br_0_295 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c295
+ bl_0_295 br_0_295 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c295
+ bl_0_295 br_0_295 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c295
+ bl_0_295 br_0_295 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c295
+ bl_0_295 br_0_295 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c295
+ bl_0_295 br_0_295 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c295
+ bl_0_295 br_0_295 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c295
+ bl_0_295 br_0_295 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c295
+ bl_0_295 br_0_295 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c295
+ bl_0_295 br_0_295 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c295
+ bl_0_295 br_0_295 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c295
+ bl_0_295 br_0_295 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c295
+ bl_0_295 br_0_295 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c295
+ bl_0_295 br_0_295 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c295
+ bl_0_295 br_0_295 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c296
+ bl_0_296 br_0_296 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c296
+ bl_0_296 br_0_296 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c296
+ bl_0_296 br_0_296 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c296
+ bl_0_296 br_0_296 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c296
+ bl_0_296 br_0_296 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c296
+ bl_0_296 br_0_296 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c296
+ bl_0_296 br_0_296 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c296
+ bl_0_296 br_0_296 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c296
+ bl_0_296 br_0_296 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c296
+ bl_0_296 br_0_296 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c296
+ bl_0_296 br_0_296 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c296
+ bl_0_296 br_0_296 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c296
+ bl_0_296 br_0_296 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c296
+ bl_0_296 br_0_296 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c296
+ bl_0_296 br_0_296 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c296
+ bl_0_296 br_0_296 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c296
+ bl_0_296 br_0_296 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c296
+ bl_0_296 br_0_296 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c296
+ bl_0_296 br_0_296 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c296
+ bl_0_296 br_0_296 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c296
+ bl_0_296 br_0_296 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c296
+ bl_0_296 br_0_296 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c296
+ bl_0_296 br_0_296 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c296
+ bl_0_296 br_0_296 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c296
+ bl_0_296 br_0_296 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c296
+ bl_0_296 br_0_296 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c296
+ bl_0_296 br_0_296 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c296
+ bl_0_296 br_0_296 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c296
+ bl_0_296 br_0_296 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c296
+ bl_0_296 br_0_296 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c296
+ bl_0_296 br_0_296 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c296
+ bl_0_296 br_0_296 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c296
+ bl_0_296 br_0_296 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c296
+ bl_0_296 br_0_296 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c296
+ bl_0_296 br_0_296 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c296
+ bl_0_296 br_0_296 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c296
+ bl_0_296 br_0_296 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c296
+ bl_0_296 br_0_296 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c296
+ bl_0_296 br_0_296 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c296
+ bl_0_296 br_0_296 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c296
+ bl_0_296 br_0_296 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c296
+ bl_0_296 br_0_296 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c296
+ bl_0_296 br_0_296 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c296
+ bl_0_296 br_0_296 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c296
+ bl_0_296 br_0_296 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c297
+ bl_0_297 br_0_297 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c297
+ bl_0_297 br_0_297 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c297
+ bl_0_297 br_0_297 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c297
+ bl_0_297 br_0_297 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c297
+ bl_0_297 br_0_297 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c297
+ bl_0_297 br_0_297 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c297
+ bl_0_297 br_0_297 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c297
+ bl_0_297 br_0_297 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c297
+ bl_0_297 br_0_297 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c297
+ bl_0_297 br_0_297 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c297
+ bl_0_297 br_0_297 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c297
+ bl_0_297 br_0_297 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c297
+ bl_0_297 br_0_297 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c297
+ bl_0_297 br_0_297 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c297
+ bl_0_297 br_0_297 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c297
+ bl_0_297 br_0_297 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c297
+ bl_0_297 br_0_297 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c297
+ bl_0_297 br_0_297 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c297
+ bl_0_297 br_0_297 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c297
+ bl_0_297 br_0_297 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c297
+ bl_0_297 br_0_297 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c297
+ bl_0_297 br_0_297 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c297
+ bl_0_297 br_0_297 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c297
+ bl_0_297 br_0_297 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c297
+ bl_0_297 br_0_297 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c297
+ bl_0_297 br_0_297 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c297
+ bl_0_297 br_0_297 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c297
+ bl_0_297 br_0_297 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c297
+ bl_0_297 br_0_297 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c297
+ bl_0_297 br_0_297 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c297
+ bl_0_297 br_0_297 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c297
+ bl_0_297 br_0_297 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c297
+ bl_0_297 br_0_297 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c297
+ bl_0_297 br_0_297 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c297
+ bl_0_297 br_0_297 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c297
+ bl_0_297 br_0_297 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c297
+ bl_0_297 br_0_297 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c297
+ bl_0_297 br_0_297 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c297
+ bl_0_297 br_0_297 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c297
+ bl_0_297 br_0_297 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c297
+ bl_0_297 br_0_297 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c297
+ bl_0_297 br_0_297 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c297
+ bl_0_297 br_0_297 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c297
+ bl_0_297 br_0_297 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c297
+ bl_0_297 br_0_297 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c298
+ bl_0_298 br_0_298 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c298
+ bl_0_298 br_0_298 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c298
+ bl_0_298 br_0_298 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c298
+ bl_0_298 br_0_298 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c298
+ bl_0_298 br_0_298 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c298
+ bl_0_298 br_0_298 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c298
+ bl_0_298 br_0_298 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c298
+ bl_0_298 br_0_298 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c298
+ bl_0_298 br_0_298 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c298
+ bl_0_298 br_0_298 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c298
+ bl_0_298 br_0_298 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c298
+ bl_0_298 br_0_298 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c298
+ bl_0_298 br_0_298 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c298
+ bl_0_298 br_0_298 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c298
+ bl_0_298 br_0_298 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c298
+ bl_0_298 br_0_298 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c298
+ bl_0_298 br_0_298 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c298
+ bl_0_298 br_0_298 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c298
+ bl_0_298 br_0_298 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c298
+ bl_0_298 br_0_298 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c298
+ bl_0_298 br_0_298 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c298
+ bl_0_298 br_0_298 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c298
+ bl_0_298 br_0_298 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c298
+ bl_0_298 br_0_298 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c298
+ bl_0_298 br_0_298 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c298
+ bl_0_298 br_0_298 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c298
+ bl_0_298 br_0_298 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c298
+ bl_0_298 br_0_298 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c298
+ bl_0_298 br_0_298 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c298
+ bl_0_298 br_0_298 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c298
+ bl_0_298 br_0_298 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c298
+ bl_0_298 br_0_298 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c298
+ bl_0_298 br_0_298 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c298
+ bl_0_298 br_0_298 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c298
+ bl_0_298 br_0_298 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c298
+ bl_0_298 br_0_298 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c298
+ bl_0_298 br_0_298 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c298
+ bl_0_298 br_0_298 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c298
+ bl_0_298 br_0_298 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c298
+ bl_0_298 br_0_298 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c298
+ bl_0_298 br_0_298 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c298
+ bl_0_298 br_0_298 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c298
+ bl_0_298 br_0_298 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c298
+ bl_0_298 br_0_298 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c298
+ bl_0_298 br_0_298 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c299
+ bl_0_299 br_0_299 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c299
+ bl_0_299 br_0_299 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c299
+ bl_0_299 br_0_299 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c299
+ bl_0_299 br_0_299 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c299
+ bl_0_299 br_0_299 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c299
+ bl_0_299 br_0_299 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c299
+ bl_0_299 br_0_299 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c299
+ bl_0_299 br_0_299 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c299
+ bl_0_299 br_0_299 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c299
+ bl_0_299 br_0_299 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c299
+ bl_0_299 br_0_299 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c299
+ bl_0_299 br_0_299 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c299
+ bl_0_299 br_0_299 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c299
+ bl_0_299 br_0_299 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c299
+ bl_0_299 br_0_299 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c299
+ bl_0_299 br_0_299 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c299
+ bl_0_299 br_0_299 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c299
+ bl_0_299 br_0_299 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c299
+ bl_0_299 br_0_299 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c299
+ bl_0_299 br_0_299 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c299
+ bl_0_299 br_0_299 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c299
+ bl_0_299 br_0_299 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c299
+ bl_0_299 br_0_299 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c299
+ bl_0_299 br_0_299 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c299
+ bl_0_299 br_0_299 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c299
+ bl_0_299 br_0_299 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c299
+ bl_0_299 br_0_299 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c299
+ bl_0_299 br_0_299 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c299
+ bl_0_299 br_0_299 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c299
+ bl_0_299 br_0_299 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c299
+ bl_0_299 br_0_299 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c299
+ bl_0_299 br_0_299 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c299
+ bl_0_299 br_0_299 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c299
+ bl_0_299 br_0_299 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c299
+ bl_0_299 br_0_299 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c299
+ bl_0_299 br_0_299 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c299
+ bl_0_299 br_0_299 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c299
+ bl_0_299 br_0_299 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c299
+ bl_0_299 br_0_299 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c299
+ bl_0_299 br_0_299 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c299
+ bl_0_299 br_0_299 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c299
+ bl_0_299 br_0_299 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c299
+ bl_0_299 br_0_299 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c299
+ bl_0_299 br_0_299 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c299
+ bl_0_299 br_0_299 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c300
+ bl_0_300 br_0_300 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c300
+ bl_0_300 br_0_300 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c300
+ bl_0_300 br_0_300 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c300
+ bl_0_300 br_0_300 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c300
+ bl_0_300 br_0_300 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c300
+ bl_0_300 br_0_300 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c300
+ bl_0_300 br_0_300 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c300
+ bl_0_300 br_0_300 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c300
+ bl_0_300 br_0_300 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c300
+ bl_0_300 br_0_300 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c300
+ bl_0_300 br_0_300 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c300
+ bl_0_300 br_0_300 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c300
+ bl_0_300 br_0_300 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c300
+ bl_0_300 br_0_300 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c300
+ bl_0_300 br_0_300 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c300
+ bl_0_300 br_0_300 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c300
+ bl_0_300 br_0_300 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c300
+ bl_0_300 br_0_300 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c300
+ bl_0_300 br_0_300 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c300
+ bl_0_300 br_0_300 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c300
+ bl_0_300 br_0_300 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c300
+ bl_0_300 br_0_300 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c300
+ bl_0_300 br_0_300 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c300
+ bl_0_300 br_0_300 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c300
+ bl_0_300 br_0_300 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c300
+ bl_0_300 br_0_300 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c300
+ bl_0_300 br_0_300 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c300
+ bl_0_300 br_0_300 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c300
+ bl_0_300 br_0_300 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c300
+ bl_0_300 br_0_300 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c300
+ bl_0_300 br_0_300 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c300
+ bl_0_300 br_0_300 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c300
+ bl_0_300 br_0_300 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c300
+ bl_0_300 br_0_300 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c300
+ bl_0_300 br_0_300 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c300
+ bl_0_300 br_0_300 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c300
+ bl_0_300 br_0_300 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c300
+ bl_0_300 br_0_300 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c300
+ bl_0_300 br_0_300 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c300
+ bl_0_300 br_0_300 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c300
+ bl_0_300 br_0_300 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c300
+ bl_0_300 br_0_300 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c300
+ bl_0_300 br_0_300 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c300
+ bl_0_300 br_0_300 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c300
+ bl_0_300 br_0_300 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c301
+ bl_0_301 br_0_301 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c301
+ bl_0_301 br_0_301 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c301
+ bl_0_301 br_0_301 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c301
+ bl_0_301 br_0_301 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c301
+ bl_0_301 br_0_301 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c301
+ bl_0_301 br_0_301 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c301
+ bl_0_301 br_0_301 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c301
+ bl_0_301 br_0_301 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c301
+ bl_0_301 br_0_301 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c301
+ bl_0_301 br_0_301 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c301
+ bl_0_301 br_0_301 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c301
+ bl_0_301 br_0_301 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c301
+ bl_0_301 br_0_301 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c301
+ bl_0_301 br_0_301 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c301
+ bl_0_301 br_0_301 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c301
+ bl_0_301 br_0_301 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c301
+ bl_0_301 br_0_301 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c301
+ bl_0_301 br_0_301 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c301
+ bl_0_301 br_0_301 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c301
+ bl_0_301 br_0_301 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c301
+ bl_0_301 br_0_301 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c301
+ bl_0_301 br_0_301 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c301
+ bl_0_301 br_0_301 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c301
+ bl_0_301 br_0_301 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c301
+ bl_0_301 br_0_301 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c301
+ bl_0_301 br_0_301 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c301
+ bl_0_301 br_0_301 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c301
+ bl_0_301 br_0_301 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c301
+ bl_0_301 br_0_301 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c301
+ bl_0_301 br_0_301 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c301
+ bl_0_301 br_0_301 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c301
+ bl_0_301 br_0_301 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c301
+ bl_0_301 br_0_301 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c301
+ bl_0_301 br_0_301 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c301
+ bl_0_301 br_0_301 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c301
+ bl_0_301 br_0_301 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c301
+ bl_0_301 br_0_301 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c301
+ bl_0_301 br_0_301 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c301
+ bl_0_301 br_0_301 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c301
+ bl_0_301 br_0_301 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c301
+ bl_0_301 br_0_301 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c301
+ bl_0_301 br_0_301 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c301
+ bl_0_301 br_0_301 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c301
+ bl_0_301 br_0_301 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c301
+ bl_0_301 br_0_301 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c302
+ bl_0_302 br_0_302 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c302
+ bl_0_302 br_0_302 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c302
+ bl_0_302 br_0_302 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c302
+ bl_0_302 br_0_302 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c302
+ bl_0_302 br_0_302 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c302
+ bl_0_302 br_0_302 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c302
+ bl_0_302 br_0_302 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c302
+ bl_0_302 br_0_302 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c302
+ bl_0_302 br_0_302 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c302
+ bl_0_302 br_0_302 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c302
+ bl_0_302 br_0_302 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c302
+ bl_0_302 br_0_302 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c302
+ bl_0_302 br_0_302 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c302
+ bl_0_302 br_0_302 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c302
+ bl_0_302 br_0_302 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c302
+ bl_0_302 br_0_302 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c302
+ bl_0_302 br_0_302 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c302
+ bl_0_302 br_0_302 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c302
+ bl_0_302 br_0_302 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c302
+ bl_0_302 br_0_302 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c302
+ bl_0_302 br_0_302 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c302
+ bl_0_302 br_0_302 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c302
+ bl_0_302 br_0_302 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c302
+ bl_0_302 br_0_302 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c302
+ bl_0_302 br_0_302 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c302
+ bl_0_302 br_0_302 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c302
+ bl_0_302 br_0_302 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c302
+ bl_0_302 br_0_302 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c302
+ bl_0_302 br_0_302 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c302
+ bl_0_302 br_0_302 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c302
+ bl_0_302 br_0_302 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c302
+ bl_0_302 br_0_302 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c302
+ bl_0_302 br_0_302 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c302
+ bl_0_302 br_0_302 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c302
+ bl_0_302 br_0_302 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c302
+ bl_0_302 br_0_302 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c302
+ bl_0_302 br_0_302 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c302
+ bl_0_302 br_0_302 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c302
+ bl_0_302 br_0_302 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c302
+ bl_0_302 br_0_302 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c302
+ bl_0_302 br_0_302 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c302
+ bl_0_302 br_0_302 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c302
+ bl_0_302 br_0_302 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c302
+ bl_0_302 br_0_302 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c302
+ bl_0_302 br_0_302 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c303
+ bl_0_303 br_0_303 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c303
+ bl_0_303 br_0_303 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c303
+ bl_0_303 br_0_303 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c303
+ bl_0_303 br_0_303 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c303
+ bl_0_303 br_0_303 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c303
+ bl_0_303 br_0_303 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c303
+ bl_0_303 br_0_303 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c303
+ bl_0_303 br_0_303 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c303
+ bl_0_303 br_0_303 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c303
+ bl_0_303 br_0_303 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c303
+ bl_0_303 br_0_303 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c303
+ bl_0_303 br_0_303 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c303
+ bl_0_303 br_0_303 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c303
+ bl_0_303 br_0_303 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c303
+ bl_0_303 br_0_303 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c303
+ bl_0_303 br_0_303 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c303
+ bl_0_303 br_0_303 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c303
+ bl_0_303 br_0_303 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c303
+ bl_0_303 br_0_303 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c303
+ bl_0_303 br_0_303 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c303
+ bl_0_303 br_0_303 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c303
+ bl_0_303 br_0_303 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c303
+ bl_0_303 br_0_303 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c303
+ bl_0_303 br_0_303 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c303
+ bl_0_303 br_0_303 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c303
+ bl_0_303 br_0_303 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c303
+ bl_0_303 br_0_303 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c303
+ bl_0_303 br_0_303 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c303
+ bl_0_303 br_0_303 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c303
+ bl_0_303 br_0_303 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c303
+ bl_0_303 br_0_303 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c303
+ bl_0_303 br_0_303 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c303
+ bl_0_303 br_0_303 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c303
+ bl_0_303 br_0_303 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c303
+ bl_0_303 br_0_303 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c303
+ bl_0_303 br_0_303 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c303
+ bl_0_303 br_0_303 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c303
+ bl_0_303 br_0_303 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c303
+ bl_0_303 br_0_303 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c303
+ bl_0_303 br_0_303 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c303
+ bl_0_303 br_0_303 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c303
+ bl_0_303 br_0_303 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c303
+ bl_0_303 br_0_303 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c303
+ bl_0_303 br_0_303 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c303
+ bl_0_303 br_0_303 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c304
+ bl_0_304 br_0_304 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c304
+ bl_0_304 br_0_304 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c304
+ bl_0_304 br_0_304 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c304
+ bl_0_304 br_0_304 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c304
+ bl_0_304 br_0_304 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c304
+ bl_0_304 br_0_304 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c304
+ bl_0_304 br_0_304 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c304
+ bl_0_304 br_0_304 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c304
+ bl_0_304 br_0_304 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c304
+ bl_0_304 br_0_304 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c304
+ bl_0_304 br_0_304 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c304
+ bl_0_304 br_0_304 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c304
+ bl_0_304 br_0_304 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c304
+ bl_0_304 br_0_304 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c304
+ bl_0_304 br_0_304 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c304
+ bl_0_304 br_0_304 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c304
+ bl_0_304 br_0_304 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c304
+ bl_0_304 br_0_304 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c304
+ bl_0_304 br_0_304 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c304
+ bl_0_304 br_0_304 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c304
+ bl_0_304 br_0_304 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c304
+ bl_0_304 br_0_304 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c304
+ bl_0_304 br_0_304 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c304
+ bl_0_304 br_0_304 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c304
+ bl_0_304 br_0_304 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c304
+ bl_0_304 br_0_304 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c304
+ bl_0_304 br_0_304 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c304
+ bl_0_304 br_0_304 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c304
+ bl_0_304 br_0_304 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c304
+ bl_0_304 br_0_304 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c304
+ bl_0_304 br_0_304 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c304
+ bl_0_304 br_0_304 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c304
+ bl_0_304 br_0_304 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c304
+ bl_0_304 br_0_304 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c304
+ bl_0_304 br_0_304 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c304
+ bl_0_304 br_0_304 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c304
+ bl_0_304 br_0_304 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c304
+ bl_0_304 br_0_304 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c304
+ bl_0_304 br_0_304 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c304
+ bl_0_304 br_0_304 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c304
+ bl_0_304 br_0_304 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c304
+ bl_0_304 br_0_304 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c304
+ bl_0_304 br_0_304 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c304
+ bl_0_304 br_0_304 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c304
+ bl_0_304 br_0_304 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c305
+ bl_0_305 br_0_305 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c305
+ bl_0_305 br_0_305 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c305
+ bl_0_305 br_0_305 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c305
+ bl_0_305 br_0_305 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c305
+ bl_0_305 br_0_305 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c305
+ bl_0_305 br_0_305 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c305
+ bl_0_305 br_0_305 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c305
+ bl_0_305 br_0_305 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c305
+ bl_0_305 br_0_305 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c305
+ bl_0_305 br_0_305 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c305
+ bl_0_305 br_0_305 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c305
+ bl_0_305 br_0_305 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c305
+ bl_0_305 br_0_305 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c305
+ bl_0_305 br_0_305 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c305
+ bl_0_305 br_0_305 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c305
+ bl_0_305 br_0_305 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c305
+ bl_0_305 br_0_305 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c305
+ bl_0_305 br_0_305 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c305
+ bl_0_305 br_0_305 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c305
+ bl_0_305 br_0_305 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c305
+ bl_0_305 br_0_305 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c305
+ bl_0_305 br_0_305 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c305
+ bl_0_305 br_0_305 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c305
+ bl_0_305 br_0_305 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c305
+ bl_0_305 br_0_305 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c305
+ bl_0_305 br_0_305 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c305
+ bl_0_305 br_0_305 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c305
+ bl_0_305 br_0_305 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c305
+ bl_0_305 br_0_305 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c305
+ bl_0_305 br_0_305 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c305
+ bl_0_305 br_0_305 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c305
+ bl_0_305 br_0_305 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c305
+ bl_0_305 br_0_305 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c305
+ bl_0_305 br_0_305 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c305
+ bl_0_305 br_0_305 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c305
+ bl_0_305 br_0_305 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c305
+ bl_0_305 br_0_305 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c305
+ bl_0_305 br_0_305 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c305
+ bl_0_305 br_0_305 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c305
+ bl_0_305 br_0_305 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c305
+ bl_0_305 br_0_305 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c305
+ bl_0_305 br_0_305 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c305
+ bl_0_305 br_0_305 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c305
+ bl_0_305 br_0_305 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c305
+ bl_0_305 br_0_305 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c306
+ bl_0_306 br_0_306 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c306
+ bl_0_306 br_0_306 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c306
+ bl_0_306 br_0_306 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c306
+ bl_0_306 br_0_306 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c306
+ bl_0_306 br_0_306 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c306
+ bl_0_306 br_0_306 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c306
+ bl_0_306 br_0_306 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c306
+ bl_0_306 br_0_306 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c306
+ bl_0_306 br_0_306 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c306
+ bl_0_306 br_0_306 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c306
+ bl_0_306 br_0_306 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c306
+ bl_0_306 br_0_306 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c306
+ bl_0_306 br_0_306 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c306
+ bl_0_306 br_0_306 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c306
+ bl_0_306 br_0_306 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c306
+ bl_0_306 br_0_306 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c306
+ bl_0_306 br_0_306 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c306
+ bl_0_306 br_0_306 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c306
+ bl_0_306 br_0_306 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c306
+ bl_0_306 br_0_306 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c306
+ bl_0_306 br_0_306 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c306
+ bl_0_306 br_0_306 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c306
+ bl_0_306 br_0_306 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c306
+ bl_0_306 br_0_306 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c306
+ bl_0_306 br_0_306 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c306
+ bl_0_306 br_0_306 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c306
+ bl_0_306 br_0_306 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c306
+ bl_0_306 br_0_306 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c306
+ bl_0_306 br_0_306 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c306
+ bl_0_306 br_0_306 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c306
+ bl_0_306 br_0_306 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c306
+ bl_0_306 br_0_306 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c306
+ bl_0_306 br_0_306 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c306
+ bl_0_306 br_0_306 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c306
+ bl_0_306 br_0_306 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c306
+ bl_0_306 br_0_306 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c306
+ bl_0_306 br_0_306 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c306
+ bl_0_306 br_0_306 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c306
+ bl_0_306 br_0_306 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c306
+ bl_0_306 br_0_306 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c306
+ bl_0_306 br_0_306 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c306
+ bl_0_306 br_0_306 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c306
+ bl_0_306 br_0_306 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c306
+ bl_0_306 br_0_306 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c306
+ bl_0_306 br_0_306 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c307
+ bl_0_307 br_0_307 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c307
+ bl_0_307 br_0_307 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c307
+ bl_0_307 br_0_307 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c307
+ bl_0_307 br_0_307 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c307
+ bl_0_307 br_0_307 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c307
+ bl_0_307 br_0_307 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c307
+ bl_0_307 br_0_307 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c307
+ bl_0_307 br_0_307 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c307
+ bl_0_307 br_0_307 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c307
+ bl_0_307 br_0_307 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c307
+ bl_0_307 br_0_307 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c307
+ bl_0_307 br_0_307 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c307
+ bl_0_307 br_0_307 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c307
+ bl_0_307 br_0_307 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c307
+ bl_0_307 br_0_307 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c307
+ bl_0_307 br_0_307 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c307
+ bl_0_307 br_0_307 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c307
+ bl_0_307 br_0_307 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c307
+ bl_0_307 br_0_307 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c307
+ bl_0_307 br_0_307 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c307
+ bl_0_307 br_0_307 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c307
+ bl_0_307 br_0_307 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c307
+ bl_0_307 br_0_307 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c307
+ bl_0_307 br_0_307 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c307
+ bl_0_307 br_0_307 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c307
+ bl_0_307 br_0_307 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c307
+ bl_0_307 br_0_307 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c307
+ bl_0_307 br_0_307 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c307
+ bl_0_307 br_0_307 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c307
+ bl_0_307 br_0_307 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c307
+ bl_0_307 br_0_307 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c307
+ bl_0_307 br_0_307 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c307
+ bl_0_307 br_0_307 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c307
+ bl_0_307 br_0_307 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c307
+ bl_0_307 br_0_307 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c307
+ bl_0_307 br_0_307 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c307
+ bl_0_307 br_0_307 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c307
+ bl_0_307 br_0_307 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c307
+ bl_0_307 br_0_307 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c307
+ bl_0_307 br_0_307 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c307
+ bl_0_307 br_0_307 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c307
+ bl_0_307 br_0_307 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c307
+ bl_0_307 br_0_307 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c307
+ bl_0_307 br_0_307 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c307
+ bl_0_307 br_0_307 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c308
+ bl_0_308 br_0_308 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c308
+ bl_0_308 br_0_308 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c308
+ bl_0_308 br_0_308 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c308
+ bl_0_308 br_0_308 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c308
+ bl_0_308 br_0_308 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c308
+ bl_0_308 br_0_308 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c308
+ bl_0_308 br_0_308 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c308
+ bl_0_308 br_0_308 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c308
+ bl_0_308 br_0_308 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c308
+ bl_0_308 br_0_308 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c308
+ bl_0_308 br_0_308 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c308
+ bl_0_308 br_0_308 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c308
+ bl_0_308 br_0_308 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c308
+ bl_0_308 br_0_308 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c308
+ bl_0_308 br_0_308 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c308
+ bl_0_308 br_0_308 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c308
+ bl_0_308 br_0_308 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c308
+ bl_0_308 br_0_308 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c308
+ bl_0_308 br_0_308 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c308
+ bl_0_308 br_0_308 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c308
+ bl_0_308 br_0_308 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c308
+ bl_0_308 br_0_308 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c308
+ bl_0_308 br_0_308 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c308
+ bl_0_308 br_0_308 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c308
+ bl_0_308 br_0_308 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c308
+ bl_0_308 br_0_308 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c308
+ bl_0_308 br_0_308 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c308
+ bl_0_308 br_0_308 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c308
+ bl_0_308 br_0_308 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c308
+ bl_0_308 br_0_308 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c308
+ bl_0_308 br_0_308 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c308
+ bl_0_308 br_0_308 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c308
+ bl_0_308 br_0_308 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c308
+ bl_0_308 br_0_308 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c308
+ bl_0_308 br_0_308 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c308
+ bl_0_308 br_0_308 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c308
+ bl_0_308 br_0_308 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c308
+ bl_0_308 br_0_308 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c308
+ bl_0_308 br_0_308 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c308
+ bl_0_308 br_0_308 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c308
+ bl_0_308 br_0_308 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c308
+ bl_0_308 br_0_308 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c308
+ bl_0_308 br_0_308 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c308
+ bl_0_308 br_0_308 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c308
+ bl_0_308 br_0_308 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c309
+ bl_0_309 br_0_309 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c309
+ bl_0_309 br_0_309 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c309
+ bl_0_309 br_0_309 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c309
+ bl_0_309 br_0_309 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c309
+ bl_0_309 br_0_309 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c309
+ bl_0_309 br_0_309 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c309
+ bl_0_309 br_0_309 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c309
+ bl_0_309 br_0_309 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c309
+ bl_0_309 br_0_309 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c309
+ bl_0_309 br_0_309 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c309
+ bl_0_309 br_0_309 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c309
+ bl_0_309 br_0_309 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c309
+ bl_0_309 br_0_309 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c309
+ bl_0_309 br_0_309 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c309
+ bl_0_309 br_0_309 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c309
+ bl_0_309 br_0_309 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c309
+ bl_0_309 br_0_309 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c309
+ bl_0_309 br_0_309 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c309
+ bl_0_309 br_0_309 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c309
+ bl_0_309 br_0_309 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c309
+ bl_0_309 br_0_309 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c309
+ bl_0_309 br_0_309 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c309
+ bl_0_309 br_0_309 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c309
+ bl_0_309 br_0_309 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c309
+ bl_0_309 br_0_309 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c309
+ bl_0_309 br_0_309 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c309
+ bl_0_309 br_0_309 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c309
+ bl_0_309 br_0_309 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c309
+ bl_0_309 br_0_309 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c309
+ bl_0_309 br_0_309 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c309
+ bl_0_309 br_0_309 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c309
+ bl_0_309 br_0_309 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c309
+ bl_0_309 br_0_309 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c309
+ bl_0_309 br_0_309 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c309
+ bl_0_309 br_0_309 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c309
+ bl_0_309 br_0_309 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c309
+ bl_0_309 br_0_309 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c309
+ bl_0_309 br_0_309 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c309
+ bl_0_309 br_0_309 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c309
+ bl_0_309 br_0_309 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c309
+ bl_0_309 br_0_309 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c309
+ bl_0_309 br_0_309 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c309
+ bl_0_309 br_0_309 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c309
+ bl_0_309 br_0_309 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c309
+ bl_0_309 br_0_309 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c310
+ bl_0_310 br_0_310 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c310
+ bl_0_310 br_0_310 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c310
+ bl_0_310 br_0_310 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c310
+ bl_0_310 br_0_310 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c310
+ bl_0_310 br_0_310 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c310
+ bl_0_310 br_0_310 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c310
+ bl_0_310 br_0_310 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c310
+ bl_0_310 br_0_310 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c310
+ bl_0_310 br_0_310 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c310
+ bl_0_310 br_0_310 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c310
+ bl_0_310 br_0_310 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c310
+ bl_0_310 br_0_310 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c310
+ bl_0_310 br_0_310 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c310
+ bl_0_310 br_0_310 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c310
+ bl_0_310 br_0_310 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c310
+ bl_0_310 br_0_310 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c310
+ bl_0_310 br_0_310 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c310
+ bl_0_310 br_0_310 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c310
+ bl_0_310 br_0_310 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c310
+ bl_0_310 br_0_310 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c310
+ bl_0_310 br_0_310 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c310
+ bl_0_310 br_0_310 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c310
+ bl_0_310 br_0_310 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c310
+ bl_0_310 br_0_310 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c310
+ bl_0_310 br_0_310 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c310
+ bl_0_310 br_0_310 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c310
+ bl_0_310 br_0_310 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c310
+ bl_0_310 br_0_310 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c310
+ bl_0_310 br_0_310 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c310
+ bl_0_310 br_0_310 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c310
+ bl_0_310 br_0_310 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c310
+ bl_0_310 br_0_310 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c310
+ bl_0_310 br_0_310 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c310
+ bl_0_310 br_0_310 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c310
+ bl_0_310 br_0_310 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c310
+ bl_0_310 br_0_310 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c310
+ bl_0_310 br_0_310 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c310
+ bl_0_310 br_0_310 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c310
+ bl_0_310 br_0_310 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c310
+ bl_0_310 br_0_310 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c310
+ bl_0_310 br_0_310 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c310
+ bl_0_310 br_0_310 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c310
+ bl_0_310 br_0_310 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c310
+ bl_0_310 br_0_310 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c310
+ bl_0_310 br_0_310 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c311
+ bl_0_311 br_0_311 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c311
+ bl_0_311 br_0_311 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c311
+ bl_0_311 br_0_311 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c311
+ bl_0_311 br_0_311 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c311
+ bl_0_311 br_0_311 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c311
+ bl_0_311 br_0_311 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c311
+ bl_0_311 br_0_311 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c311
+ bl_0_311 br_0_311 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c311
+ bl_0_311 br_0_311 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c311
+ bl_0_311 br_0_311 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c311
+ bl_0_311 br_0_311 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c311
+ bl_0_311 br_0_311 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c311
+ bl_0_311 br_0_311 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c311
+ bl_0_311 br_0_311 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c311
+ bl_0_311 br_0_311 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c311
+ bl_0_311 br_0_311 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c311
+ bl_0_311 br_0_311 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c311
+ bl_0_311 br_0_311 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c311
+ bl_0_311 br_0_311 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c311
+ bl_0_311 br_0_311 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c311
+ bl_0_311 br_0_311 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c311
+ bl_0_311 br_0_311 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c311
+ bl_0_311 br_0_311 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c311
+ bl_0_311 br_0_311 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c311
+ bl_0_311 br_0_311 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c311
+ bl_0_311 br_0_311 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c311
+ bl_0_311 br_0_311 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c311
+ bl_0_311 br_0_311 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c311
+ bl_0_311 br_0_311 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c311
+ bl_0_311 br_0_311 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c311
+ bl_0_311 br_0_311 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c311
+ bl_0_311 br_0_311 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c311
+ bl_0_311 br_0_311 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c311
+ bl_0_311 br_0_311 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c311
+ bl_0_311 br_0_311 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c311
+ bl_0_311 br_0_311 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c311
+ bl_0_311 br_0_311 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c311
+ bl_0_311 br_0_311 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c311
+ bl_0_311 br_0_311 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c311
+ bl_0_311 br_0_311 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c311
+ bl_0_311 br_0_311 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c311
+ bl_0_311 br_0_311 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c311
+ bl_0_311 br_0_311 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c311
+ bl_0_311 br_0_311 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c311
+ bl_0_311 br_0_311 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c312
+ bl_0_312 br_0_312 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c312
+ bl_0_312 br_0_312 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c312
+ bl_0_312 br_0_312 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c312
+ bl_0_312 br_0_312 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c312
+ bl_0_312 br_0_312 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c312
+ bl_0_312 br_0_312 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c312
+ bl_0_312 br_0_312 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c312
+ bl_0_312 br_0_312 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c312
+ bl_0_312 br_0_312 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c312
+ bl_0_312 br_0_312 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c312
+ bl_0_312 br_0_312 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c312
+ bl_0_312 br_0_312 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c312
+ bl_0_312 br_0_312 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c312
+ bl_0_312 br_0_312 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c312
+ bl_0_312 br_0_312 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c312
+ bl_0_312 br_0_312 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c312
+ bl_0_312 br_0_312 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c312
+ bl_0_312 br_0_312 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c312
+ bl_0_312 br_0_312 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c312
+ bl_0_312 br_0_312 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c312
+ bl_0_312 br_0_312 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c312
+ bl_0_312 br_0_312 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c312
+ bl_0_312 br_0_312 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c312
+ bl_0_312 br_0_312 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c312
+ bl_0_312 br_0_312 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c312
+ bl_0_312 br_0_312 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c312
+ bl_0_312 br_0_312 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c312
+ bl_0_312 br_0_312 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c312
+ bl_0_312 br_0_312 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c312
+ bl_0_312 br_0_312 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c312
+ bl_0_312 br_0_312 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c312
+ bl_0_312 br_0_312 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c312
+ bl_0_312 br_0_312 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c312
+ bl_0_312 br_0_312 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c312
+ bl_0_312 br_0_312 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c312
+ bl_0_312 br_0_312 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c312
+ bl_0_312 br_0_312 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c312
+ bl_0_312 br_0_312 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c312
+ bl_0_312 br_0_312 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c312
+ bl_0_312 br_0_312 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c312
+ bl_0_312 br_0_312 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c312
+ bl_0_312 br_0_312 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c312
+ bl_0_312 br_0_312 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c312
+ bl_0_312 br_0_312 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c312
+ bl_0_312 br_0_312 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c313
+ bl_0_313 br_0_313 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c313
+ bl_0_313 br_0_313 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c313
+ bl_0_313 br_0_313 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c313
+ bl_0_313 br_0_313 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c313
+ bl_0_313 br_0_313 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c313
+ bl_0_313 br_0_313 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c313
+ bl_0_313 br_0_313 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c313
+ bl_0_313 br_0_313 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c313
+ bl_0_313 br_0_313 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c313
+ bl_0_313 br_0_313 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c313
+ bl_0_313 br_0_313 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c313
+ bl_0_313 br_0_313 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c313
+ bl_0_313 br_0_313 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c313
+ bl_0_313 br_0_313 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c313
+ bl_0_313 br_0_313 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c313
+ bl_0_313 br_0_313 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c313
+ bl_0_313 br_0_313 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c313
+ bl_0_313 br_0_313 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c313
+ bl_0_313 br_0_313 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c313
+ bl_0_313 br_0_313 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c313
+ bl_0_313 br_0_313 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c313
+ bl_0_313 br_0_313 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c313
+ bl_0_313 br_0_313 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c313
+ bl_0_313 br_0_313 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c313
+ bl_0_313 br_0_313 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c313
+ bl_0_313 br_0_313 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c313
+ bl_0_313 br_0_313 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c313
+ bl_0_313 br_0_313 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c313
+ bl_0_313 br_0_313 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c313
+ bl_0_313 br_0_313 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c313
+ bl_0_313 br_0_313 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c313
+ bl_0_313 br_0_313 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c313
+ bl_0_313 br_0_313 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c313
+ bl_0_313 br_0_313 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c313
+ bl_0_313 br_0_313 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c313
+ bl_0_313 br_0_313 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c313
+ bl_0_313 br_0_313 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c313
+ bl_0_313 br_0_313 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c313
+ bl_0_313 br_0_313 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c313
+ bl_0_313 br_0_313 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c313
+ bl_0_313 br_0_313 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c313
+ bl_0_313 br_0_313 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c313
+ bl_0_313 br_0_313 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c313
+ bl_0_313 br_0_313 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c313
+ bl_0_313 br_0_313 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c314
+ bl_0_314 br_0_314 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c314
+ bl_0_314 br_0_314 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c314
+ bl_0_314 br_0_314 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c314
+ bl_0_314 br_0_314 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c314
+ bl_0_314 br_0_314 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c314
+ bl_0_314 br_0_314 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c314
+ bl_0_314 br_0_314 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c314
+ bl_0_314 br_0_314 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c314
+ bl_0_314 br_0_314 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c314
+ bl_0_314 br_0_314 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c314
+ bl_0_314 br_0_314 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c314
+ bl_0_314 br_0_314 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c314
+ bl_0_314 br_0_314 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c314
+ bl_0_314 br_0_314 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c314
+ bl_0_314 br_0_314 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c314
+ bl_0_314 br_0_314 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c314
+ bl_0_314 br_0_314 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c314
+ bl_0_314 br_0_314 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c314
+ bl_0_314 br_0_314 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c314
+ bl_0_314 br_0_314 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c314
+ bl_0_314 br_0_314 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c314
+ bl_0_314 br_0_314 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c314
+ bl_0_314 br_0_314 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c314
+ bl_0_314 br_0_314 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c314
+ bl_0_314 br_0_314 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c314
+ bl_0_314 br_0_314 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c314
+ bl_0_314 br_0_314 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c314
+ bl_0_314 br_0_314 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c314
+ bl_0_314 br_0_314 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c314
+ bl_0_314 br_0_314 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c314
+ bl_0_314 br_0_314 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c314
+ bl_0_314 br_0_314 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c314
+ bl_0_314 br_0_314 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c314
+ bl_0_314 br_0_314 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c314
+ bl_0_314 br_0_314 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c314
+ bl_0_314 br_0_314 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c314
+ bl_0_314 br_0_314 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c314
+ bl_0_314 br_0_314 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c314
+ bl_0_314 br_0_314 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c314
+ bl_0_314 br_0_314 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c314
+ bl_0_314 br_0_314 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c314
+ bl_0_314 br_0_314 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c314
+ bl_0_314 br_0_314 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c314
+ bl_0_314 br_0_314 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c314
+ bl_0_314 br_0_314 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c315
+ bl_0_315 br_0_315 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c315
+ bl_0_315 br_0_315 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c315
+ bl_0_315 br_0_315 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c315
+ bl_0_315 br_0_315 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c315
+ bl_0_315 br_0_315 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c315
+ bl_0_315 br_0_315 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c315
+ bl_0_315 br_0_315 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c315
+ bl_0_315 br_0_315 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c315
+ bl_0_315 br_0_315 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c315
+ bl_0_315 br_0_315 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c315
+ bl_0_315 br_0_315 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c315
+ bl_0_315 br_0_315 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c315
+ bl_0_315 br_0_315 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c315
+ bl_0_315 br_0_315 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c315
+ bl_0_315 br_0_315 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c315
+ bl_0_315 br_0_315 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c315
+ bl_0_315 br_0_315 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c315
+ bl_0_315 br_0_315 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c315
+ bl_0_315 br_0_315 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c315
+ bl_0_315 br_0_315 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c315
+ bl_0_315 br_0_315 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c315
+ bl_0_315 br_0_315 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c315
+ bl_0_315 br_0_315 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c315
+ bl_0_315 br_0_315 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c315
+ bl_0_315 br_0_315 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c315
+ bl_0_315 br_0_315 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c315
+ bl_0_315 br_0_315 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c315
+ bl_0_315 br_0_315 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c315
+ bl_0_315 br_0_315 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c315
+ bl_0_315 br_0_315 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c315
+ bl_0_315 br_0_315 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c315
+ bl_0_315 br_0_315 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c315
+ bl_0_315 br_0_315 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c315
+ bl_0_315 br_0_315 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c315
+ bl_0_315 br_0_315 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c315
+ bl_0_315 br_0_315 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c315
+ bl_0_315 br_0_315 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c315
+ bl_0_315 br_0_315 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c315
+ bl_0_315 br_0_315 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c315
+ bl_0_315 br_0_315 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c315
+ bl_0_315 br_0_315 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c315
+ bl_0_315 br_0_315 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c315
+ bl_0_315 br_0_315 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c315
+ bl_0_315 br_0_315 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c315
+ bl_0_315 br_0_315 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c316
+ bl_0_316 br_0_316 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c316
+ bl_0_316 br_0_316 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c316
+ bl_0_316 br_0_316 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c316
+ bl_0_316 br_0_316 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c316
+ bl_0_316 br_0_316 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c316
+ bl_0_316 br_0_316 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c316
+ bl_0_316 br_0_316 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c316
+ bl_0_316 br_0_316 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c316
+ bl_0_316 br_0_316 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c316
+ bl_0_316 br_0_316 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c316
+ bl_0_316 br_0_316 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c316
+ bl_0_316 br_0_316 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c316
+ bl_0_316 br_0_316 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c316
+ bl_0_316 br_0_316 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c316
+ bl_0_316 br_0_316 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c316
+ bl_0_316 br_0_316 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c316
+ bl_0_316 br_0_316 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c316
+ bl_0_316 br_0_316 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c316
+ bl_0_316 br_0_316 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c316
+ bl_0_316 br_0_316 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c316
+ bl_0_316 br_0_316 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c316
+ bl_0_316 br_0_316 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c316
+ bl_0_316 br_0_316 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c316
+ bl_0_316 br_0_316 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c316
+ bl_0_316 br_0_316 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c316
+ bl_0_316 br_0_316 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c316
+ bl_0_316 br_0_316 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c316
+ bl_0_316 br_0_316 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c316
+ bl_0_316 br_0_316 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c316
+ bl_0_316 br_0_316 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c316
+ bl_0_316 br_0_316 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c316
+ bl_0_316 br_0_316 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c316
+ bl_0_316 br_0_316 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c316
+ bl_0_316 br_0_316 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c316
+ bl_0_316 br_0_316 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c316
+ bl_0_316 br_0_316 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c316
+ bl_0_316 br_0_316 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c316
+ bl_0_316 br_0_316 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c316
+ bl_0_316 br_0_316 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c316
+ bl_0_316 br_0_316 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c316
+ bl_0_316 br_0_316 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c316
+ bl_0_316 br_0_316 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c316
+ bl_0_316 br_0_316 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c316
+ bl_0_316 br_0_316 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c316
+ bl_0_316 br_0_316 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c317
+ bl_0_317 br_0_317 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c317
+ bl_0_317 br_0_317 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c317
+ bl_0_317 br_0_317 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c317
+ bl_0_317 br_0_317 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c317
+ bl_0_317 br_0_317 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c317
+ bl_0_317 br_0_317 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c317
+ bl_0_317 br_0_317 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c317
+ bl_0_317 br_0_317 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c317
+ bl_0_317 br_0_317 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c317
+ bl_0_317 br_0_317 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c317
+ bl_0_317 br_0_317 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c317
+ bl_0_317 br_0_317 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c317
+ bl_0_317 br_0_317 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c317
+ bl_0_317 br_0_317 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c317
+ bl_0_317 br_0_317 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c317
+ bl_0_317 br_0_317 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c317
+ bl_0_317 br_0_317 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c317
+ bl_0_317 br_0_317 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c317
+ bl_0_317 br_0_317 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c317
+ bl_0_317 br_0_317 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c317
+ bl_0_317 br_0_317 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c317
+ bl_0_317 br_0_317 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c317
+ bl_0_317 br_0_317 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c317
+ bl_0_317 br_0_317 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c317
+ bl_0_317 br_0_317 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c317
+ bl_0_317 br_0_317 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c317
+ bl_0_317 br_0_317 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c317
+ bl_0_317 br_0_317 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c317
+ bl_0_317 br_0_317 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c317
+ bl_0_317 br_0_317 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c317
+ bl_0_317 br_0_317 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c317
+ bl_0_317 br_0_317 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c317
+ bl_0_317 br_0_317 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c317
+ bl_0_317 br_0_317 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c317
+ bl_0_317 br_0_317 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c317
+ bl_0_317 br_0_317 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c317
+ bl_0_317 br_0_317 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c317
+ bl_0_317 br_0_317 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c317
+ bl_0_317 br_0_317 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c317
+ bl_0_317 br_0_317 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c317
+ bl_0_317 br_0_317 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c317
+ bl_0_317 br_0_317 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c317
+ bl_0_317 br_0_317 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c317
+ bl_0_317 br_0_317 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c317
+ bl_0_317 br_0_317 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c318
+ bl_0_318 br_0_318 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c318
+ bl_0_318 br_0_318 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c318
+ bl_0_318 br_0_318 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c318
+ bl_0_318 br_0_318 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c318
+ bl_0_318 br_0_318 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c318
+ bl_0_318 br_0_318 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c318
+ bl_0_318 br_0_318 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c318
+ bl_0_318 br_0_318 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c318
+ bl_0_318 br_0_318 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c318
+ bl_0_318 br_0_318 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c318
+ bl_0_318 br_0_318 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c318
+ bl_0_318 br_0_318 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c318
+ bl_0_318 br_0_318 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c318
+ bl_0_318 br_0_318 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c318
+ bl_0_318 br_0_318 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c318
+ bl_0_318 br_0_318 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c318
+ bl_0_318 br_0_318 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c318
+ bl_0_318 br_0_318 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c318
+ bl_0_318 br_0_318 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c318
+ bl_0_318 br_0_318 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c318
+ bl_0_318 br_0_318 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c318
+ bl_0_318 br_0_318 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c318
+ bl_0_318 br_0_318 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c318
+ bl_0_318 br_0_318 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c318
+ bl_0_318 br_0_318 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c318
+ bl_0_318 br_0_318 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c318
+ bl_0_318 br_0_318 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c318
+ bl_0_318 br_0_318 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c318
+ bl_0_318 br_0_318 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c318
+ bl_0_318 br_0_318 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c318
+ bl_0_318 br_0_318 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c318
+ bl_0_318 br_0_318 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c318
+ bl_0_318 br_0_318 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c318
+ bl_0_318 br_0_318 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c318
+ bl_0_318 br_0_318 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c318
+ bl_0_318 br_0_318 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c318
+ bl_0_318 br_0_318 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c318
+ bl_0_318 br_0_318 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c318
+ bl_0_318 br_0_318 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c318
+ bl_0_318 br_0_318 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c318
+ bl_0_318 br_0_318 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c318
+ bl_0_318 br_0_318 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c318
+ bl_0_318 br_0_318 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c318
+ bl_0_318 br_0_318 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c318
+ bl_0_318 br_0_318 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c319
+ bl_0_319 br_0_319 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c319
+ bl_0_319 br_0_319 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c319
+ bl_0_319 br_0_319 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c319
+ bl_0_319 br_0_319 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c319
+ bl_0_319 br_0_319 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c319
+ bl_0_319 br_0_319 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c319
+ bl_0_319 br_0_319 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c319
+ bl_0_319 br_0_319 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c319
+ bl_0_319 br_0_319 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c319
+ bl_0_319 br_0_319 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c319
+ bl_0_319 br_0_319 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c319
+ bl_0_319 br_0_319 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c319
+ bl_0_319 br_0_319 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c319
+ bl_0_319 br_0_319 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c319
+ bl_0_319 br_0_319 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c319
+ bl_0_319 br_0_319 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c319
+ bl_0_319 br_0_319 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c319
+ bl_0_319 br_0_319 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c319
+ bl_0_319 br_0_319 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c319
+ bl_0_319 br_0_319 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c319
+ bl_0_319 br_0_319 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c319
+ bl_0_319 br_0_319 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c319
+ bl_0_319 br_0_319 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c319
+ bl_0_319 br_0_319 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c319
+ bl_0_319 br_0_319 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c319
+ bl_0_319 br_0_319 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c319
+ bl_0_319 br_0_319 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c319
+ bl_0_319 br_0_319 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c319
+ bl_0_319 br_0_319 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c319
+ bl_0_319 br_0_319 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c319
+ bl_0_319 br_0_319 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c319
+ bl_0_319 br_0_319 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c319
+ bl_0_319 br_0_319 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c319
+ bl_0_319 br_0_319 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c319
+ bl_0_319 br_0_319 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c319
+ bl_0_319 br_0_319 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c319
+ bl_0_319 br_0_319 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c319
+ bl_0_319 br_0_319 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c319
+ bl_0_319 br_0_319 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c319
+ bl_0_319 br_0_319 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c319
+ bl_0_319 br_0_319 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c319
+ bl_0_319 br_0_319 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c319
+ bl_0_319 br_0_319 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c319
+ bl_0_319 br_0_319 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c319
+ bl_0_319 br_0_319 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c320
+ bl_0_320 br_0_320 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c320
+ bl_0_320 br_0_320 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c320
+ bl_0_320 br_0_320 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c320
+ bl_0_320 br_0_320 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c320
+ bl_0_320 br_0_320 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c320
+ bl_0_320 br_0_320 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c320
+ bl_0_320 br_0_320 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c320
+ bl_0_320 br_0_320 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c320
+ bl_0_320 br_0_320 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c320
+ bl_0_320 br_0_320 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c320
+ bl_0_320 br_0_320 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c320
+ bl_0_320 br_0_320 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c320
+ bl_0_320 br_0_320 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c320
+ bl_0_320 br_0_320 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c320
+ bl_0_320 br_0_320 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c320
+ bl_0_320 br_0_320 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c320
+ bl_0_320 br_0_320 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c320
+ bl_0_320 br_0_320 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c320
+ bl_0_320 br_0_320 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c320
+ bl_0_320 br_0_320 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c320
+ bl_0_320 br_0_320 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c320
+ bl_0_320 br_0_320 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c320
+ bl_0_320 br_0_320 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c320
+ bl_0_320 br_0_320 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c320
+ bl_0_320 br_0_320 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c320
+ bl_0_320 br_0_320 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c320
+ bl_0_320 br_0_320 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c320
+ bl_0_320 br_0_320 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c320
+ bl_0_320 br_0_320 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c320
+ bl_0_320 br_0_320 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c320
+ bl_0_320 br_0_320 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c320
+ bl_0_320 br_0_320 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c320
+ bl_0_320 br_0_320 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c320
+ bl_0_320 br_0_320 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c320
+ bl_0_320 br_0_320 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c320
+ bl_0_320 br_0_320 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c320
+ bl_0_320 br_0_320 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c320
+ bl_0_320 br_0_320 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c320
+ bl_0_320 br_0_320 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c320
+ bl_0_320 br_0_320 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c320
+ bl_0_320 br_0_320 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c320
+ bl_0_320 br_0_320 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c320
+ bl_0_320 br_0_320 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c320
+ bl_0_320 br_0_320 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c320
+ bl_0_320 br_0_320 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c321
+ bl_0_321 br_0_321 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c321
+ bl_0_321 br_0_321 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c321
+ bl_0_321 br_0_321 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c321
+ bl_0_321 br_0_321 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c321
+ bl_0_321 br_0_321 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c321
+ bl_0_321 br_0_321 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c321
+ bl_0_321 br_0_321 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c321
+ bl_0_321 br_0_321 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c321
+ bl_0_321 br_0_321 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c321
+ bl_0_321 br_0_321 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c321
+ bl_0_321 br_0_321 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c321
+ bl_0_321 br_0_321 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c321
+ bl_0_321 br_0_321 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c321
+ bl_0_321 br_0_321 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c321
+ bl_0_321 br_0_321 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c321
+ bl_0_321 br_0_321 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c321
+ bl_0_321 br_0_321 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c321
+ bl_0_321 br_0_321 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c321
+ bl_0_321 br_0_321 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c321
+ bl_0_321 br_0_321 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c321
+ bl_0_321 br_0_321 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c321
+ bl_0_321 br_0_321 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c321
+ bl_0_321 br_0_321 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c321
+ bl_0_321 br_0_321 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c321
+ bl_0_321 br_0_321 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c321
+ bl_0_321 br_0_321 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c321
+ bl_0_321 br_0_321 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c321
+ bl_0_321 br_0_321 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c321
+ bl_0_321 br_0_321 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c321
+ bl_0_321 br_0_321 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c321
+ bl_0_321 br_0_321 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c321
+ bl_0_321 br_0_321 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c321
+ bl_0_321 br_0_321 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c321
+ bl_0_321 br_0_321 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c321
+ bl_0_321 br_0_321 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c321
+ bl_0_321 br_0_321 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c321
+ bl_0_321 br_0_321 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c321
+ bl_0_321 br_0_321 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c321
+ bl_0_321 br_0_321 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c321
+ bl_0_321 br_0_321 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c321
+ bl_0_321 br_0_321 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c321
+ bl_0_321 br_0_321 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c321
+ bl_0_321 br_0_321 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c321
+ bl_0_321 br_0_321 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c321
+ bl_0_321 br_0_321 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c322
+ bl_0_322 br_0_322 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c322
+ bl_0_322 br_0_322 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c322
+ bl_0_322 br_0_322 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c322
+ bl_0_322 br_0_322 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c322
+ bl_0_322 br_0_322 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c322
+ bl_0_322 br_0_322 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c322
+ bl_0_322 br_0_322 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c322
+ bl_0_322 br_0_322 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c322
+ bl_0_322 br_0_322 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c322
+ bl_0_322 br_0_322 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c322
+ bl_0_322 br_0_322 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c322
+ bl_0_322 br_0_322 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c322
+ bl_0_322 br_0_322 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c322
+ bl_0_322 br_0_322 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c322
+ bl_0_322 br_0_322 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c322
+ bl_0_322 br_0_322 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c322
+ bl_0_322 br_0_322 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c322
+ bl_0_322 br_0_322 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c322
+ bl_0_322 br_0_322 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c322
+ bl_0_322 br_0_322 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c322
+ bl_0_322 br_0_322 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c322
+ bl_0_322 br_0_322 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c322
+ bl_0_322 br_0_322 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c322
+ bl_0_322 br_0_322 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c322
+ bl_0_322 br_0_322 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c322
+ bl_0_322 br_0_322 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c322
+ bl_0_322 br_0_322 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c322
+ bl_0_322 br_0_322 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c322
+ bl_0_322 br_0_322 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c322
+ bl_0_322 br_0_322 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c322
+ bl_0_322 br_0_322 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c322
+ bl_0_322 br_0_322 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c322
+ bl_0_322 br_0_322 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c322
+ bl_0_322 br_0_322 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c322
+ bl_0_322 br_0_322 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c322
+ bl_0_322 br_0_322 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c322
+ bl_0_322 br_0_322 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c322
+ bl_0_322 br_0_322 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c322
+ bl_0_322 br_0_322 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c322
+ bl_0_322 br_0_322 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c322
+ bl_0_322 br_0_322 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c322
+ bl_0_322 br_0_322 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c322
+ bl_0_322 br_0_322 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c322
+ bl_0_322 br_0_322 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c322
+ bl_0_322 br_0_322 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c323
+ bl_0_323 br_0_323 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c323
+ bl_0_323 br_0_323 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c323
+ bl_0_323 br_0_323 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c323
+ bl_0_323 br_0_323 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c323
+ bl_0_323 br_0_323 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c323
+ bl_0_323 br_0_323 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c323
+ bl_0_323 br_0_323 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c323
+ bl_0_323 br_0_323 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c323
+ bl_0_323 br_0_323 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c323
+ bl_0_323 br_0_323 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c323
+ bl_0_323 br_0_323 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c323
+ bl_0_323 br_0_323 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c323
+ bl_0_323 br_0_323 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c323
+ bl_0_323 br_0_323 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c323
+ bl_0_323 br_0_323 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c323
+ bl_0_323 br_0_323 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c323
+ bl_0_323 br_0_323 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c323
+ bl_0_323 br_0_323 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c323
+ bl_0_323 br_0_323 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c323
+ bl_0_323 br_0_323 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c323
+ bl_0_323 br_0_323 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c323
+ bl_0_323 br_0_323 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c323
+ bl_0_323 br_0_323 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c323
+ bl_0_323 br_0_323 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c323
+ bl_0_323 br_0_323 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c323
+ bl_0_323 br_0_323 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c323
+ bl_0_323 br_0_323 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c323
+ bl_0_323 br_0_323 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c323
+ bl_0_323 br_0_323 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c323
+ bl_0_323 br_0_323 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c323
+ bl_0_323 br_0_323 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c323
+ bl_0_323 br_0_323 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c323
+ bl_0_323 br_0_323 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c323
+ bl_0_323 br_0_323 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c323
+ bl_0_323 br_0_323 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c323
+ bl_0_323 br_0_323 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c323
+ bl_0_323 br_0_323 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c323
+ bl_0_323 br_0_323 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c323
+ bl_0_323 br_0_323 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c323
+ bl_0_323 br_0_323 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c323
+ bl_0_323 br_0_323 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c323
+ bl_0_323 br_0_323 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c323
+ bl_0_323 br_0_323 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c323
+ bl_0_323 br_0_323 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c323
+ bl_0_323 br_0_323 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c324
+ bl_0_324 br_0_324 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c324
+ bl_0_324 br_0_324 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c324
+ bl_0_324 br_0_324 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c324
+ bl_0_324 br_0_324 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c324
+ bl_0_324 br_0_324 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c324
+ bl_0_324 br_0_324 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c324
+ bl_0_324 br_0_324 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c324
+ bl_0_324 br_0_324 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c324
+ bl_0_324 br_0_324 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c324
+ bl_0_324 br_0_324 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c324
+ bl_0_324 br_0_324 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c324
+ bl_0_324 br_0_324 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c324
+ bl_0_324 br_0_324 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c324
+ bl_0_324 br_0_324 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c324
+ bl_0_324 br_0_324 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c324
+ bl_0_324 br_0_324 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c324
+ bl_0_324 br_0_324 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c324
+ bl_0_324 br_0_324 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c324
+ bl_0_324 br_0_324 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c324
+ bl_0_324 br_0_324 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c324
+ bl_0_324 br_0_324 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c324
+ bl_0_324 br_0_324 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c324
+ bl_0_324 br_0_324 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c324
+ bl_0_324 br_0_324 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c324
+ bl_0_324 br_0_324 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c324
+ bl_0_324 br_0_324 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c324
+ bl_0_324 br_0_324 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c324
+ bl_0_324 br_0_324 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c324
+ bl_0_324 br_0_324 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c324
+ bl_0_324 br_0_324 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c324
+ bl_0_324 br_0_324 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c324
+ bl_0_324 br_0_324 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c324
+ bl_0_324 br_0_324 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c324
+ bl_0_324 br_0_324 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c324
+ bl_0_324 br_0_324 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c324
+ bl_0_324 br_0_324 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c324
+ bl_0_324 br_0_324 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c324
+ bl_0_324 br_0_324 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c324
+ bl_0_324 br_0_324 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c324
+ bl_0_324 br_0_324 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c324
+ bl_0_324 br_0_324 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c324
+ bl_0_324 br_0_324 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c324
+ bl_0_324 br_0_324 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c324
+ bl_0_324 br_0_324 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c324
+ bl_0_324 br_0_324 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c325
+ bl_0_325 br_0_325 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c325
+ bl_0_325 br_0_325 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c325
+ bl_0_325 br_0_325 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c325
+ bl_0_325 br_0_325 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c325
+ bl_0_325 br_0_325 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c325
+ bl_0_325 br_0_325 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c325
+ bl_0_325 br_0_325 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c325
+ bl_0_325 br_0_325 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c325
+ bl_0_325 br_0_325 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c325
+ bl_0_325 br_0_325 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c325
+ bl_0_325 br_0_325 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c325
+ bl_0_325 br_0_325 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c325
+ bl_0_325 br_0_325 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c325
+ bl_0_325 br_0_325 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c325
+ bl_0_325 br_0_325 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c325
+ bl_0_325 br_0_325 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c325
+ bl_0_325 br_0_325 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c325
+ bl_0_325 br_0_325 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c325
+ bl_0_325 br_0_325 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c325
+ bl_0_325 br_0_325 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c325
+ bl_0_325 br_0_325 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c325
+ bl_0_325 br_0_325 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c325
+ bl_0_325 br_0_325 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c325
+ bl_0_325 br_0_325 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c325
+ bl_0_325 br_0_325 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c325
+ bl_0_325 br_0_325 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c325
+ bl_0_325 br_0_325 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c325
+ bl_0_325 br_0_325 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c325
+ bl_0_325 br_0_325 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c325
+ bl_0_325 br_0_325 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c325
+ bl_0_325 br_0_325 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c325
+ bl_0_325 br_0_325 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c325
+ bl_0_325 br_0_325 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c325
+ bl_0_325 br_0_325 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c325
+ bl_0_325 br_0_325 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c325
+ bl_0_325 br_0_325 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c325
+ bl_0_325 br_0_325 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c325
+ bl_0_325 br_0_325 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c325
+ bl_0_325 br_0_325 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c325
+ bl_0_325 br_0_325 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c325
+ bl_0_325 br_0_325 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c325
+ bl_0_325 br_0_325 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c325
+ bl_0_325 br_0_325 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c325
+ bl_0_325 br_0_325 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c325
+ bl_0_325 br_0_325 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c326
+ bl_0_326 br_0_326 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c326
+ bl_0_326 br_0_326 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c326
+ bl_0_326 br_0_326 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c326
+ bl_0_326 br_0_326 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c326
+ bl_0_326 br_0_326 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c326
+ bl_0_326 br_0_326 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c326
+ bl_0_326 br_0_326 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c326
+ bl_0_326 br_0_326 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c326
+ bl_0_326 br_0_326 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c326
+ bl_0_326 br_0_326 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c326
+ bl_0_326 br_0_326 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c326
+ bl_0_326 br_0_326 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c326
+ bl_0_326 br_0_326 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c326
+ bl_0_326 br_0_326 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c326
+ bl_0_326 br_0_326 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c326
+ bl_0_326 br_0_326 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c326
+ bl_0_326 br_0_326 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c326
+ bl_0_326 br_0_326 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c326
+ bl_0_326 br_0_326 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c326
+ bl_0_326 br_0_326 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c326
+ bl_0_326 br_0_326 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c326
+ bl_0_326 br_0_326 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c326
+ bl_0_326 br_0_326 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c326
+ bl_0_326 br_0_326 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c326
+ bl_0_326 br_0_326 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c326
+ bl_0_326 br_0_326 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c326
+ bl_0_326 br_0_326 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c326
+ bl_0_326 br_0_326 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c326
+ bl_0_326 br_0_326 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c326
+ bl_0_326 br_0_326 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c326
+ bl_0_326 br_0_326 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c326
+ bl_0_326 br_0_326 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c326
+ bl_0_326 br_0_326 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c326
+ bl_0_326 br_0_326 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c326
+ bl_0_326 br_0_326 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c326
+ bl_0_326 br_0_326 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c326
+ bl_0_326 br_0_326 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c326
+ bl_0_326 br_0_326 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c326
+ bl_0_326 br_0_326 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c326
+ bl_0_326 br_0_326 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c326
+ bl_0_326 br_0_326 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c326
+ bl_0_326 br_0_326 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c326
+ bl_0_326 br_0_326 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c326
+ bl_0_326 br_0_326 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c326
+ bl_0_326 br_0_326 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c327
+ bl_0_327 br_0_327 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c327
+ bl_0_327 br_0_327 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c327
+ bl_0_327 br_0_327 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c327
+ bl_0_327 br_0_327 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c327
+ bl_0_327 br_0_327 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c327
+ bl_0_327 br_0_327 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c327
+ bl_0_327 br_0_327 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c327
+ bl_0_327 br_0_327 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c327
+ bl_0_327 br_0_327 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c327
+ bl_0_327 br_0_327 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c327
+ bl_0_327 br_0_327 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c327
+ bl_0_327 br_0_327 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c327
+ bl_0_327 br_0_327 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c327
+ bl_0_327 br_0_327 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c327
+ bl_0_327 br_0_327 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c327
+ bl_0_327 br_0_327 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c327
+ bl_0_327 br_0_327 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c327
+ bl_0_327 br_0_327 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c327
+ bl_0_327 br_0_327 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c327
+ bl_0_327 br_0_327 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c327
+ bl_0_327 br_0_327 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c327
+ bl_0_327 br_0_327 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c327
+ bl_0_327 br_0_327 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c327
+ bl_0_327 br_0_327 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c327
+ bl_0_327 br_0_327 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c327
+ bl_0_327 br_0_327 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c327
+ bl_0_327 br_0_327 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c327
+ bl_0_327 br_0_327 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c327
+ bl_0_327 br_0_327 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c327
+ bl_0_327 br_0_327 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c327
+ bl_0_327 br_0_327 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c327
+ bl_0_327 br_0_327 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c327
+ bl_0_327 br_0_327 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c327
+ bl_0_327 br_0_327 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c327
+ bl_0_327 br_0_327 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c327
+ bl_0_327 br_0_327 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c327
+ bl_0_327 br_0_327 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c327
+ bl_0_327 br_0_327 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c327
+ bl_0_327 br_0_327 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c327
+ bl_0_327 br_0_327 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c327
+ bl_0_327 br_0_327 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c327
+ bl_0_327 br_0_327 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c327
+ bl_0_327 br_0_327 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c327
+ bl_0_327 br_0_327 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c327
+ bl_0_327 br_0_327 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c328
+ bl_0_328 br_0_328 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c328
+ bl_0_328 br_0_328 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c328
+ bl_0_328 br_0_328 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c328
+ bl_0_328 br_0_328 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c328
+ bl_0_328 br_0_328 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c328
+ bl_0_328 br_0_328 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c328
+ bl_0_328 br_0_328 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c328
+ bl_0_328 br_0_328 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c328
+ bl_0_328 br_0_328 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c328
+ bl_0_328 br_0_328 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c328
+ bl_0_328 br_0_328 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c328
+ bl_0_328 br_0_328 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c328
+ bl_0_328 br_0_328 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c328
+ bl_0_328 br_0_328 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c328
+ bl_0_328 br_0_328 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c328
+ bl_0_328 br_0_328 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c328
+ bl_0_328 br_0_328 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c328
+ bl_0_328 br_0_328 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c328
+ bl_0_328 br_0_328 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c328
+ bl_0_328 br_0_328 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c328
+ bl_0_328 br_0_328 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c328
+ bl_0_328 br_0_328 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c328
+ bl_0_328 br_0_328 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c328
+ bl_0_328 br_0_328 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c328
+ bl_0_328 br_0_328 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c328
+ bl_0_328 br_0_328 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c328
+ bl_0_328 br_0_328 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c328
+ bl_0_328 br_0_328 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c328
+ bl_0_328 br_0_328 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c328
+ bl_0_328 br_0_328 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c328
+ bl_0_328 br_0_328 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c328
+ bl_0_328 br_0_328 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c328
+ bl_0_328 br_0_328 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c328
+ bl_0_328 br_0_328 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c328
+ bl_0_328 br_0_328 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c328
+ bl_0_328 br_0_328 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c328
+ bl_0_328 br_0_328 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c328
+ bl_0_328 br_0_328 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c328
+ bl_0_328 br_0_328 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c328
+ bl_0_328 br_0_328 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c328
+ bl_0_328 br_0_328 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c328
+ bl_0_328 br_0_328 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c328
+ bl_0_328 br_0_328 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c328
+ bl_0_328 br_0_328 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c328
+ bl_0_328 br_0_328 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c329
+ bl_0_329 br_0_329 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c329
+ bl_0_329 br_0_329 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c329
+ bl_0_329 br_0_329 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c329
+ bl_0_329 br_0_329 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c329
+ bl_0_329 br_0_329 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c329
+ bl_0_329 br_0_329 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c329
+ bl_0_329 br_0_329 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c329
+ bl_0_329 br_0_329 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c329
+ bl_0_329 br_0_329 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c329
+ bl_0_329 br_0_329 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c329
+ bl_0_329 br_0_329 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c329
+ bl_0_329 br_0_329 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c329
+ bl_0_329 br_0_329 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c329
+ bl_0_329 br_0_329 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c329
+ bl_0_329 br_0_329 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c329
+ bl_0_329 br_0_329 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c329
+ bl_0_329 br_0_329 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c329
+ bl_0_329 br_0_329 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c329
+ bl_0_329 br_0_329 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c329
+ bl_0_329 br_0_329 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c329
+ bl_0_329 br_0_329 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c329
+ bl_0_329 br_0_329 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c329
+ bl_0_329 br_0_329 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c329
+ bl_0_329 br_0_329 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c329
+ bl_0_329 br_0_329 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c329
+ bl_0_329 br_0_329 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c329
+ bl_0_329 br_0_329 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c329
+ bl_0_329 br_0_329 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c329
+ bl_0_329 br_0_329 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c329
+ bl_0_329 br_0_329 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c329
+ bl_0_329 br_0_329 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c329
+ bl_0_329 br_0_329 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c329
+ bl_0_329 br_0_329 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c329
+ bl_0_329 br_0_329 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c329
+ bl_0_329 br_0_329 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c329
+ bl_0_329 br_0_329 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c329
+ bl_0_329 br_0_329 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c329
+ bl_0_329 br_0_329 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c329
+ bl_0_329 br_0_329 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c329
+ bl_0_329 br_0_329 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c329
+ bl_0_329 br_0_329 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c329
+ bl_0_329 br_0_329 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c329
+ bl_0_329 br_0_329 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c329
+ bl_0_329 br_0_329 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c329
+ bl_0_329 br_0_329 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c330
+ bl_0_330 br_0_330 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c330
+ bl_0_330 br_0_330 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c330
+ bl_0_330 br_0_330 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c330
+ bl_0_330 br_0_330 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c330
+ bl_0_330 br_0_330 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c330
+ bl_0_330 br_0_330 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c330
+ bl_0_330 br_0_330 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c330
+ bl_0_330 br_0_330 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c330
+ bl_0_330 br_0_330 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c330
+ bl_0_330 br_0_330 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c330
+ bl_0_330 br_0_330 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c330
+ bl_0_330 br_0_330 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c330
+ bl_0_330 br_0_330 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c330
+ bl_0_330 br_0_330 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c330
+ bl_0_330 br_0_330 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c330
+ bl_0_330 br_0_330 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c330
+ bl_0_330 br_0_330 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c330
+ bl_0_330 br_0_330 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c330
+ bl_0_330 br_0_330 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c330
+ bl_0_330 br_0_330 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c330
+ bl_0_330 br_0_330 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c330
+ bl_0_330 br_0_330 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c330
+ bl_0_330 br_0_330 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c330
+ bl_0_330 br_0_330 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c330
+ bl_0_330 br_0_330 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c330
+ bl_0_330 br_0_330 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c330
+ bl_0_330 br_0_330 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c330
+ bl_0_330 br_0_330 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c330
+ bl_0_330 br_0_330 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c330
+ bl_0_330 br_0_330 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c330
+ bl_0_330 br_0_330 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c330
+ bl_0_330 br_0_330 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c330
+ bl_0_330 br_0_330 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c330
+ bl_0_330 br_0_330 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c330
+ bl_0_330 br_0_330 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c330
+ bl_0_330 br_0_330 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c330
+ bl_0_330 br_0_330 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c330
+ bl_0_330 br_0_330 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c330
+ bl_0_330 br_0_330 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c330
+ bl_0_330 br_0_330 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c330
+ bl_0_330 br_0_330 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c330
+ bl_0_330 br_0_330 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c330
+ bl_0_330 br_0_330 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c330
+ bl_0_330 br_0_330 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c330
+ bl_0_330 br_0_330 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c331
+ bl_0_331 br_0_331 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c331
+ bl_0_331 br_0_331 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c331
+ bl_0_331 br_0_331 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c331
+ bl_0_331 br_0_331 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c331
+ bl_0_331 br_0_331 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c331
+ bl_0_331 br_0_331 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c331
+ bl_0_331 br_0_331 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c331
+ bl_0_331 br_0_331 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c331
+ bl_0_331 br_0_331 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c331
+ bl_0_331 br_0_331 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c331
+ bl_0_331 br_0_331 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c331
+ bl_0_331 br_0_331 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c331
+ bl_0_331 br_0_331 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c331
+ bl_0_331 br_0_331 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c331
+ bl_0_331 br_0_331 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c331
+ bl_0_331 br_0_331 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c331
+ bl_0_331 br_0_331 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c331
+ bl_0_331 br_0_331 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c331
+ bl_0_331 br_0_331 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c331
+ bl_0_331 br_0_331 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c331
+ bl_0_331 br_0_331 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c331
+ bl_0_331 br_0_331 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c331
+ bl_0_331 br_0_331 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c331
+ bl_0_331 br_0_331 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c331
+ bl_0_331 br_0_331 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c331
+ bl_0_331 br_0_331 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c331
+ bl_0_331 br_0_331 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c331
+ bl_0_331 br_0_331 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c331
+ bl_0_331 br_0_331 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c331
+ bl_0_331 br_0_331 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c331
+ bl_0_331 br_0_331 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c331
+ bl_0_331 br_0_331 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c331
+ bl_0_331 br_0_331 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c331
+ bl_0_331 br_0_331 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c331
+ bl_0_331 br_0_331 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c331
+ bl_0_331 br_0_331 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c331
+ bl_0_331 br_0_331 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c331
+ bl_0_331 br_0_331 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c331
+ bl_0_331 br_0_331 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c331
+ bl_0_331 br_0_331 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c331
+ bl_0_331 br_0_331 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c331
+ bl_0_331 br_0_331 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c331
+ bl_0_331 br_0_331 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c331
+ bl_0_331 br_0_331 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c331
+ bl_0_331 br_0_331 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c332
+ bl_0_332 br_0_332 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c332
+ bl_0_332 br_0_332 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c332
+ bl_0_332 br_0_332 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c332
+ bl_0_332 br_0_332 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c332
+ bl_0_332 br_0_332 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c332
+ bl_0_332 br_0_332 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c332
+ bl_0_332 br_0_332 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c332
+ bl_0_332 br_0_332 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c332
+ bl_0_332 br_0_332 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c332
+ bl_0_332 br_0_332 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c332
+ bl_0_332 br_0_332 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c332
+ bl_0_332 br_0_332 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c332
+ bl_0_332 br_0_332 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c332
+ bl_0_332 br_0_332 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c332
+ bl_0_332 br_0_332 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c332
+ bl_0_332 br_0_332 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c332
+ bl_0_332 br_0_332 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c332
+ bl_0_332 br_0_332 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c332
+ bl_0_332 br_0_332 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c332
+ bl_0_332 br_0_332 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c332
+ bl_0_332 br_0_332 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c332
+ bl_0_332 br_0_332 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c332
+ bl_0_332 br_0_332 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c332
+ bl_0_332 br_0_332 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c332
+ bl_0_332 br_0_332 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c332
+ bl_0_332 br_0_332 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c332
+ bl_0_332 br_0_332 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c332
+ bl_0_332 br_0_332 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c332
+ bl_0_332 br_0_332 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c332
+ bl_0_332 br_0_332 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c332
+ bl_0_332 br_0_332 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c332
+ bl_0_332 br_0_332 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c332
+ bl_0_332 br_0_332 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c332
+ bl_0_332 br_0_332 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c332
+ bl_0_332 br_0_332 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c332
+ bl_0_332 br_0_332 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c332
+ bl_0_332 br_0_332 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c332
+ bl_0_332 br_0_332 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c332
+ bl_0_332 br_0_332 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c332
+ bl_0_332 br_0_332 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c332
+ bl_0_332 br_0_332 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c332
+ bl_0_332 br_0_332 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c332
+ bl_0_332 br_0_332 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c332
+ bl_0_332 br_0_332 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c332
+ bl_0_332 br_0_332 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c333
+ bl_0_333 br_0_333 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c333
+ bl_0_333 br_0_333 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c333
+ bl_0_333 br_0_333 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c333
+ bl_0_333 br_0_333 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c333
+ bl_0_333 br_0_333 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c333
+ bl_0_333 br_0_333 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c333
+ bl_0_333 br_0_333 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c333
+ bl_0_333 br_0_333 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c333
+ bl_0_333 br_0_333 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c333
+ bl_0_333 br_0_333 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c333
+ bl_0_333 br_0_333 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c333
+ bl_0_333 br_0_333 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c333
+ bl_0_333 br_0_333 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c333
+ bl_0_333 br_0_333 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c333
+ bl_0_333 br_0_333 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c333
+ bl_0_333 br_0_333 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c333
+ bl_0_333 br_0_333 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c333
+ bl_0_333 br_0_333 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c333
+ bl_0_333 br_0_333 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c333
+ bl_0_333 br_0_333 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c333
+ bl_0_333 br_0_333 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c333
+ bl_0_333 br_0_333 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c333
+ bl_0_333 br_0_333 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c333
+ bl_0_333 br_0_333 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c333
+ bl_0_333 br_0_333 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c333
+ bl_0_333 br_0_333 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c333
+ bl_0_333 br_0_333 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c333
+ bl_0_333 br_0_333 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c333
+ bl_0_333 br_0_333 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c333
+ bl_0_333 br_0_333 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c333
+ bl_0_333 br_0_333 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c333
+ bl_0_333 br_0_333 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c333
+ bl_0_333 br_0_333 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c333
+ bl_0_333 br_0_333 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c333
+ bl_0_333 br_0_333 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c333
+ bl_0_333 br_0_333 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c333
+ bl_0_333 br_0_333 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c333
+ bl_0_333 br_0_333 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c333
+ bl_0_333 br_0_333 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c333
+ bl_0_333 br_0_333 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c333
+ bl_0_333 br_0_333 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c333
+ bl_0_333 br_0_333 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c333
+ bl_0_333 br_0_333 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c333
+ bl_0_333 br_0_333 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c333
+ bl_0_333 br_0_333 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c334
+ bl_0_334 br_0_334 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c334
+ bl_0_334 br_0_334 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c334
+ bl_0_334 br_0_334 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c334
+ bl_0_334 br_0_334 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c334
+ bl_0_334 br_0_334 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c334
+ bl_0_334 br_0_334 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c334
+ bl_0_334 br_0_334 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c334
+ bl_0_334 br_0_334 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c334
+ bl_0_334 br_0_334 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c334
+ bl_0_334 br_0_334 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c334
+ bl_0_334 br_0_334 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c334
+ bl_0_334 br_0_334 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c334
+ bl_0_334 br_0_334 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c334
+ bl_0_334 br_0_334 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c334
+ bl_0_334 br_0_334 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c334
+ bl_0_334 br_0_334 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c334
+ bl_0_334 br_0_334 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c334
+ bl_0_334 br_0_334 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c334
+ bl_0_334 br_0_334 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c334
+ bl_0_334 br_0_334 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c334
+ bl_0_334 br_0_334 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c334
+ bl_0_334 br_0_334 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c334
+ bl_0_334 br_0_334 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c334
+ bl_0_334 br_0_334 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c334
+ bl_0_334 br_0_334 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c334
+ bl_0_334 br_0_334 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c334
+ bl_0_334 br_0_334 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c334
+ bl_0_334 br_0_334 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c334
+ bl_0_334 br_0_334 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c334
+ bl_0_334 br_0_334 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c334
+ bl_0_334 br_0_334 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c334
+ bl_0_334 br_0_334 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c334
+ bl_0_334 br_0_334 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c334
+ bl_0_334 br_0_334 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c334
+ bl_0_334 br_0_334 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c334
+ bl_0_334 br_0_334 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c334
+ bl_0_334 br_0_334 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c334
+ bl_0_334 br_0_334 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c334
+ bl_0_334 br_0_334 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c334
+ bl_0_334 br_0_334 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c334
+ bl_0_334 br_0_334 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c334
+ bl_0_334 br_0_334 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c334
+ bl_0_334 br_0_334 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c334
+ bl_0_334 br_0_334 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c334
+ bl_0_334 br_0_334 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c335
+ bl_0_335 br_0_335 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c335
+ bl_0_335 br_0_335 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c335
+ bl_0_335 br_0_335 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c335
+ bl_0_335 br_0_335 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c335
+ bl_0_335 br_0_335 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c335
+ bl_0_335 br_0_335 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c335
+ bl_0_335 br_0_335 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c335
+ bl_0_335 br_0_335 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c335
+ bl_0_335 br_0_335 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c335
+ bl_0_335 br_0_335 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c335
+ bl_0_335 br_0_335 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c335
+ bl_0_335 br_0_335 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c335
+ bl_0_335 br_0_335 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c335
+ bl_0_335 br_0_335 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c335
+ bl_0_335 br_0_335 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c335
+ bl_0_335 br_0_335 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c335
+ bl_0_335 br_0_335 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c335
+ bl_0_335 br_0_335 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c335
+ bl_0_335 br_0_335 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c335
+ bl_0_335 br_0_335 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c335
+ bl_0_335 br_0_335 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c335
+ bl_0_335 br_0_335 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c335
+ bl_0_335 br_0_335 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c335
+ bl_0_335 br_0_335 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c335
+ bl_0_335 br_0_335 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c335
+ bl_0_335 br_0_335 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c335
+ bl_0_335 br_0_335 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c335
+ bl_0_335 br_0_335 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c335
+ bl_0_335 br_0_335 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c335
+ bl_0_335 br_0_335 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c335
+ bl_0_335 br_0_335 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c335
+ bl_0_335 br_0_335 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c335
+ bl_0_335 br_0_335 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c335
+ bl_0_335 br_0_335 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c335
+ bl_0_335 br_0_335 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c335
+ bl_0_335 br_0_335 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c335
+ bl_0_335 br_0_335 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c335
+ bl_0_335 br_0_335 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c335
+ bl_0_335 br_0_335 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c335
+ bl_0_335 br_0_335 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c335
+ bl_0_335 br_0_335 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c335
+ bl_0_335 br_0_335 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c335
+ bl_0_335 br_0_335 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c335
+ bl_0_335 br_0_335 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c335
+ bl_0_335 br_0_335 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c336
+ bl_0_336 br_0_336 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c336
+ bl_0_336 br_0_336 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c336
+ bl_0_336 br_0_336 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c336
+ bl_0_336 br_0_336 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c336
+ bl_0_336 br_0_336 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c336
+ bl_0_336 br_0_336 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c336
+ bl_0_336 br_0_336 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c336
+ bl_0_336 br_0_336 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c336
+ bl_0_336 br_0_336 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c336
+ bl_0_336 br_0_336 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c336
+ bl_0_336 br_0_336 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c336
+ bl_0_336 br_0_336 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c336
+ bl_0_336 br_0_336 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c336
+ bl_0_336 br_0_336 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c336
+ bl_0_336 br_0_336 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c336
+ bl_0_336 br_0_336 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c336
+ bl_0_336 br_0_336 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c336
+ bl_0_336 br_0_336 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c336
+ bl_0_336 br_0_336 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c336
+ bl_0_336 br_0_336 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c336
+ bl_0_336 br_0_336 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c336
+ bl_0_336 br_0_336 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c336
+ bl_0_336 br_0_336 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c336
+ bl_0_336 br_0_336 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c336
+ bl_0_336 br_0_336 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c336
+ bl_0_336 br_0_336 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c336
+ bl_0_336 br_0_336 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c336
+ bl_0_336 br_0_336 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c336
+ bl_0_336 br_0_336 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c336
+ bl_0_336 br_0_336 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c336
+ bl_0_336 br_0_336 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c336
+ bl_0_336 br_0_336 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c336
+ bl_0_336 br_0_336 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c336
+ bl_0_336 br_0_336 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c336
+ bl_0_336 br_0_336 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c336
+ bl_0_336 br_0_336 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c336
+ bl_0_336 br_0_336 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c336
+ bl_0_336 br_0_336 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c336
+ bl_0_336 br_0_336 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c336
+ bl_0_336 br_0_336 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c336
+ bl_0_336 br_0_336 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c336
+ bl_0_336 br_0_336 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c336
+ bl_0_336 br_0_336 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c336
+ bl_0_336 br_0_336 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c336
+ bl_0_336 br_0_336 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c337
+ bl_0_337 br_0_337 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c337
+ bl_0_337 br_0_337 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c337
+ bl_0_337 br_0_337 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c337
+ bl_0_337 br_0_337 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c337
+ bl_0_337 br_0_337 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c337
+ bl_0_337 br_0_337 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c337
+ bl_0_337 br_0_337 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c337
+ bl_0_337 br_0_337 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c337
+ bl_0_337 br_0_337 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c337
+ bl_0_337 br_0_337 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c337
+ bl_0_337 br_0_337 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c337
+ bl_0_337 br_0_337 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c337
+ bl_0_337 br_0_337 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c337
+ bl_0_337 br_0_337 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c337
+ bl_0_337 br_0_337 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c337
+ bl_0_337 br_0_337 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c337
+ bl_0_337 br_0_337 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c337
+ bl_0_337 br_0_337 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c337
+ bl_0_337 br_0_337 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c337
+ bl_0_337 br_0_337 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c337
+ bl_0_337 br_0_337 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c337
+ bl_0_337 br_0_337 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c337
+ bl_0_337 br_0_337 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c337
+ bl_0_337 br_0_337 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c337
+ bl_0_337 br_0_337 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c337
+ bl_0_337 br_0_337 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c337
+ bl_0_337 br_0_337 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c337
+ bl_0_337 br_0_337 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c337
+ bl_0_337 br_0_337 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c337
+ bl_0_337 br_0_337 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c337
+ bl_0_337 br_0_337 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c337
+ bl_0_337 br_0_337 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c337
+ bl_0_337 br_0_337 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c337
+ bl_0_337 br_0_337 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c337
+ bl_0_337 br_0_337 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c337
+ bl_0_337 br_0_337 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c337
+ bl_0_337 br_0_337 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c337
+ bl_0_337 br_0_337 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c337
+ bl_0_337 br_0_337 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c337
+ bl_0_337 br_0_337 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c337
+ bl_0_337 br_0_337 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c337
+ bl_0_337 br_0_337 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c337
+ bl_0_337 br_0_337 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c337
+ bl_0_337 br_0_337 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c337
+ bl_0_337 br_0_337 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c338
+ bl_0_338 br_0_338 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c338
+ bl_0_338 br_0_338 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c338
+ bl_0_338 br_0_338 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c338
+ bl_0_338 br_0_338 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c338
+ bl_0_338 br_0_338 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c338
+ bl_0_338 br_0_338 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c338
+ bl_0_338 br_0_338 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c338
+ bl_0_338 br_0_338 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c338
+ bl_0_338 br_0_338 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c338
+ bl_0_338 br_0_338 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c338
+ bl_0_338 br_0_338 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c338
+ bl_0_338 br_0_338 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c338
+ bl_0_338 br_0_338 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c338
+ bl_0_338 br_0_338 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c338
+ bl_0_338 br_0_338 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c338
+ bl_0_338 br_0_338 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c338
+ bl_0_338 br_0_338 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c338
+ bl_0_338 br_0_338 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c338
+ bl_0_338 br_0_338 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c338
+ bl_0_338 br_0_338 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c338
+ bl_0_338 br_0_338 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c338
+ bl_0_338 br_0_338 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c338
+ bl_0_338 br_0_338 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c338
+ bl_0_338 br_0_338 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c338
+ bl_0_338 br_0_338 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c338
+ bl_0_338 br_0_338 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c338
+ bl_0_338 br_0_338 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c338
+ bl_0_338 br_0_338 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c338
+ bl_0_338 br_0_338 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c338
+ bl_0_338 br_0_338 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c338
+ bl_0_338 br_0_338 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c338
+ bl_0_338 br_0_338 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c338
+ bl_0_338 br_0_338 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c338
+ bl_0_338 br_0_338 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c338
+ bl_0_338 br_0_338 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c338
+ bl_0_338 br_0_338 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c338
+ bl_0_338 br_0_338 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c338
+ bl_0_338 br_0_338 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c338
+ bl_0_338 br_0_338 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c338
+ bl_0_338 br_0_338 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c338
+ bl_0_338 br_0_338 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c338
+ bl_0_338 br_0_338 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c338
+ bl_0_338 br_0_338 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c338
+ bl_0_338 br_0_338 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c338
+ bl_0_338 br_0_338 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c339
+ bl_0_339 br_0_339 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c339
+ bl_0_339 br_0_339 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c339
+ bl_0_339 br_0_339 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c339
+ bl_0_339 br_0_339 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c339
+ bl_0_339 br_0_339 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c339
+ bl_0_339 br_0_339 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c339
+ bl_0_339 br_0_339 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c339
+ bl_0_339 br_0_339 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c339
+ bl_0_339 br_0_339 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c339
+ bl_0_339 br_0_339 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c339
+ bl_0_339 br_0_339 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c339
+ bl_0_339 br_0_339 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c339
+ bl_0_339 br_0_339 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c339
+ bl_0_339 br_0_339 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c339
+ bl_0_339 br_0_339 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c339
+ bl_0_339 br_0_339 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c339
+ bl_0_339 br_0_339 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c339
+ bl_0_339 br_0_339 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c339
+ bl_0_339 br_0_339 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c339
+ bl_0_339 br_0_339 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c339
+ bl_0_339 br_0_339 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c339
+ bl_0_339 br_0_339 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c339
+ bl_0_339 br_0_339 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c339
+ bl_0_339 br_0_339 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c339
+ bl_0_339 br_0_339 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c339
+ bl_0_339 br_0_339 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c339
+ bl_0_339 br_0_339 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c339
+ bl_0_339 br_0_339 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c339
+ bl_0_339 br_0_339 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c339
+ bl_0_339 br_0_339 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c339
+ bl_0_339 br_0_339 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c339
+ bl_0_339 br_0_339 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c339
+ bl_0_339 br_0_339 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c339
+ bl_0_339 br_0_339 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c339
+ bl_0_339 br_0_339 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c339
+ bl_0_339 br_0_339 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c339
+ bl_0_339 br_0_339 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c339
+ bl_0_339 br_0_339 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c339
+ bl_0_339 br_0_339 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c339
+ bl_0_339 br_0_339 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c339
+ bl_0_339 br_0_339 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c339
+ bl_0_339 br_0_339 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c339
+ bl_0_339 br_0_339 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c339
+ bl_0_339 br_0_339 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c339
+ bl_0_339 br_0_339 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c340
+ bl_0_340 br_0_340 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c340
+ bl_0_340 br_0_340 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c340
+ bl_0_340 br_0_340 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c340
+ bl_0_340 br_0_340 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c340
+ bl_0_340 br_0_340 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c340
+ bl_0_340 br_0_340 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c340
+ bl_0_340 br_0_340 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c340
+ bl_0_340 br_0_340 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c340
+ bl_0_340 br_0_340 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c340
+ bl_0_340 br_0_340 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c340
+ bl_0_340 br_0_340 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c340
+ bl_0_340 br_0_340 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c340
+ bl_0_340 br_0_340 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c340
+ bl_0_340 br_0_340 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c340
+ bl_0_340 br_0_340 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c340
+ bl_0_340 br_0_340 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c340
+ bl_0_340 br_0_340 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c340
+ bl_0_340 br_0_340 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c340
+ bl_0_340 br_0_340 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c340
+ bl_0_340 br_0_340 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c340
+ bl_0_340 br_0_340 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c340
+ bl_0_340 br_0_340 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c340
+ bl_0_340 br_0_340 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c340
+ bl_0_340 br_0_340 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c340
+ bl_0_340 br_0_340 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c340
+ bl_0_340 br_0_340 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c340
+ bl_0_340 br_0_340 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c340
+ bl_0_340 br_0_340 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c340
+ bl_0_340 br_0_340 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c340
+ bl_0_340 br_0_340 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c340
+ bl_0_340 br_0_340 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c340
+ bl_0_340 br_0_340 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c340
+ bl_0_340 br_0_340 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c340
+ bl_0_340 br_0_340 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c340
+ bl_0_340 br_0_340 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c340
+ bl_0_340 br_0_340 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c340
+ bl_0_340 br_0_340 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c340
+ bl_0_340 br_0_340 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c340
+ bl_0_340 br_0_340 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c340
+ bl_0_340 br_0_340 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c340
+ bl_0_340 br_0_340 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c340
+ bl_0_340 br_0_340 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c340
+ bl_0_340 br_0_340 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c340
+ bl_0_340 br_0_340 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c340
+ bl_0_340 br_0_340 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c341
+ bl_0_341 br_0_341 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c341
+ bl_0_341 br_0_341 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c341
+ bl_0_341 br_0_341 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c341
+ bl_0_341 br_0_341 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c341
+ bl_0_341 br_0_341 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c341
+ bl_0_341 br_0_341 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c341
+ bl_0_341 br_0_341 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c341
+ bl_0_341 br_0_341 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c341
+ bl_0_341 br_0_341 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c341
+ bl_0_341 br_0_341 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c341
+ bl_0_341 br_0_341 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c341
+ bl_0_341 br_0_341 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c341
+ bl_0_341 br_0_341 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c341
+ bl_0_341 br_0_341 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c341
+ bl_0_341 br_0_341 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c341
+ bl_0_341 br_0_341 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c341
+ bl_0_341 br_0_341 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c341
+ bl_0_341 br_0_341 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c341
+ bl_0_341 br_0_341 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c341
+ bl_0_341 br_0_341 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c341
+ bl_0_341 br_0_341 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c341
+ bl_0_341 br_0_341 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c341
+ bl_0_341 br_0_341 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c341
+ bl_0_341 br_0_341 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c341
+ bl_0_341 br_0_341 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c341
+ bl_0_341 br_0_341 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c341
+ bl_0_341 br_0_341 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c341
+ bl_0_341 br_0_341 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c341
+ bl_0_341 br_0_341 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c341
+ bl_0_341 br_0_341 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c341
+ bl_0_341 br_0_341 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c341
+ bl_0_341 br_0_341 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c341
+ bl_0_341 br_0_341 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c341
+ bl_0_341 br_0_341 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c341
+ bl_0_341 br_0_341 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c341
+ bl_0_341 br_0_341 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c341
+ bl_0_341 br_0_341 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c341
+ bl_0_341 br_0_341 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c341
+ bl_0_341 br_0_341 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c341
+ bl_0_341 br_0_341 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c341
+ bl_0_341 br_0_341 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c341
+ bl_0_341 br_0_341 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c341
+ bl_0_341 br_0_341 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c341
+ bl_0_341 br_0_341 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c341
+ bl_0_341 br_0_341 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c342
+ bl_0_342 br_0_342 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c342
+ bl_0_342 br_0_342 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c342
+ bl_0_342 br_0_342 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c342
+ bl_0_342 br_0_342 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c342
+ bl_0_342 br_0_342 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c342
+ bl_0_342 br_0_342 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c342
+ bl_0_342 br_0_342 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c342
+ bl_0_342 br_0_342 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c342
+ bl_0_342 br_0_342 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c342
+ bl_0_342 br_0_342 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c342
+ bl_0_342 br_0_342 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c342
+ bl_0_342 br_0_342 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c342
+ bl_0_342 br_0_342 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c342
+ bl_0_342 br_0_342 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c342
+ bl_0_342 br_0_342 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c342
+ bl_0_342 br_0_342 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c342
+ bl_0_342 br_0_342 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c342
+ bl_0_342 br_0_342 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c342
+ bl_0_342 br_0_342 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c342
+ bl_0_342 br_0_342 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c342
+ bl_0_342 br_0_342 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c342
+ bl_0_342 br_0_342 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c342
+ bl_0_342 br_0_342 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c342
+ bl_0_342 br_0_342 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c342
+ bl_0_342 br_0_342 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c342
+ bl_0_342 br_0_342 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c342
+ bl_0_342 br_0_342 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c342
+ bl_0_342 br_0_342 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c342
+ bl_0_342 br_0_342 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c342
+ bl_0_342 br_0_342 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c342
+ bl_0_342 br_0_342 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c342
+ bl_0_342 br_0_342 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c342
+ bl_0_342 br_0_342 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c342
+ bl_0_342 br_0_342 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c342
+ bl_0_342 br_0_342 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c342
+ bl_0_342 br_0_342 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c342
+ bl_0_342 br_0_342 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c342
+ bl_0_342 br_0_342 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c342
+ bl_0_342 br_0_342 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c342
+ bl_0_342 br_0_342 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c342
+ bl_0_342 br_0_342 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c342
+ bl_0_342 br_0_342 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c342
+ bl_0_342 br_0_342 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c342
+ bl_0_342 br_0_342 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c342
+ bl_0_342 br_0_342 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c343
+ bl_0_343 br_0_343 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c343
+ bl_0_343 br_0_343 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c343
+ bl_0_343 br_0_343 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c343
+ bl_0_343 br_0_343 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c343
+ bl_0_343 br_0_343 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c343
+ bl_0_343 br_0_343 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c343
+ bl_0_343 br_0_343 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c343
+ bl_0_343 br_0_343 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c343
+ bl_0_343 br_0_343 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c343
+ bl_0_343 br_0_343 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c343
+ bl_0_343 br_0_343 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c343
+ bl_0_343 br_0_343 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c343
+ bl_0_343 br_0_343 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c343
+ bl_0_343 br_0_343 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c343
+ bl_0_343 br_0_343 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c343
+ bl_0_343 br_0_343 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c343
+ bl_0_343 br_0_343 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c343
+ bl_0_343 br_0_343 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c343
+ bl_0_343 br_0_343 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c343
+ bl_0_343 br_0_343 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c343
+ bl_0_343 br_0_343 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c343
+ bl_0_343 br_0_343 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c343
+ bl_0_343 br_0_343 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c343
+ bl_0_343 br_0_343 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c343
+ bl_0_343 br_0_343 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c343
+ bl_0_343 br_0_343 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c343
+ bl_0_343 br_0_343 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c343
+ bl_0_343 br_0_343 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c343
+ bl_0_343 br_0_343 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c343
+ bl_0_343 br_0_343 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c343
+ bl_0_343 br_0_343 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c343
+ bl_0_343 br_0_343 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c343
+ bl_0_343 br_0_343 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c343
+ bl_0_343 br_0_343 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c343
+ bl_0_343 br_0_343 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c343
+ bl_0_343 br_0_343 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c343
+ bl_0_343 br_0_343 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c343
+ bl_0_343 br_0_343 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c343
+ bl_0_343 br_0_343 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c343
+ bl_0_343 br_0_343 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c343
+ bl_0_343 br_0_343 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c343
+ bl_0_343 br_0_343 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c343
+ bl_0_343 br_0_343 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c343
+ bl_0_343 br_0_343 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c343
+ bl_0_343 br_0_343 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c344
+ bl_0_344 br_0_344 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c344
+ bl_0_344 br_0_344 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c344
+ bl_0_344 br_0_344 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c344
+ bl_0_344 br_0_344 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c344
+ bl_0_344 br_0_344 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c344
+ bl_0_344 br_0_344 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c344
+ bl_0_344 br_0_344 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c344
+ bl_0_344 br_0_344 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c344
+ bl_0_344 br_0_344 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c344
+ bl_0_344 br_0_344 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c344
+ bl_0_344 br_0_344 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c344
+ bl_0_344 br_0_344 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c344
+ bl_0_344 br_0_344 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c344
+ bl_0_344 br_0_344 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c344
+ bl_0_344 br_0_344 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c344
+ bl_0_344 br_0_344 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c344
+ bl_0_344 br_0_344 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c344
+ bl_0_344 br_0_344 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c344
+ bl_0_344 br_0_344 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c344
+ bl_0_344 br_0_344 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c344
+ bl_0_344 br_0_344 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c344
+ bl_0_344 br_0_344 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c344
+ bl_0_344 br_0_344 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c344
+ bl_0_344 br_0_344 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c344
+ bl_0_344 br_0_344 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c344
+ bl_0_344 br_0_344 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c344
+ bl_0_344 br_0_344 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c344
+ bl_0_344 br_0_344 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c344
+ bl_0_344 br_0_344 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c344
+ bl_0_344 br_0_344 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c344
+ bl_0_344 br_0_344 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c344
+ bl_0_344 br_0_344 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c344
+ bl_0_344 br_0_344 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c344
+ bl_0_344 br_0_344 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c344
+ bl_0_344 br_0_344 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c344
+ bl_0_344 br_0_344 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c344
+ bl_0_344 br_0_344 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c344
+ bl_0_344 br_0_344 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c344
+ bl_0_344 br_0_344 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c344
+ bl_0_344 br_0_344 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c344
+ bl_0_344 br_0_344 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c344
+ bl_0_344 br_0_344 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c344
+ bl_0_344 br_0_344 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c344
+ bl_0_344 br_0_344 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c344
+ bl_0_344 br_0_344 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c345
+ bl_0_345 br_0_345 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c345
+ bl_0_345 br_0_345 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c345
+ bl_0_345 br_0_345 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c345
+ bl_0_345 br_0_345 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c345
+ bl_0_345 br_0_345 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c345
+ bl_0_345 br_0_345 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c345
+ bl_0_345 br_0_345 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c345
+ bl_0_345 br_0_345 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c345
+ bl_0_345 br_0_345 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c345
+ bl_0_345 br_0_345 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c345
+ bl_0_345 br_0_345 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c345
+ bl_0_345 br_0_345 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c345
+ bl_0_345 br_0_345 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c345
+ bl_0_345 br_0_345 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c345
+ bl_0_345 br_0_345 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c345
+ bl_0_345 br_0_345 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c345
+ bl_0_345 br_0_345 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c345
+ bl_0_345 br_0_345 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c345
+ bl_0_345 br_0_345 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c345
+ bl_0_345 br_0_345 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c345
+ bl_0_345 br_0_345 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c345
+ bl_0_345 br_0_345 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c345
+ bl_0_345 br_0_345 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c345
+ bl_0_345 br_0_345 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c345
+ bl_0_345 br_0_345 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c345
+ bl_0_345 br_0_345 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c345
+ bl_0_345 br_0_345 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c345
+ bl_0_345 br_0_345 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c345
+ bl_0_345 br_0_345 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c345
+ bl_0_345 br_0_345 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c345
+ bl_0_345 br_0_345 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c345
+ bl_0_345 br_0_345 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c345
+ bl_0_345 br_0_345 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c345
+ bl_0_345 br_0_345 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c345
+ bl_0_345 br_0_345 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c345
+ bl_0_345 br_0_345 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c345
+ bl_0_345 br_0_345 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c345
+ bl_0_345 br_0_345 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c345
+ bl_0_345 br_0_345 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c345
+ bl_0_345 br_0_345 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c345
+ bl_0_345 br_0_345 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c345
+ bl_0_345 br_0_345 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c345
+ bl_0_345 br_0_345 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c345
+ bl_0_345 br_0_345 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c345
+ bl_0_345 br_0_345 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c346
+ bl_0_346 br_0_346 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c346
+ bl_0_346 br_0_346 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c346
+ bl_0_346 br_0_346 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c346
+ bl_0_346 br_0_346 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c346
+ bl_0_346 br_0_346 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c346
+ bl_0_346 br_0_346 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c346
+ bl_0_346 br_0_346 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c346
+ bl_0_346 br_0_346 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c346
+ bl_0_346 br_0_346 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c346
+ bl_0_346 br_0_346 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c346
+ bl_0_346 br_0_346 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c346
+ bl_0_346 br_0_346 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c346
+ bl_0_346 br_0_346 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c346
+ bl_0_346 br_0_346 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c346
+ bl_0_346 br_0_346 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c346
+ bl_0_346 br_0_346 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c346
+ bl_0_346 br_0_346 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c346
+ bl_0_346 br_0_346 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c346
+ bl_0_346 br_0_346 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c346
+ bl_0_346 br_0_346 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c346
+ bl_0_346 br_0_346 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c346
+ bl_0_346 br_0_346 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c346
+ bl_0_346 br_0_346 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c346
+ bl_0_346 br_0_346 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c346
+ bl_0_346 br_0_346 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c346
+ bl_0_346 br_0_346 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c346
+ bl_0_346 br_0_346 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c346
+ bl_0_346 br_0_346 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c346
+ bl_0_346 br_0_346 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c346
+ bl_0_346 br_0_346 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c346
+ bl_0_346 br_0_346 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c346
+ bl_0_346 br_0_346 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c346
+ bl_0_346 br_0_346 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c346
+ bl_0_346 br_0_346 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c346
+ bl_0_346 br_0_346 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c346
+ bl_0_346 br_0_346 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c346
+ bl_0_346 br_0_346 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c346
+ bl_0_346 br_0_346 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c346
+ bl_0_346 br_0_346 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c346
+ bl_0_346 br_0_346 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c346
+ bl_0_346 br_0_346 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c346
+ bl_0_346 br_0_346 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c346
+ bl_0_346 br_0_346 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c346
+ bl_0_346 br_0_346 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c346
+ bl_0_346 br_0_346 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c347
+ bl_0_347 br_0_347 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c347
+ bl_0_347 br_0_347 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c347
+ bl_0_347 br_0_347 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c347
+ bl_0_347 br_0_347 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c347
+ bl_0_347 br_0_347 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c347
+ bl_0_347 br_0_347 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c347
+ bl_0_347 br_0_347 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c347
+ bl_0_347 br_0_347 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c347
+ bl_0_347 br_0_347 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c347
+ bl_0_347 br_0_347 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c347
+ bl_0_347 br_0_347 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c347
+ bl_0_347 br_0_347 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c347
+ bl_0_347 br_0_347 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c347
+ bl_0_347 br_0_347 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c347
+ bl_0_347 br_0_347 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c347
+ bl_0_347 br_0_347 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c347
+ bl_0_347 br_0_347 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c347
+ bl_0_347 br_0_347 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c347
+ bl_0_347 br_0_347 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c347
+ bl_0_347 br_0_347 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c347
+ bl_0_347 br_0_347 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c347
+ bl_0_347 br_0_347 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c347
+ bl_0_347 br_0_347 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c347
+ bl_0_347 br_0_347 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c347
+ bl_0_347 br_0_347 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c347
+ bl_0_347 br_0_347 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c347
+ bl_0_347 br_0_347 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c347
+ bl_0_347 br_0_347 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c347
+ bl_0_347 br_0_347 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c347
+ bl_0_347 br_0_347 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c347
+ bl_0_347 br_0_347 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c347
+ bl_0_347 br_0_347 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c347
+ bl_0_347 br_0_347 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c347
+ bl_0_347 br_0_347 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c347
+ bl_0_347 br_0_347 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c347
+ bl_0_347 br_0_347 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c347
+ bl_0_347 br_0_347 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c347
+ bl_0_347 br_0_347 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c347
+ bl_0_347 br_0_347 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c347
+ bl_0_347 br_0_347 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c347
+ bl_0_347 br_0_347 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c347
+ bl_0_347 br_0_347 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c347
+ bl_0_347 br_0_347 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c347
+ bl_0_347 br_0_347 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c347
+ bl_0_347 br_0_347 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c348
+ bl_0_348 br_0_348 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c348
+ bl_0_348 br_0_348 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c348
+ bl_0_348 br_0_348 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c348
+ bl_0_348 br_0_348 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c348
+ bl_0_348 br_0_348 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c348
+ bl_0_348 br_0_348 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c348
+ bl_0_348 br_0_348 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c348
+ bl_0_348 br_0_348 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c348
+ bl_0_348 br_0_348 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c348
+ bl_0_348 br_0_348 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c348
+ bl_0_348 br_0_348 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c348
+ bl_0_348 br_0_348 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c348
+ bl_0_348 br_0_348 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c348
+ bl_0_348 br_0_348 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c348
+ bl_0_348 br_0_348 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c348
+ bl_0_348 br_0_348 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c348
+ bl_0_348 br_0_348 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c348
+ bl_0_348 br_0_348 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c348
+ bl_0_348 br_0_348 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c348
+ bl_0_348 br_0_348 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c348
+ bl_0_348 br_0_348 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c348
+ bl_0_348 br_0_348 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c348
+ bl_0_348 br_0_348 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c348
+ bl_0_348 br_0_348 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c348
+ bl_0_348 br_0_348 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c348
+ bl_0_348 br_0_348 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c348
+ bl_0_348 br_0_348 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c348
+ bl_0_348 br_0_348 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c348
+ bl_0_348 br_0_348 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c348
+ bl_0_348 br_0_348 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c348
+ bl_0_348 br_0_348 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c348
+ bl_0_348 br_0_348 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c348
+ bl_0_348 br_0_348 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c348
+ bl_0_348 br_0_348 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c348
+ bl_0_348 br_0_348 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c348
+ bl_0_348 br_0_348 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c348
+ bl_0_348 br_0_348 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c348
+ bl_0_348 br_0_348 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c348
+ bl_0_348 br_0_348 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c348
+ bl_0_348 br_0_348 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c348
+ bl_0_348 br_0_348 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c348
+ bl_0_348 br_0_348 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c348
+ bl_0_348 br_0_348 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c348
+ bl_0_348 br_0_348 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c348
+ bl_0_348 br_0_348 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c349
+ bl_0_349 br_0_349 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c349
+ bl_0_349 br_0_349 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c349
+ bl_0_349 br_0_349 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c349
+ bl_0_349 br_0_349 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c349
+ bl_0_349 br_0_349 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c349
+ bl_0_349 br_0_349 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c349
+ bl_0_349 br_0_349 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c349
+ bl_0_349 br_0_349 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c349
+ bl_0_349 br_0_349 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c349
+ bl_0_349 br_0_349 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c349
+ bl_0_349 br_0_349 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c349
+ bl_0_349 br_0_349 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c349
+ bl_0_349 br_0_349 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c349
+ bl_0_349 br_0_349 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c349
+ bl_0_349 br_0_349 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c349
+ bl_0_349 br_0_349 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c349
+ bl_0_349 br_0_349 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c349
+ bl_0_349 br_0_349 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c349
+ bl_0_349 br_0_349 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c349
+ bl_0_349 br_0_349 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c349
+ bl_0_349 br_0_349 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c349
+ bl_0_349 br_0_349 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c349
+ bl_0_349 br_0_349 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c349
+ bl_0_349 br_0_349 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c349
+ bl_0_349 br_0_349 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c349
+ bl_0_349 br_0_349 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c349
+ bl_0_349 br_0_349 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c349
+ bl_0_349 br_0_349 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c349
+ bl_0_349 br_0_349 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c349
+ bl_0_349 br_0_349 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c349
+ bl_0_349 br_0_349 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c349
+ bl_0_349 br_0_349 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c349
+ bl_0_349 br_0_349 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c349
+ bl_0_349 br_0_349 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c349
+ bl_0_349 br_0_349 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c349
+ bl_0_349 br_0_349 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c349
+ bl_0_349 br_0_349 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c349
+ bl_0_349 br_0_349 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c349
+ bl_0_349 br_0_349 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c349
+ bl_0_349 br_0_349 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c349
+ bl_0_349 br_0_349 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c349
+ bl_0_349 br_0_349 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c349
+ bl_0_349 br_0_349 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c349
+ bl_0_349 br_0_349 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c349
+ bl_0_349 br_0_349 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c350
+ bl_0_350 br_0_350 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c350
+ bl_0_350 br_0_350 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c350
+ bl_0_350 br_0_350 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c350
+ bl_0_350 br_0_350 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c350
+ bl_0_350 br_0_350 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c350
+ bl_0_350 br_0_350 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c350
+ bl_0_350 br_0_350 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c350
+ bl_0_350 br_0_350 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c350
+ bl_0_350 br_0_350 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c350
+ bl_0_350 br_0_350 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c350
+ bl_0_350 br_0_350 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c350
+ bl_0_350 br_0_350 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c350
+ bl_0_350 br_0_350 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c350
+ bl_0_350 br_0_350 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c350
+ bl_0_350 br_0_350 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c350
+ bl_0_350 br_0_350 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c350
+ bl_0_350 br_0_350 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c350
+ bl_0_350 br_0_350 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c350
+ bl_0_350 br_0_350 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c350
+ bl_0_350 br_0_350 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c350
+ bl_0_350 br_0_350 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c350
+ bl_0_350 br_0_350 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c350
+ bl_0_350 br_0_350 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c350
+ bl_0_350 br_0_350 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c350
+ bl_0_350 br_0_350 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c350
+ bl_0_350 br_0_350 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c350
+ bl_0_350 br_0_350 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c350
+ bl_0_350 br_0_350 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c350
+ bl_0_350 br_0_350 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c350
+ bl_0_350 br_0_350 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c350
+ bl_0_350 br_0_350 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c350
+ bl_0_350 br_0_350 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c350
+ bl_0_350 br_0_350 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c350
+ bl_0_350 br_0_350 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c350
+ bl_0_350 br_0_350 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c350
+ bl_0_350 br_0_350 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c350
+ bl_0_350 br_0_350 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c350
+ bl_0_350 br_0_350 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c350
+ bl_0_350 br_0_350 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c350
+ bl_0_350 br_0_350 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c350
+ bl_0_350 br_0_350 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c350
+ bl_0_350 br_0_350 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c350
+ bl_0_350 br_0_350 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c350
+ bl_0_350 br_0_350 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c350
+ bl_0_350 br_0_350 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c351
+ bl_0_351 br_0_351 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c351
+ bl_0_351 br_0_351 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c351
+ bl_0_351 br_0_351 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c351
+ bl_0_351 br_0_351 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c351
+ bl_0_351 br_0_351 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c351
+ bl_0_351 br_0_351 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c351
+ bl_0_351 br_0_351 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c351
+ bl_0_351 br_0_351 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c351
+ bl_0_351 br_0_351 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c351
+ bl_0_351 br_0_351 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c351
+ bl_0_351 br_0_351 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c351
+ bl_0_351 br_0_351 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c351
+ bl_0_351 br_0_351 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c351
+ bl_0_351 br_0_351 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c351
+ bl_0_351 br_0_351 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c351
+ bl_0_351 br_0_351 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c351
+ bl_0_351 br_0_351 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c351
+ bl_0_351 br_0_351 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c351
+ bl_0_351 br_0_351 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c351
+ bl_0_351 br_0_351 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c351
+ bl_0_351 br_0_351 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c351
+ bl_0_351 br_0_351 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c351
+ bl_0_351 br_0_351 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c351
+ bl_0_351 br_0_351 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c351
+ bl_0_351 br_0_351 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c351
+ bl_0_351 br_0_351 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c351
+ bl_0_351 br_0_351 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c351
+ bl_0_351 br_0_351 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c351
+ bl_0_351 br_0_351 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c351
+ bl_0_351 br_0_351 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c351
+ bl_0_351 br_0_351 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c351
+ bl_0_351 br_0_351 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c351
+ bl_0_351 br_0_351 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c351
+ bl_0_351 br_0_351 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c351
+ bl_0_351 br_0_351 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c351
+ bl_0_351 br_0_351 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c351
+ bl_0_351 br_0_351 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c351
+ bl_0_351 br_0_351 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c351
+ bl_0_351 br_0_351 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c351
+ bl_0_351 br_0_351 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c351
+ bl_0_351 br_0_351 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c351
+ bl_0_351 br_0_351 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c351
+ bl_0_351 br_0_351 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c351
+ bl_0_351 br_0_351 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c351
+ bl_0_351 br_0_351 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c352
+ bl_0_352 br_0_352 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c352
+ bl_0_352 br_0_352 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c352
+ bl_0_352 br_0_352 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c352
+ bl_0_352 br_0_352 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c352
+ bl_0_352 br_0_352 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c352
+ bl_0_352 br_0_352 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c352
+ bl_0_352 br_0_352 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c352
+ bl_0_352 br_0_352 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c352
+ bl_0_352 br_0_352 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c352
+ bl_0_352 br_0_352 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c352
+ bl_0_352 br_0_352 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c352
+ bl_0_352 br_0_352 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c352
+ bl_0_352 br_0_352 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c352
+ bl_0_352 br_0_352 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c352
+ bl_0_352 br_0_352 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c352
+ bl_0_352 br_0_352 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c352
+ bl_0_352 br_0_352 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c352
+ bl_0_352 br_0_352 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c352
+ bl_0_352 br_0_352 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c352
+ bl_0_352 br_0_352 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c352
+ bl_0_352 br_0_352 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c352
+ bl_0_352 br_0_352 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c352
+ bl_0_352 br_0_352 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c352
+ bl_0_352 br_0_352 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c352
+ bl_0_352 br_0_352 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c352
+ bl_0_352 br_0_352 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c352
+ bl_0_352 br_0_352 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c352
+ bl_0_352 br_0_352 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c352
+ bl_0_352 br_0_352 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c352
+ bl_0_352 br_0_352 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c352
+ bl_0_352 br_0_352 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c352
+ bl_0_352 br_0_352 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c352
+ bl_0_352 br_0_352 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c352
+ bl_0_352 br_0_352 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c352
+ bl_0_352 br_0_352 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c352
+ bl_0_352 br_0_352 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c352
+ bl_0_352 br_0_352 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c352
+ bl_0_352 br_0_352 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c352
+ bl_0_352 br_0_352 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c352
+ bl_0_352 br_0_352 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c352
+ bl_0_352 br_0_352 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c352
+ bl_0_352 br_0_352 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c352
+ bl_0_352 br_0_352 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c352
+ bl_0_352 br_0_352 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c352
+ bl_0_352 br_0_352 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c353
+ bl_0_353 br_0_353 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c353
+ bl_0_353 br_0_353 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c353
+ bl_0_353 br_0_353 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c353
+ bl_0_353 br_0_353 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c353
+ bl_0_353 br_0_353 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c353
+ bl_0_353 br_0_353 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c353
+ bl_0_353 br_0_353 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c353
+ bl_0_353 br_0_353 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c353
+ bl_0_353 br_0_353 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c353
+ bl_0_353 br_0_353 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c353
+ bl_0_353 br_0_353 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c353
+ bl_0_353 br_0_353 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c353
+ bl_0_353 br_0_353 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c353
+ bl_0_353 br_0_353 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c353
+ bl_0_353 br_0_353 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c353
+ bl_0_353 br_0_353 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c353
+ bl_0_353 br_0_353 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c353
+ bl_0_353 br_0_353 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c353
+ bl_0_353 br_0_353 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c353
+ bl_0_353 br_0_353 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c353
+ bl_0_353 br_0_353 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c353
+ bl_0_353 br_0_353 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c353
+ bl_0_353 br_0_353 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c353
+ bl_0_353 br_0_353 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c353
+ bl_0_353 br_0_353 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c353
+ bl_0_353 br_0_353 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c353
+ bl_0_353 br_0_353 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c353
+ bl_0_353 br_0_353 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c353
+ bl_0_353 br_0_353 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c353
+ bl_0_353 br_0_353 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c353
+ bl_0_353 br_0_353 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c353
+ bl_0_353 br_0_353 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c353
+ bl_0_353 br_0_353 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c353
+ bl_0_353 br_0_353 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c353
+ bl_0_353 br_0_353 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c353
+ bl_0_353 br_0_353 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c353
+ bl_0_353 br_0_353 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c353
+ bl_0_353 br_0_353 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c353
+ bl_0_353 br_0_353 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c353
+ bl_0_353 br_0_353 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c353
+ bl_0_353 br_0_353 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c353
+ bl_0_353 br_0_353 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c353
+ bl_0_353 br_0_353 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c353
+ bl_0_353 br_0_353 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c353
+ bl_0_353 br_0_353 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c354
+ bl_0_354 br_0_354 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c354
+ bl_0_354 br_0_354 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c354
+ bl_0_354 br_0_354 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c354
+ bl_0_354 br_0_354 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c354
+ bl_0_354 br_0_354 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c354
+ bl_0_354 br_0_354 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c354
+ bl_0_354 br_0_354 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c354
+ bl_0_354 br_0_354 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c354
+ bl_0_354 br_0_354 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c354
+ bl_0_354 br_0_354 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c354
+ bl_0_354 br_0_354 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c354
+ bl_0_354 br_0_354 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c354
+ bl_0_354 br_0_354 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c354
+ bl_0_354 br_0_354 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c354
+ bl_0_354 br_0_354 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c354
+ bl_0_354 br_0_354 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c354
+ bl_0_354 br_0_354 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c354
+ bl_0_354 br_0_354 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c354
+ bl_0_354 br_0_354 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c354
+ bl_0_354 br_0_354 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c354
+ bl_0_354 br_0_354 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c354
+ bl_0_354 br_0_354 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c354
+ bl_0_354 br_0_354 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c354
+ bl_0_354 br_0_354 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c354
+ bl_0_354 br_0_354 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c354
+ bl_0_354 br_0_354 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c354
+ bl_0_354 br_0_354 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c354
+ bl_0_354 br_0_354 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c354
+ bl_0_354 br_0_354 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c354
+ bl_0_354 br_0_354 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c354
+ bl_0_354 br_0_354 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c354
+ bl_0_354 br_0_354 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c354
+ bl_0_354 br_0_354 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c354
+ bl_0_354 br_0_354 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c354
+ bl_0_354 br_0_354 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c354
+ bl_0_354 br_0_354 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c354
+ bl_0_354 br_0_354 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c354
+ bl_0_354 br_0_354 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c354
+ bl_0_354 br_0_354 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c354
+ bl_0_354 br_0_354 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c354
+ bl_0_354 br_0_354 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c354
+ bl_0_354 br_0_354 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c354
+ bl_0_354 br_0_354 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c354
+ bl_0_354 br_0_354 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c354
+ bl_0_354 br_0_354 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c355
+ bl_0_355 br_0_355 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c355
+ bl_0_355 br_0_355 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c355
+ bl_0_355 br_0_355 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c355
+ bl_0_355 br_0_355 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c355
+ bl_0_355 br_0_355 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c355
+ bl_0_355 br_0_355 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c355
+ bl_0_355 br_0_355 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c355
+ bl_0_355 br_0_355 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c355
+ bl_0_355 br_0_355 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c355
+ bl_0_355 br_0_355 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c355
+ bl_0_355 br_0_355 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c355
+ bl_0_355 br_0_355 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c355
+ bl_0_355 br_0_355 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c355
+ bl_0_355 br_0_355 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c355
+ bl_0_355 br_0_355 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c355
+ bl_0_355 br_0_355 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c355
+ bl_0_355 br_0_355 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c355
+ bl_0_355 br_0_355 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c355
+ bl_0_355 br_0_355 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c355
+ bl_0_355 br_0_355 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c355
+ bl_0_355 br_0_355 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c355
+ bl_0_355 br_0_355 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c355
+ bl_0_355 br_0_355 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c355
+ bl_0_355 br_0_355 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c355
+ bl_0_355 br_0_355 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c355
+ bl_0_355 br_0_355 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c355
+ bl_0_355 br_0_355 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c355
+ bl_0_355 br_0_355 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c355
+ bl_0_355 br_0_355 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c355
+ bl_0_355 br_0_355 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c355
+ bl_0_355 br_0_355 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c355
+ bl_0_355 br_0_355 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c355
+ bl_0_355 br_0_355 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c355
+ bl_0_355 br_0_355 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c355
+ bl_0_355 br_0_355 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c355
+ bl_0_355 br_0_355 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c355
+ bl_0_355 br_0_355 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c355
+ bl_0_355 br_0_355 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c355
+ bl_0_355 br_0_355 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c355
+ bl_0_355 br_0_355 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c355
+ bl_0_355 br_0_355 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c355
+ bl_0_355 br_0_355 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c355
+ bl_0_355 br_0_355 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c355
+ bl_0_355 br_0_355 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c355
+ bl_0_355 br_0_355 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c356
+ bl_0_356 br_0_356 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c356
+ bl_0_356 br_0_356 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c356
+ bl_0_356 br_0_356 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c356
+ bl_0_356 br_0_356 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c356
+ bl_0_356 br_0_356 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c356
+ bl_0_356 br_0_356 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c356
+ bl_0_356 br_0_356 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c356
+ bl_0_356 br_0_356 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c356
+ bl_0_356 br_0_356 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c356
+ bl_0_356 br_0_356 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c356
+ bl_0_356 br_0_356 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c356
+ bl_0_356 br_0_356 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c356
+ bl_0_356 br_0_356 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c356
+ bl_0_356 br_0_356 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c356
+ bl_0_356 br_0_356 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c356
+ bl_0_356 br_0_356 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c356
+ bl_0_356 br_0_356 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c356
+ bl_0_356 br_0_356 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c356
+ bl_0_356 br_0_356 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c356
+ bl_0_356 br_0_356 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c356
+ bl_0_356 br_0_356 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c356
+ bl_0_356 br_0_356 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c356
+ bl_0_356 br_0_356 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c356
+ bl_0_356 br_0_356 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c356
+ bl_0_356 br_0_356 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c356
+ bl_0_356 br_0_356 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c356
+ bl_0_356 br_0_356 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c356
+ bl_0_356 br_0_356 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c356
+ bl_0_356 br_0_356 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c356
+ bl_0_356 br_0_356 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c356
+ bl_0_356 br_0_356 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c356
+ bl_0_356 br_0_356 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c356
+ bl_0_356 br_0_356 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c356
+ bl_0_356 br_0_356 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c356
+ bl_0_356 br_0_356 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c356
+ bl_0_356 br_0_356 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c356
+ bl_0_356 br_0_356 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c356
+ bl_0_356 br_0_356 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c356
+ bl_0_356 br_0_356 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c356
+ bl_0_356 br_0_356 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c356
+ bl_0_356 br_0_356 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c356
+ bl_0_356 br_0_356 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c356
+ bl_0_356 br_0_356 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c356
+ bl_0_356 br_0_356 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c356
+ bl_0_356 br_0_356 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c357
+ bl_0_357 br_0_357 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c357
+ bl_0_357 br_0_357 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c357
+ bl_0_357 br_0_357 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c357
+ bl_0_357 br_0_357 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c357
+ bl_0_357 br_0_357 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c357
+ bl_0_357 br_0_357 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c357
+ bl_0_357 br_0_357 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c357
+ bl_0_357 br_0_357 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c357
+ bl_0_357 br_0_357 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c357
+ bl_0_357 br_0_357 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c357
+ bl_0_357 br_0_357 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c357
+ bl_0_357 br_0_357 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c357
+ bl_0_357 br_0_357 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c357
+ bl_0_357 br_0_357 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c357
+ bl_0_357 br_0_357 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c357
+ bl_0_357 br_0_357 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c357
+ bl_0_357 br_0_357 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c357
+ bl_0_357 br_0_357 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c357
+ bl_0_357 br_0_357 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c357
+ bl_0_357 br_0_357 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c357
+ bl_0_357 br_0_357 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c357
+ bl_0_357 br_0_357 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c357
+ bl_0_357 br_0_357 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c357
+ bl_0_357 br_0_357 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c357
+ bl_0_357 br_0_357 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c357
+ bl_0_357 br_0_357 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c357
+ bl_0_357 br_0_357 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c357
+ bl_0_357 br_0_357 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c357
+ bl_0_357 br_0_357 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c357
+ bl_0_357 br_0_357 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c357
+ bl_0_357 br_0_357 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c357
+ bl_0_357 br_0_357 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c357
+ bl_0_357 br_0_357 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c357
+ bl_0_357 br_0_357 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c357
+ bl_0_357 br_0_357 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c357
+ bl_0_357 br_0_357 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c357
+ bl_0_357 br_0_357 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c357
+ bl_0_357 br_0_357 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c357
+ bl_0_357 br_0_357 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c357
+ bl_0_357 br_0_357 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c357
+ bl_0_357 br_0_357 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c357
+ bl_0_357 br_0_357 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c357
+ bl_0_357 br_0_357 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c357
+ bl_0_357 br_0_357 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c357
+ bl_0_357 br_0_357 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c358
+ bl_0_358 br_0_358 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c358
+ bl_0_358 br_0_358 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c358
+ bl_0_358 br_0_358 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c358
+ bl_0_358 br_0_358 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c358
+ bl_0_358 br_0_358 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c358
+ bl_0_358 br_0_358 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c358
+ bl_0_358 br_0_358 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c358
+ bl_0_358 br_0_358 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c358
+ bl_0_358 br_0_358 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c358
+ bl_0_358 br_0_358 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c358
+ bl_0_358 br_0_358 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c358
+ bl_0_358 br_0_358 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c358
+ bl_0_358 br_0_358 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c358
+ bl_0_358 br_0_358 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c358
+ bl_0_358 br_0_358 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c358
+ bl_0_358 br_0_358 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c358
+ bl_0_358 br_0_358 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c358
+ bl_0_358 br_0_358 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c358
+ bl_0_358 br_0_358 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c358
+ bl_0_358 br_0_358 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c358
+ bl_0_358 br_0_358 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c358
+ bl_0_358 br_0_358 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c358
+ bl_0_358 br_0_358 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c358
+ bl_0_358 br_0_358 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c358
+ bl_0_358 br_0_358 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c358
+ bl_0_358 br_0_358 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c358
+ bl_0_358 br_0_358 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c358
+ bl_0_358 br_0_358 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c358
+ bl_0_358 br_0_358 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c358
+ bl_0_358 br_0_358 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c358
+ bl_0_358 br_0_358 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c358
+ bl_0_358 br_0_358 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c358
+ bl_0_358 br_0_358 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c358
+ bl_0_358 br_0_358 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c358
+ bl_0_358 br_0_358 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c358
+ bl_0_358 br_0_358 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c358
+ bl_0_358 br_0_358 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c358
+ bl_0_358 br_0_358 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c358
+ bl_0_358 br_0_358 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c358
+ bl_0_358 br_0_358 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c358
+ bl_0_358 br_0_358 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c358
+ bl_0_358 br_0_358 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c358
+ bl_0_358 br_0_358 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c358
+ bl_0_358 br_0_358 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c358
+ bl_0_358 br_0_358 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c359
+ bl_0_359 br_0_359 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c359
+ bl_0_359 br_0_359 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c359
+ bl_0_359 br_0_359 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c359
+ bl_0_359 br_0_359 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c359
+ bl_0_359 br_0_359 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c359
+ bl_0_359 br_0_359 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c359
+ bl_0_359 br_0_359 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c359
+ bl_0_359 br_0_359 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c359
+ bl_0_359 br_0_359 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c359
+ bl_0_359 br_0_359 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c359
+ bl_0_359 br_0_359 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c359
+ bl_0_359 br_0_359 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c359
+ bl_0_359 br_0_359 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c359
+ bl_0_359 br_0_359 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c359
+ bl_0_359 br_0_359 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c359
+ bl_0_359 br_0_359 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c359
+ bl_0_359 br_0_359 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c359
+ bl_0_359 br_0_359 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c359
+ bl_0_359 br_0_359 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c359
+ bl_0_359 br_0_359 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c359
+ bl_0_359 br_0_359 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c359
+ bl_0_359 br_0_359 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c359
+ bl_0_359 br_0_359 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c359
+ bl_0_359 br_0_359 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c359
+ bl_0_359 br_0_359 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c359
+ bl_0_359 br_0_359 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c359
+ bl_0_359 br_0_359 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c359
+ bl_0_359 br_0_359 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c359
+ bl_0_359 br_0_359 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c359
+ bl_0_359 br_0_359 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c359
+ bl_0_359 br_0_359 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c359
+ bl_0_359 br_0_359 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c359
+ bl_0_359 br_0_359 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c359
+ bl_0_359 br_0_359 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c359
+ bl_0_359 br_0_359 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c359
+ bl_0_359 br_0_359 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c359
+ bl_0_359 br_0_359 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c359
+ bl_0_359 br_0_359 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c359
+ bl_0_359 br_0_359 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c359
+ bl_0_359 br_0_359 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c359
+ bl_0_359 br_0_359 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c359
+ bl_0_359 br_0_359 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c359
+ bl_0_359 br_0_359 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c359
+ bl_0_359 br_0_359 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c359
+ bl_0_359 br_0_359 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c360
+ bl_0_360 br_0_360 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c360
+ bl_0_360 br_0_360 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c360
+ bl_0_360 br_0_360 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c360
+ bl_0_360 br_0_360 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c360
+ bl_0_360 br_0_360 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c360
+ bl_0_360 br_0_360 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c360
+ bl_0_360 br_0_360 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c360
+ bl_0_360 br_0_360 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c360
+ bl_0_360 br_0_360 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c360
+ bl_0_360 br_0_360 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c360
+ bl_0_360 br_0_360 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c360
+ bl_0_360 br_0_360 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c360
+ bl_0_360 br_0_360 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c360
+ bl_0_360 br_0_360 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c360
+ bl_0_360 br_0_360 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c360
+ bl_0_360 br_0_360 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c360
+ bl_0_360 br_0_360 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c360
+ bl_0_360 br_0_360 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c360
+ bl_0_360 br_0_360 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c360
+ bl_0_360 br_0_360 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c360
+ bl_0_360 br_0_360 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c360
+ bl_0_360 br_0_360 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c360
+ bl_0_360 br_0_360 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c360
+ bl_0_360 br_0_360 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c360
+ bl_0_360 br_0_360 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c360
+ bl_0_360 br_0_360 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c360
+ bl_0_360 br_0_360 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c360
+ bl_0_360 br_0_360 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c360
+ bl_0_360 br_0_360 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c360
+ bl_0_360 br_0_360 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c360
+ bl_0_360 br_0_360 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c360
+ bl_0_360 br_0_360 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c360
+ bl_0_360 br_0_360 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c360
+ bl_0_360 br_0_360 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c360
+ bl_0_360 br_0_360 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c360
+ bl_0_360 br_0_360 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c360
+ bl_0_360 br_0_360 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c360
+ bl_0_360 br_0_360 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c360
+ bl_0_360 br_0_360 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c360
+ bl_0_360 br_0_360 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c360
+ bl_0_360 br_0_360 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c360
+ bl_0_360 br_0_360 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c360
+ bl_0_360 br_0_360 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c360
+ bl_0_360 br_0_360 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c360
+ bl_0_360 br_0_360 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c361
+ bl_0_361 br_0_361 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c361
+ bl_0_361 br_0_361 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c361
+ bl_0_361 br_0_361 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c361
+ bl_0_361 br_0_361 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c361
+ bl_0_361 br_0_361 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c361
+ bl_0_361 br_0_361 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c361
+ bl_0_361 br_0_361 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c361
+ bl_0_361 br_0_361 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c361
+ bl_0_361 br_0_361 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c361
+ bl_0_361 br_0_361 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c361
+ bl_0_361 br_0_361 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c361
+ bl_0_361 br_0_361 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c361
+ bl_0_361 br_0_361 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c361
+ bl_0_361 br_0_361 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c361
+ bl_0_361 br_0_361 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c361
+ bl_0_361 br_0_361 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c361
+ bl_0_361 br_0_361 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c361
+ bl_0_361 br_0_361 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c361
+ bl_0_361 br_0_361 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c361
+ bl_0_361 br_0_361 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c361
+ bl_0_361 br_0_361 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c361
+ bl_0_361 br_0_361 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c361
+ bl_0_361 br_0_361 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c361
+ bl_0_361 br_0_361 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c361
+ bl_0_361 br_0_361 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c361
+ bl_0_361 br_0_361 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c361
+ bl_0_361 br_0_361 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c361
+ bl_0_361 br_0_361 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c361
+ bl_0_361 br_0_361 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c361
+ bl_0_361 br_0_361 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c361
+ bl_0_361 br_0_361 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c361
+ bl_0_361 br_0_361 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c361
+ bl_0_361 br_0_361 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c361
+ bl_0_361 br_0_361 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c361
+ bl_0_361 br_0_361 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c361
+ bl_0_361 br_0_361 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c361
+ bl_0_361 br_0_361 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c361
+ bl_0_361 br_0_361 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c361
+ bl_0_361 br_0_361 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c361
+ bl_0_361 br_0_361 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c361
+ bl_0_361 br_0_361 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c361
+ bl_0_361 br_0_361 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c361
+ bl_0_361 br_0_361 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c361
+ bl_0_361 br_0_361 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c361
+ bl_0_361 br_0_361 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c362
+ bl_0_362 br_0_362 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c362
+ bl_0_362 br_0_362 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c362
+ bl_0_362 br_0_362 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c362
+ bl_0_362 br_0_362 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c362
+ bl_0_362 br_0_362 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c362
+ bl_0_362 br_0_362 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c362
+ bl_0_362 br_0_362 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c362
+ bl_0_362 br_0_362 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c362
+ bl_0_362 br_0_362 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c362
+ bl_0_362 br_0_362 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c362
+ bl_0_362 br_0_362 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c362
+ bl_0_362 br_0_362 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c362
+ bl_0_362 br_0_362 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c362
+ bl_0_362 br_0_362 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c362
+ bl_0_362 br_0_362 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c362
+ bl_0_362 br_0_362 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c362
+ bl_0_362 br_0_362 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c362
+ bl_0_362 br_0_362 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c362
+ bl_0_362 br_0_362 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c362
+ bl_0_362 br_0_362 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c362
+ bl_0_362 br_0_362 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c362
+ bl_0_362 br_0_362 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c362
+ bl_0_362 br_0_362 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c362
+ bl_0_362 br_0_362 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c362
+ bl_0_362 br_0_362 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c362
+ bl_0_362 br_0_362 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c362
+ bl_0_362 br_0_362 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c362
+ bl_0_362 br_0_362 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c362
+ bl_0_362 br_0_362 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c362
+ bl_0_362 br_0_362 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c362
+ bl_0_362 br_0_362 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c362
+ bl_0_362 br_0_362 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c362
+ bl_0_362 br_0_362 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c362
+ bl_0_362 br_0_362 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c362
+ bl_0_362 br_0_362 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c362
+ bl_0_362 br_0_362 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c362
+ bl_0_362 br_0_362 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c362
+ bl_0_362 br_0_362 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c362
+ bl_0_362 br_0_362 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c362
+ bl_0_362 br_0_362 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c362
+ bl_0_362 br_0_362 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c362
+ bl_0_362 br_0_362 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c362
+ bl_0_362 br_0_362 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c362
+ bl_0_362 br_0_362 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c362
+ bl_0_362 br_0_362 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c363
+ bl_0_363 br_0_363 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c363
+ bl_0_363 br_0_363 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c363
+ bl_0_363 br_0_363 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c363
+ bl_0_363 br_0_363 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c363
+ bl_0_363 br_0_363 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c363
+ bl_0_363 br_0_363 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c363
+ bl_0_363 br_0_363 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c363
+ bl_0_363 br_0_363 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c363
+ bl_0_363 br_0_363 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c363
+ bl_0_363 br_0_363 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c363
+ bl_0_363 br_0_363 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c363
+ bl_0_363 br_0_363 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c363
+ bl_0_363 br_0_363 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c363
+ bl_0_363 br_0_363 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c363
+ bl_0_363 br_0_363 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c363
+ bl_0_363 br_0_363 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c363
+ bl_0_363 br_0_363 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c363
+ bl_0_363 br_0_363 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c363
+ bl_0_363 br_0_363 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c363
+ bl_0_363 br_0_363 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c363
+ bl_0_363 br_0_363 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c363
+ bl_0_363 br_0_363 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c363
+ bl_0_363 br_0_363 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c363
+ bl_0_363 br_0_363 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c363
+ bl_0_363 br_0_363 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c363
+ bl_0_363 br_0_363 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c363
+ bl_0_363 br_0_363 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c363
+ bl_0_363 br_0_363 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c363
+ bl_0_363 br_0_363 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c363
+ bl_0_363 br_0_363 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c363
+ bl_0_363 br_0_363 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c363
+ bl_0_363 br_0_363 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c363
+ bl_0_363 br_0_363 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c363
+ bl_0_363 br_0_363 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c363
+ bl_0_363 br_0_363 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c363
+ bl_0_363 br_0_363 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c363
+ bl_0_363 br_0_363 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c363
+ bl_0_363 br_0_363 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c363
+ bl_0_363 br_0_363 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c363
+ bl_0_363 br_0_363 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c363
+ bl_0_363 br_0_363 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c363
+ bl_0_363 br_0_363 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c363
+ bl_0_363 br_0_363 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c363
+ bl_0_363 br_0_363 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c363
+ bl_0_363 br_0_363 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c364
+ bl_0_364 br_0_364 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c364
+ bl_0_364 br_0_364 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c364
+ bl_0_364 br_0_364 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c364
+ bl_0_364 br_0_364 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c364
+ bl_0_364 br_0_364 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c364
+ bl_0_364 br_0_364 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c364
+ bl_0_364 br_0_364 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c364
+ bl_0_364 br_0_364 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c364
+ bl_0_364 br_0_364 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c364
+ bl_0_364 br_0_364 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c364
+ bl_0_364 br_0_364 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c364
+ bl_0_364 br_0_364 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c364
+ bl_0_364 br_0_364 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c364
+ bl_0_364 br_0_364 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c364
+ bl_0_364 br_0_364 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c364
+ bl_0_364 br_0_364 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c364
+ bl_0_364 br_0_364 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c364
+ bl_0_364 br_0_364 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c364
+ bl_0_364 br_0_364 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c364
+ bl_0_364 br_0_364 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c364
+ bl_0_364 br_0_364 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c364
+ bl_0_364 br_0_364 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c364
+ bl_0_364 br_0_364 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c364
+ bl_0_364 br_0_364 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c364
+ bl_0_364 br_0_364 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c364
+ bl_0_364 br_0_364 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c364
+ bl_0_364 br_0_364 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c364
+ bl_0_364 br_0_364 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c364
+ bl_0_364 br_0_364 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c364
+ bl_0_364 br_0_364 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c364
+ bl_0_364 br_0_364 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c364
+ bl_0_364 br_0_364 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c364
+ bl_0_364 br_0_364 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c364
+ bl_0_364 br_0_364 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c364
+ bl_0_364 br_0_364 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c364
+ bl_0_364 br_0_364 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c364
+ bl_0_364 br_0_364 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c364
+ bl_0_364 br_0_364 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c364
+ bl_0_364 br_0_364 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c364
+ bl_0_364 br_0_364 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c364
+ bl_0_364 br_0_364 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c364
+ bl_0_364 br_0_364 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c364
+ bl_0_364 br_0_364 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c364
+ bl_0_364 br_0_364 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c364
+ bl_0_364 br_0_364 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c365
+ bl_0_365 br_0_365 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c365
+ bl_0_365 br_0_365 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c365
+ bl_0_365 br_0_365 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c365
+ bl_0_365 br_0_365 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c365
+ bl_0_365 br_0_365 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c365
+ bl_0_365 br_0_365 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c365
+ bl_0_365 br_0_365 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c365
+ bl_0_365 br_0_365 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c365
+ bl_0_365 br_0_365 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c365
+ bl_0_365 br_0_365 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c365
+ bl_0_365 br_0_365 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c365
+ bl_0_365 br_0_365 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c365
+ bl_0_365 br_0_365 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c365
+ bl_0_365 br_0_365 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c365
+ bl_0_365 br_0_365 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c365
+ bl_0_365 br_0_365 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c365
+ bl_0_365 br_0_365 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c365
+ bl_0_365 br_0_365 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c365
+ bl_0_365 br_0_365 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c365
+ bl_0_365 br_0_365 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c365
+ bl_0_365 br_0_365 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c365
+ bl_0_365 br_0_365 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c365
+ bl_0_365 br_0_365 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c365
+ bl_0_365 br_0_365 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c365
+ bl_0_365 br_0_365 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c365
+ bl_0_365 br_0_365 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c365
+ bl_0_365 br_0_365 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c365
+ bl_0_365 br_0_365 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c365
+ bl_0_365 br_0_365 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c365
+ bl_0_365 br_0_365 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c365
+ bl_0_365 br_0_365 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c365
+ bl_0_365 br_0_365 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c365
+ bl_0_365 br_0_365 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c365
+ bl_0_365 br_0_365 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c365
+ bl_0_365 br_0_365 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c365
+ bl_0_365 br_0_365 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c365
+ bl_0_365 br_0_365 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c365
+ bl_0_365 br_0_365 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c365
+ bl_0_365 br_0_365 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c365
+ bl_0_365 br_0_365 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c365
+ bl_0_365 br_0_365 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c365
+ bl_0_365 br_0_365 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c365
+ bl_0_365 br_0_365 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c365
+ bl_0_365 br_0_365 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c365
+ bl_0_365 br_0_365 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c366
+ bl_0_366 br_0_366 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c366
+ bl_0_366 br_0_366 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c366
+ bl_0_366 br_0_366 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c366
+ bl_0_366 br_0_366 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c366
+ bl_0_366 br_0_366 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c366
+ bl_0_366 br_0_366 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c366
+ bl_0_366 br_0_366 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c366
+ bl_0_366 br_0_366 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c366
+ bl_0_366 br_0_366 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c366
+ bl_0_366 br_0_366 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c366
+ bl_0_366 br_0_366 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c366
+ bl_0_366 br_0_366 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c366
+ bl_0_366 br_0_366 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c366
+ bl_0_366 br_0_366 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c366
+ bl_0_366 br_0_366 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c366
+ bl_0_366 br_0_366 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c366
+ bl_0_366 br_0_366 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c366
+ bl_0_366 br_0_366 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c366
+ bl_0_366 br_0_366 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c366
+ bl_0_366 br_0_366 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c366
+ bl_0_366 br_0_366 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c366
+ bl_0_366 br_0_366 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c366
+ bl_0_366 br_0_366 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c366
+ bl_0_366 br_0_366 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c366
+ bl_0_366 br_0_366 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c366
+ bl_0_366 br_0_366 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c366
+ bl_0_366 br_0_366 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c366
+ bl_0_366 br_0_366 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c366
+ bl_0_366 br_0_366 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c366
+ bl_0_366 br_0_366 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c366
+ bl_0_366 br_0_366 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c366
+ bl_0_366 br_0_366 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c366
+ bl_0_366 br_0_366 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c366
+ bl_0_366 br_0_366 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c366
+ bl_0_366 br_0_366 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c366
+ bl_0_366 br_0_366 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c366
+ bl_0_366 br_0_366 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c366
+ bl_0_366 br_0_366 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c366
+ bl_0_366 br_0_366 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c366
+ bl_0_366 br_0_366 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c366
+ bl_0_366 br_0_366 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c366
+ bl_0_366 br_0_366 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c366
+ bl_0_366 br_0_366 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c366
+ bl_0_366 br_0_366 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c366
+ bl_0_366 br_0_366 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c367
+ bl_0_367 br_0_367 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c367
+ bl_0_367 br_0_367 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c367
+ bl_0_367 br_0_367 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c367
+ bl_0_367 br_0_367 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c367
+ bl_0_367 br_0_367 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c367
+ bl_0_367 br_0_367 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c367
+ bl_0_367 br_0_367 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c367
+ bl_0_367 br_0_367 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c367
+ bl_0_367 br_0_367 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c367
+ bl_0_367 br_0_367 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c367
+ bl_0_367 br_0_367 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c367
+ bl_0_367 br_0_367 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c367
+ bl_0_367 br_0_367 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c367
+ bl_0_367 br_0_367 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c367
+ bl_0_367 br_0_367 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c367
+ bl_0_367 br_0_367 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c367
+ bl_0_367 br_0_367 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c367
+ bl_0_367 br_0_367 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c367
+ bl_0_367 br_0_367 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c367
+ bl_0_367 br_0_367 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c367
+ bl_0_367 br_0_367 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c367
+ bl_0_367 br_0_367 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c367
+ bl_0_367 br_0_367 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c367
+ bl_0_367 br_0_367 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c367
+ bl_0_367 br_0_367 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c367
+ bl_0_367 br_0_367 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c367
+ bl_0_367 br_0_367 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c367
+ bl_0_367 br_0_367 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c367
+ bl_0_367 br_0_367 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c367
+ bl_0_367 br_0_367 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c367
+ bl_0_367 br_0_367 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c367
+ bl_0_367 br_0_367 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c367
+ bl_0_367 br_0_367 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c367
+ bl_0_367 br_0_367 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c367
+ bl_0_367 br_0_367 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c367
+ bl_0_367 br_0_367 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c367
+ bl_0_367 br_0_367 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c367
+ bl_0_367 br_0_367 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c367
+ bl_0_367 br_0_367 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c367
+ bl_0_367 br_0_367 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c367
+ bl_0_367 br_0_367 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c367
+ bl_0_367 br_0_367 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c367
+ bl_0_367 br_0_367 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c367
+ bl_0_367 br_0_367 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c367
+ bl_0_367 br_0_367 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c368
+ bl_0_368 br_0_368 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c368
+ bl_0_368 br_0_368 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c368
+ bl_0_368 br_0_368 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c368
+ bl_0_368 br_0_368 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c368
+ bl_0_368 br_0_368 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c368
+ bl_0_368 br_0_368 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c368
+ bl_0_368 br_0_368 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c368
+ bl_0_368 br_0_368 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c368
+ bl_0_368 br_0_368 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c368
+ bl_0_368 br_0_368 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c368
+ bl_0_368 br_0_368 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c368
+ bl_0_368 br_0_368 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c368
+ bl_0_368 br_0_368 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c368
+ bl_0_368 br_0_368 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c368
+ bl_0_368 br_0_368 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c368
+ bl_0_368 br_0_368 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c368
+ bl_0_368 br_0_368 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c368
+ bl_0_368 br_0_368 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c368
+ bl_0_368 br_0_368 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c368
+ bl_0_368 br_0_368 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c368
+ bl_0_368 br_0_368 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c368
+ bl_0_368 br_0_368 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c368
+ bl_0_368 br_0_368 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c368
+ bl_0_368 br_0_368 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c368
+ bl_0_368 br_0_368 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c368
+ bl_0_368 br_0_368 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c368
+ bl_0_368 br_0_368 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c368
+ bl_0_368 br_0_368 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c368
+ bl_0_368 br_0_368 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c368
+ bl_0_368 br_0_368 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c368
+ bl_0_368 br_0_368 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c368
+ bl_0_368 br_0_368 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c368
+ bl_0_368 br_0_368 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c368
+ bl_0_368 br_0_368 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c368
+ bl_0_368 br_0_368 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c368
+ bl_0_368 br_0_368 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c368
+ bl_0_368 br_0_368 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c368
+ bl_0_368 br_0_368 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c368
+ bl_0_368 br_0_368 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c368
+ bl_0_368 br_0_368 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c368
+ bl_0_368 br_0_368 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c368
+ bl_0_368 br_0_368 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c368
+ bl_0_368 br_0_368 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c368
+ bl_0_368 br_0_368 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c368
+ bl_0_368 br_0_368 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c369
+ bl_0_369 br_0_369 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c369
+ bl_0_369 br_0_369 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c369
+ bl_0_369 br_0_369 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c369
+ bl_0_369 br_0_369 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c369
+ bl_0_369 br_0_369 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c369
+ bl_0_369 br_0_369 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c369
+ bl_0_369 br_0_369 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c369
+ bl_0_369 br_0_369 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c369
+ bl_0_369 br_0_369 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c369
+ bl_0_369 br_0_369 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c369
+ bl_0_369 br_0_369 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c369
+ bl_0_369 br_0_369 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c369
+ bl_0_369 br_0_369 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c369
+ bl_0_369 br_0_369 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c369
+ bl_0_369 br_0_369 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c369
+ bl_0_369 br_0_369 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c369
+ bl_0_369 br_0_369 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c369
+ bl_0_369 br_0_369 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c369
+ bl_0_369 br_0_369 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c369
+ bl_0_369 br_0_369 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c369
+ bl_0_369 br_0_369 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c369
+ bl_0_369 br_0_369 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c369
+ bl_0_369 br_0_369 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c369
+ bl_0_369 br_0_369 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c369
+ bl_0_369 br_0_369 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c369
+ bl_0_369 br_0_369 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c369
+ bl_0_369 br_0_369 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c369
+ bl_0_369 br_0_369 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c369
+ bl_0_369 br_0_369 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c369
+ bl_0_369 br_0_369 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c369
+ bl_0_369 br_0_369 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c369
+ bl_0_369 br_0_369 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c369
+ bl_0_369 br_0_369 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c369
+ bl_0_369 br_0_369 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c369
+ bl_0_369 br_0_369 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c369
+ bl_0_369 br_0_369 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c369
+ bl_0_369 br_0_369 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c369
+ bl_0_369 br_0_369 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c369
+ bl_0_369 br_0_369 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c369
+ bl_0_369 br_0_369 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c369
+ bl_0_369 br_0_369 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c369
+ bl_0_369 br_0_369 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c369
+ bl_0_369 br_0_369 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c369
+ bl_0_369 br_0_369 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c369
+ bl_0_369 br_0_369 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c370
+ bl_0_370 br_0_370 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c370
+ bl_0_370 br_0_370 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c370
+ bl_0_370 br_0_370 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c370
+ bl_0_370 br_0_370 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c370
+ bl_0_370 br_0_370 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c370
+ bl_0_370 br_0_370 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c370
+ bl_0_370 br_0_370 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c370
+ bl_0_370 br_0_370 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c370
+ bl_0_370 br_0_370 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c370
+ bl_0_370 br_0_370 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c370
+ bl_0_370 br_0_370 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c370
+ bl_0_370 br_0_370 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c370
+ bl_0_370 br_0_370 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c370
+ bl_0_370 br_0_370 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c370
+ bl_0_370 br_0_370 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c370
+ bl_0_370 br_0_370 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c370
+ bl_0_370 br_0_370 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c370
+ bl_0_370 br_0_370 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c370
+ bl_0_370 br_0_370 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c370
+ bl_0_370 br_0_370 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c370
+ bl_0_370 br_0_370 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c370
+ bl_0_370 br_0_370 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c370
+ bl_0_370 br_0_370 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c370
+ bl_0_370 br_0_370 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c370
+ bl_0_370 br_0_370 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c370
+ bl_0_370 br_0_370 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c370
+ bl_0_370 br_0_370 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c370
+ bl_0_370 br_0_370 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c370
+ bl_0_370 br_0_370 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c370
+ bl_0_370 br_0_370 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c370
+ bl_0_370 br_0_370 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c370
+ bl_0_370 br_0_370 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c370
+ bl_0_370 br_0_370 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c370
+ bl_0_370 br_0_370 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c370
+ bl_0_370 br_0_370 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c370
+ bl_0_370 br_0_370 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c370
+ bl_0_370 br_0_370 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c370
+ bl_0_370 br_0_370 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c370
+ bl_0_370 br_0_370 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c370
+ bl_0_370 br_0_370 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c370
+ bl_0_370 br_0_370 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c370
+ bl_0_370 br_0_370 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c370
+ bl_0_370 br_0_370 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c370
+ bl_0_370 br_0_370 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c370
+ bl_0_370 br_0_370 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c371
+ bl_0_371 br_0_371 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c371
+ bl_0_371 br_0_371 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c371
+ bl_0_371 br_0_371 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c371
+ bl_0_371 br_0_371 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c371
+ bl_0_371 br_0_371 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c371
+ bl_0_371 br_0_371 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c371
+ bl_0_371 br_0_371 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c371
+ bl_0_371 br_0_371 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c371
+ bl_0_371 br_0_371 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c371
+ bl_0_371 br_0_371 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c371
+ bl_0_371 br_0_371 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c371
+ bl_0_371 br_0_371 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c371
+ bl_0_371 br_0_371 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c371
+ bl_0_371 br_0_371 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c371
+ bl_0_371 br_0_371 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c371
+ bl_0_371 br_0_371 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c371
+ bl_0_371 br_0_371 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c371
+ bl_0_371 br_0_371 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c371
+ bl_0_371 br_0_371 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c371
+ bl_0_371 br_0_371 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c371
+ bl_0_371 br_0_371 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c371
+ bl_0_371 br_0_371 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c371
+ bl_0_371 br_0_371 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c371
+ bl_0_371 br_0_371 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c371
+ bl_0_371 br_0_371 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c371
+ bl_0_371 br_0_371 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c371
+ bl_0_371 br_0_371 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c371
+ bl_0_371 br_0_371 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c371
+ bl_0_371 br_0_371 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c371
+ bl_0_371 br_0_371 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c371
+ bl_0_371 br_0_371 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c371
+ bl_0_371 br_0_371 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c371
+ bl_0_371 br_0_371 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c371
+ bl_0_371 br_0_371 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c371
+ bl_0_371 br_0_371 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c371
+ bl_0_371 br_0_371 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c371
+ bl_0_371 br_0_371 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c371
+ bl_0_371 br_0_371 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c371
+ bl_0_371 br_0_371 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c371
+ bl_0_371 br_0_371 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c371
+ bl_0_371 br_0_371 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c371
+ bl_0_371 br_0_371 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c371
+ bl_0_371 br_0_371 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c371
+ bl_0_371 br_0_371 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c371
+ bl_0_371 br_0_371 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c372
+ bl_0_372 br_0_372 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c372
+ bl_0_372 br_0_372 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c372
+ bl_0_372 br_0_372 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c372
+ bl_0_372 br_0_372 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c372
+ bl_0_372 br_0_372 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c372
+ bl_0_372 br_0_372 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c372
+ bl_0_372 br_0_372 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c372
+ bl_0_372 br_0_372 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c372
+ bl_0_372 br_0_372 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c372
+ bl_0_372 br_0_372 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c372
+ bl_0_372 br_0_372 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c372
+ bl_0_372 br_0_372 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c372
+ bl_0_372 br_0_372 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c372
+ bl_0_372 br_0_372 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c372
+ bl_0_372 br_0_372 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c372
+ bl_0_372 br_0_372 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c372
+ bl_0_372 br_0_372 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c372
+ bl_0_372 br_0_372 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c372
+ bl_0_372 br_0_372 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c372
+ bl_0_372 br_0_372 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c372
+ bl_0_372 br_0_372 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c372
+ bl_0_372 br_0_372 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c372
+ bl_0_372 br_0_372 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c372
+ bl_0_372 br_0_372 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c372
+ bl_0_372 br_0_372 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c372
+ bl_0_372 br_0_372 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c372
+ bl_0_372 br_0_372 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c372
+ bl_0_372 br_0_372 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c372
+ bl_0_372 br_0_372 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c372
+ bl_0_372 br_0_372 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c372
+ bl_0_372 br_0_372 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c372
+ bl_0_372 br_0_372 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c372
+ bl_0_372 br_0_372 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c372
+ bl_0_372 br_0_372 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c372
+ bl_0_372 br_0_372 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c372
+ bl_0_372 br_0_372 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c372
+ bl_0_372 br_0_372 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c372
+ bl_0_372 br_0_372 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c372
+ bl_0_372 br_0_372 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c372
+ bl_0_372 br_0_372 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c372
+ bl_0_372 br_0_372 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c372
+ bl_0_372 br_0_372 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c372
+ bl_0_372 br_0_372 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c372
+ bl_0_372 br_0_372 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c372
+ bl_0_372 br_0_372 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c373
+ bl_0_373 br_0_373 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c373
+ bl_0_373 br_0_373 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c373
+ bl_0_373 br_0_373 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c373
+ bl_0_373 br_0_373 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c373
+ bl_0_373 br_0_373 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c373
+ bl_0_373 br_0_373 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c373
+ bl_0_373 br_0_373 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c373
+ bl_0_373 br_0_373 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c373
+ bl_0_373 br_0_373 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c373
+ bl_0_373 br_0_373 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c373
+ bl_0_373 br_0_373 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c373
+ bl_0_373 br_0_373 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c373
+ bl_0_373 br_0_373 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c373
+ bl_0_373 br_0_373 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c373
+ bl_0_373 br_0_373 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c373
+ bl_0_373 br_0_373 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c373
+ bl_0_373 br_0_373 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c373
+ bl_0_373 br_0_373 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c373
+ bl_0_373 br_0_373 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c373
+ bl_0_373 br_0_373 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c373
+ bl_0_373 br_0_373 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c373
+ bl_0_373 br_0_373 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c373
+ bl_0_373 br_0_373 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c373
+ bl_0_373 br_0_373 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c373
+ bl_0_373 br_0_373 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c373
+ bl_0_373 br_0_373 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c373
+ bl_0_373 br_0_373 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c373
+ bl_0_373 br_0_373 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c373
+ bl_0_373 br_0_373 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c373
+ bl_0_373 br_0_373 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c373
+ bl_0_373 br_0_373 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c373
+ bl_0_373 br_0_373 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c373
+ bl_0_373 br_0_373 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c373
+ bl_0_373 br_0_373 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c373
+ bl_0_373 br_0_373 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c373
+ bl_0_373 br_0_373 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c373
+ bl_0_373 br_0_373 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c373
+ bl_0_373 br_0_373 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c373
+ bl_0_373 br_0_373 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c373
+ bl_0_373 br_0_373 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c373
+ bl_0_373 br_0_373 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c373
+ bl_0_373 br_0_373 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c373
+ bl_0_373 br_0_373 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c373
+ bl_0_373 br_0_373 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c373
+ bl_0_373 br_0_373 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c374
+ bl_0_374 br_0_374 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c374
+ bl_0_374 br_0_374 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c374
+ bl_0_374 br_0_374 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c374
+ bl_0_374 br_0_374 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c374
+ bl_0_374 br_0_374 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c374
+ bl_0_374 br_0_374 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c374
+ bl_0_374 br_0_374 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c374
+ bl_0_374 br_0_374 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c374
+ bl_0_374 br_0_374 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c374
+ bl_0_374 br_0_374 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c374
+ bl_0_374 br_0_374 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c374
+ bl_0_374 br_0_374 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c374
+ bl_0_374 br_0_374 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c374
+ bl_0_374 br_0_374 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c374
+ bl_0_374 br_0_374 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c374
+ bl_0_374 br_0_374 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c374
+ bl_0_374 br_0_374 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c374
+ bl_0_374 br_0_374 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c374
+ bl_0_374 br_0_374 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c374
+ bl_0_374 br_0_374 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c374
+ bl_0_374 br_0_374 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c374
+ bl_0_374 br_0_374 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c374
+ bl_0_374 br_0_374 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c374
+ bl_0_374 br_0_374 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c374
+ bl_0_374 br_0_374 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c374
+ bl_0_374 br_0_374 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c374
+ bl_0_374 br_0_374 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c374
+ bl_0_374 br_0_374 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c374
+ bl_0_374 br_0_374 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c374
+ bl_0_374 br_0_374 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c374
+ bl_0_374 br_0_374 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c374
+ bl_0_374 br_0_374 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c374
+ bl_0_374 br_0_374 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c374
+ bl_0_374 br_0_374 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c374
+ bl_0_374 br_0_374 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c374
+ bl_0_374 br_0_374 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c374
+ bl_0_374 br_0_374 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c374
+ bl_0_374 br_0_374 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c374
+ bl_0_374 br_0_374 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c374
+ bl_0_374 br_0_374 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c374
+ bl_0_374 br_0_374 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c374
+ bl_0_374 br_0_374 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c374
+ bl_0_374 br_0_374 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c374
+ bl_0_374 br_0_374 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c374
+ bl_0_374 br_0_374 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c375
+ bl_0_375 br_0_375 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c375
+ bl_0_375 br_0_375 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c375
+ bl_0_375 br_0_375 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c375
+ bl_0_375 br_0_375 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c375
+ bl_0_375 br_0_375 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c375
+ bl_0_375 br_0_375 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c375
+ bl_0_375 br_0_375 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c375
+ bl_0_375 br_0_375 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c375
+ bl_0_375 br_0_375 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c375
+ bl_0_375 br_0_375 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c375
+ bl_0_375 br_0_375 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c375
+ bl_0_375 br_0_375 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c375
+ bl_0_375 br_0_375 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c375
+ bl_0_375 br_0_375 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c375
+ bl_0_375 br_0_375 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c375
+ bl_0_375 br_0_375 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c375
+ bl_0_375 br_0_375 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c375
+ bl_0_375 br_0_375 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c375
+ bl_0_375 br_0_375 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c375
+ bl_0_375 br_0_375 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c375
+ bl_0_375 br_0_375 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c375
+ bl_0_375 br_0_375 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c375
+ bl_0_375 br_0_375 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c375
+ bl_0_375 br_0_375 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c375
+ bl_0_375 br_0_375 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c375
+ bl_0_375 br_0_375 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c375
+ bl_0_375 br_0_375 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c375
+ bl_0_375 br_0_375 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c375
+ bl_0_375 br_0_375 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c375
+ bl_0_375 br_0_375 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c375
+ bl_0_375 br_0_375 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c375
+ bl_0_375 br_0_375 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c375
+ bl_0_375 br_0_375 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c375
+ bl_0_375 br_0_375 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c375
+ bl_0_375 br_0_375 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c375
+ bl_0_375 br_0_375 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c375
+ bl_0_375 br_0_375 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c375
+ bl_0_375 br_0_375 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c375
+ bl_0_375 br_0_375 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c375
+ bl_0_375 br_0_375 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c375
+ bl_0_375 br_0_375 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c375
+ bl_0_375 br_0_375 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c375
+ bl_0_375 br_0_375 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c375
+ bl_0_375 br_0_375 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c375
+ bl_0_375 br_0_375 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c376
+ bl_0_376 br_0_376 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c376
+ bl_0_376 br_0_376 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c376
+ bl_0_376 br_0_376 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c376
+ bl_0_376 br_0_376 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c376
+ bl_0_376 br_0_376 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c376
+ bl_0_376 br_0_376 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c376
+ bl_0_376 br_0_376 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c376
+ bl_0_376 br_0_376 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c376
+ bl_0_376 br_0_376 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c376
+ bl_0_376 br_0_376 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c376
+ bl_0_376 br_0_376 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c376
+ bl_0_376 br_0_376 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c376
+ bl_0_376 br_0_376 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c376
+ bl_0_376 br_0_376 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c376
+ bl_0_376 br_0_376 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c376
+ bl_0_376 br_0_376 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c376
+ bl_0_376 br_0_376 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c376
+ bl_0_376 br_0_376 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c376
+ bl_0_376 br_0_376 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c376
+ bl_0_376 br_0_376 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c376
+ bl_0_376 br_0_376 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c376
+ bl_0_376 br_0_376 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c376
+ bl_0_376 br_0_376 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c376
+ bl_0_376 br_0_376 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c376
+ bl_0_376 br_0_376 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c376
+ bl_0_376 br_0_376 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c376
+ bl_0_376 br_0_376 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c376
+ bl_0_376 br_0_376 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c376
+ bl_0_376 br_0_376 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c376
+ bl_0_376 br_0_376 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c376
+ bl_0_376 br_0_376 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c376
+ bl_0_376 br_0_376 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c376
+ bl_0_376 br_0_376 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c376
+ bl_0_376 br_0_376 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c376
+ bl_0_376 br_0_376 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c376
+ bl_0_376 br_0_376 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c376
+ bl_0_376 br_0_376 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c376
+ bl_0_376 br_0_376 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c376
+ bl_0_376 br_0_376 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c376
+ bl_0_376 br_0_376 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c376
+ bl_0_376 br_0_376 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c376
+ bl_0_376 br_0_376 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c376
+ bl_0_376 br_0_376 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c376
+ bl_0_376 br_0_376 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c376
+ bl_0_376 br_0_376 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c377
+ bl_0_377 br_0_377 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c377
+ bl_0_377 br_0_377 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c377
+ bl_0_377 br_0_377 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c377
+ bl_0_377 br_0_377 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c377
+ bl_0_377 br_0_377 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c377
+ bl_0_377 br_0_377 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c377
+ bl_0_377 br_0_377 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c377
+ bl_0_377 br_0_377 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c377
+ bl_0_377 br_0_377 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c377
+ bl_0_377 br_0_377 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c377
+ bl_0_377 br_0_377 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c377
+ bl_0_377 br_0_377 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c377
+ bl_0_377 br_0_377 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c377
+ bl_0_377 br_0_377 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c377
+ bl_0_377 br_0_377 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c377
+ bl_0_377 br_0_377 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c377
+ bl_0_377 br_0_377 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c377
+ bl_0_377 br_0_377 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c377
+ bl_0_377 br_0_377 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c377
+ bl_0_377 br_0_377 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c377
+ bl_0_377 br_0_377 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c377
+ bl_0_377 br_0_377 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c377
+ bl_0_377 br_0_377 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c377
+ bl_0_377 br_0_377 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c377
+ bl_0_377 br_0_377 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c377
+ bl_0_377 br_0_377 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c377
+ bl_0_377 br_0_377 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c377
+ bl_0_377 br_0_377 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c377
+ bl_0_377 br_0_377 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c377
+ bl_0_377 br_0_377 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c377
+ bl_0_377 br_0_377 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c377
+ bl_0_377 br_0_377 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c377
+ bl_0_377 br_0_377 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c377
+ bl_0_377 br_0_377 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c377
+ bl_0_377 br_0_377 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c377
+ bl_0_377 br_0_377 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c377
+ bl_0_377 br_0_377 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c377
+ bl_0_377 br_0_377 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c377
+ bl_0_377 br_0_377 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c377
+ bl_0_377 br_0_377 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c377
+ bl_0_377 br_0_377 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c377
+ bl_0_377 br_0_377 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c377
+ bl_0_377 br_0_377 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c377
+ bl_0_377 br_0_377 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c377
+ bl_0_377 br_0_377 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c378
+ bl_0_378 br_0_378 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c378
+ bl_0_378 br_0_378 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c378
+ bl_0_378 br_0_378 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c378
+ bl_0_378 br_0_378 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c378
+ bl_0_378 br_0_378 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c378
+ bl_0_378 br_0_378 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c378
+ bl_0_378 br_0_378 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c378
+ bl_0_378 br_0_378 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c378
+ bl_0_378 br_0_378 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c378
+ bl_0_378 br_0_378 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c378
+ bl_0_378 br_0_378 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c378
+ bl_0_378 br_0_378 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c378
+ bl_0_378 br_0_378 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c378
+ bl_0_378 br_0_378 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c378
+ bl_0_378 br_0_378 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c378
+ bl_0_378 br_0_378 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c378
+ bl_0_378 br_0_378 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c378
+ bl_0_378 br_0_378 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c378
+ bl_0_378 br_0_378 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c378
+ bl_0_378 br_0_378 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c378
+ bl_0_378 br_0_378 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c378
+ bl_0_378 br_0_378 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c378
+ bl_0_378 br_0_378 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c378
+ bl_0_378 br_0_378 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c378
+ bl_0_378 br_0_378 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c378
+ bl_0_378 br_0_378 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c378
+ bl_0_378 br_0_378 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c378
+ bl_0_378 br_0_378 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c378
+ bl_0_378 br_0_378 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c378
+ bl_0_378 br_0_378 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c378
+ bl_0_378 br_0_378 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c378
+ bl_0_378 br_0_378 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c378
+ bl_0_378 br_0_378 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c378
+ bl_0_378 br_0_378 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c378
+ bl_0_378 br_0_378 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c378
+ bl_0_378 br_0_378 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c378
+ bl_0_378 br_0_378 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c378
+ bl_0_378 br_0_378 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c378
+ bl_0_378 br_0_378 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c378
+ bl_0_378 br_0_378 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c378
+ bl_0_378 br_0_378 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c378
+ bl_0_378 br_0_378 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c378
+ bl_0_378 br_0_378 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c378
+ bl_0_378 br_0_378 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c378
+ bl_0_378 br_0_378 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c379
+ bl_0_379 br_0_379 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c379
+ bl_0_379 br_0_379 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c379
+ bl_0_379 br_0_379 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c379
+ bl_0_379 br_0_379 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c379
+ bl_0_379 br_0_379 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c379
+ bl_0_379 br_0_379 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c379
+ bl_0_379 br_0_379 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c379
+ bl_0_379 br_0_379 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c379
+ bl_0_379 br_0_379 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c379
+ bl_0_379 br_0_379 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c379
+ bl_0_379 br_0_379 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c379
+ bl_0_379 br_0_379 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c379
+ bl_0_379 br_0_379 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c379
+ bl_0_379 br_0_379 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c379
+ bl_0_379 br_0_379 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c379
+ bl_0_379 br_0_379 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c379
+ bl_0_379 br_0_379 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c379
+ bl_0_379 br_0_379 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c379
+ bl_0_379 br_0_379 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c379
+ bl_0_379 br_0_379 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c379
+ bl_0_379 br_0_379 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c379
+ bl_0_379 br_0_379 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c379
+ bl_0_379 br_0_379 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c379
+ bl_0_379 br_0_379 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c379
+ bl_0_379 br_0_379 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c379
+ bl_0_379 br_0_379 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c379
+ bl_0_379 br_0_379 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c379
+ bl_0_379 br_0_379 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c379
+ bl_0_379 br_0_379 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c379
+ bl_0_379 br_0_379 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c379
+ bl_0_379 br_0_379 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c379
+ bl_0_379 br_0_379 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c379
+ bl_0_379 br_0_379 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c379
+ bl_0_379 br_0_379 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c379
+ bl_0_379 br_0_379 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c379
+ bl_0_379 br_0_379 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c379
+ bl_0_379 br_0_379 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c379
+ bl_0_379 br_0_379 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c379
+ bl_0_379 br_0_379 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c379
+ bl_0_379 br_0_379 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c379
+ bl_0_379 br_0_379 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c379
+ bl_0_379 br_0_379 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c379
+ bl_0_379 br_0_379 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c379
+ bl_0_379 br_0_379 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c379
+ bl_0_379 br_0_379 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c380
+ bl_0_380 br_0_380 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c380
+ bl_0_380 br_0_380 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c380
+ bl_0_380 br_0_380 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c380
+ bl_0_380 br_0_380 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c380
+ bl_0_380 br_0_380 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c380
+ bl_0_380 br_0_380 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c380
+ bl_0_380 br_0_380 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c380
+ bl_0_380 br_0_380 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c380
+ bl_0_380 br_0_380 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c380
+ bl_0_380 br_0_380 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c380
+ bl_0_380 br_0_380 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c380
+ bl_0_380 br_0_380 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c380
+ bl_0_380 br_0_380 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c380
+ bl_0_380 br_0_380 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c380
+ bl_0_380 br_0_380 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c380
+ bl_0_380 br_0_380 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c380
+ bl_0_380 br_0_380 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c380
+ bl_0_380 br_0_380 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c380
+ bl_0_380 br_0_380 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c380
+ bl_0_380 br_0_380 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c380
+ bl_0_380 br_0_380 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c380
+ bl_0_380 br_0_380 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c380
+ bl_0_380 br_0_380 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c380
+ bl_0_380 br_0_380 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c380
+ bl_0_380 br_0_380 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c380
+ bl_0_380 br_0_380 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c380
+ bl_0_380 br_0_380 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c380
+ bl_0_380 br_0_380 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c380
+ bl_0_380 br_0_380 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c380
+ bl_0_380 br_0_380 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c380
+ bl_0_380 br_0_380 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c380
+ bl_0_380 br_0_380 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c380
+ bl_0_380 br_0_380 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c380
+ bl_0_380 br_0_380 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c380
+ bl_0_380 br_0_380 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c380
+ bl_0_380 br_0_380 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c380
+ bl_0_380 br_0_380 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c380
+ bl_0_380 br_0_380 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c380
+ bl_0_380 br_0_380 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c380
+ bl_0_380 br_0_380 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c380
+ bl_0_380 br_0_380 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c380
+ bl_0_380 br_0_380 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c380
+ bl_0_380 br_0_380 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c380
+ bl_0_380 br_0_380 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c380
+ bl_0_380 br_0_380 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c381
+ bl_0_381 br_0_381 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c381
+ bl_0_381 br_0_381 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c381
+ bl_0_381 br_0_381 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c381
+ bl_0_381 br_0_381 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c381
+ bl_0_381 br_0_381 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c381
+ bl_0_381 br_0_381 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c381
+ bl_0_381 br_0_381 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c381
+ bl_0_381 br_0_381 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c381
+ bl_0_381 br_0_381 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c381
+ bl_0_381 br_0_381 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c381
+ bl_0_381 br_0_381 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c381
+ bl_0_381 br_0_381 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c381
+ bl_0_381 br_0_381 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c381
+ bl_0_381 br_0_381 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c381
+ bl_0_381 br_0_381 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c381
+ bl_0_381 br_0_381 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c381
+ bl_0_381 br_0_381 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c381
+ bl_0_381 br_0_381 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c381
+ bl_0_381 br_0_381 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c381
+ bl_0_381 br_0_381 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c381
+ bl_0_381 br_0_381 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c381
+ bl_0_381 br_0_381 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c381
+ bl_0_381 br_0_381 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c381
+ bl_0_381 br_0_381 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c381
+ bl_0_381 br_0_381 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c381
+ bl_0_381 br_0_381 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c381
+ bl_0_381 br_0_381 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c381
+ bl_0_381 br_0_381 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c381
+ bl_0_381 br_0_381 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c381
+ bl_0_381 br_0_381 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c381
+ bl_0_381 br_0_381 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c381
+ bl_0_381 br_0_381 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c381
+ bl_0_381 br_0_381 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c381
+ bl_0_381 br_0_381 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c381
+ bl_0_381 br_0_381 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c381
+ bl_0_381 br_0_381 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c381
+ bl_0_381 br_0_381 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c381
+ bl_0_381 br_0_381 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c381
+ bl_0_381 br_0_381 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c381
+ bl_0_381 br_0_381 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c381
+ bl_0_381 br_0_381 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c381
+ bl_0_381 br_0_381 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c381
+ bl_0_381 br_0_381 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c381
+ bl_0_381 br_0_381 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c381
+ bl_0_381 br_0_381 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c382
+ bl_0_382 br_0_382 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c382
+ bl_0_382 br_0_382 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c382
+ bl_0_382 br_0_382 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c382
+ bl_0_382 br_0_382 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c382
+ bl_0_382 br_0_382 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c382
+ bl_0_382 br_0_382 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c382
+ bl_0_382 br_0_382 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c382
+ bl_0_382 br_0_382 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c382
+ bl_0_382 br_0_382 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c382
+ bl_0_382 br_0_382 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c382
+ bl_0_382 br_0_382 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c382
+ bl_0_382 br_0_382 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c382
+ bl_0_382 br_0_382 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c382
+ bl_0_382 br_0_382 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c382
+ bl_0_382 br_0_382 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c382
+ bl_0_382 br_0_382 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c382
+ bl_0_382 br_0_382 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c382
+ bl_0_382 br_0_382 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c382
+ bl_0_382 br_0_382 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c382
+ bl_0_382 br_0_382 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c382
+ bl_0_382 br_0_382 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c382
+ bl_0_382 br_0_382 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c382
+ bl_0_382 br_0_382 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c382
+ bl_0_382 br_0_382 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c382
+ bl_0_382 br_0_382 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c382
+ bl_0_382 br_0_382 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c382
+ bl_0_382 br_0_382 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c382
+ bl_0_382 br_0_382 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c382
+ bl_0_382 br_0_382 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c382
+ bl_0_382 br_0_382 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c382
+ bl_0_382 br_0_382 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c382
+ bl_0_382 br_0_382 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c382
+ bl_0_382 br_0_382 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c382
+ bl_0_382 br_0_382 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c382
+ bl_0_382 br_0_382 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c382
+ bl_0_382 br_0_382 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c382
+ bl_0_382 br_0_382 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c382
+ bl_0_382 br_0_382 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c382
+ bl_0_382 br_0_382 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c382
+ bl_0_382 br_0_382 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c382
+ bl_0_382 br_0_382 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c382
+ bl_0_382 br_0_382 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c382
+ bl_0_382 br_0_382 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c382
+ bl_0_382 br_0_382 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c382
+ bl_0_382 br_0_382 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c383
+ bl_0_383 br_0_383 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c383
+ bl_0_383 br_0_383 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c383
+ bl_0_383 br_0_383 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c383
+ bl_0_383 br_0_383 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c383
+ bl_0_383 br_0_383 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c383
+ bl_0_383 br_0_383 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c383
+ bl_0_383 br_0_383 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c383
+ bl_0_383 br_0_383 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c383
+ bl_0_383 br_0_383 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c383
+ bl_0_383 br_0_383 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c383
+ bl_0_383 br_0_383 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c383
+ bl_0_383 br_0_383 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c383
+ bl_0_383 br_0_383 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c383
+ bl_0_383 br_0_383 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c383
+ bl_0_383 br_0_383 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c383
+ bl_0_383 br_0_383 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c383
+ bl_0_383 br_0_383 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c383
+ bl_0_383 br_0_383 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c383
+ bl_0_383 br_0_383 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c383
+ bl_0_383 br_0_383 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c383
+ bl_0_383 br_0_383 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c383
+ bl_0_383 br_0_383 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c383
+ bl_0_383 br_0_383 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c383
+ bl_0_383 br_0_383 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c383
+ bl_0_383 br_0_383 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c383
+ bl_0_383 br_0_383 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c383
+ bl_0_383 br_0_383 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c383
+ bl_0_383 br_0_383 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c383
+ bl_0_383 br_0_383 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c383
+ bl_0_383 br_0_383 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c383
+ bl_0_383 br_0_383 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c383
+ bl_0_383 br_0_383 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c383
+ bl_0_383 br_0_383 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c383
+ bl_0_383 br_0_383 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c383
+ bl_0_383 br_0_383 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c383
+ bl_0_383 br_0_383 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c383
+ bl_0_383 br_0_383 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c383
+ bl_0_383 br_0_383 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c383
+ bl_0_383 br_0_383 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c383
+ bl_0_383 br_0_383 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c383
+ bl_0_383 br_0_383 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c383
+ bl_0_383 br_0_383 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c383
+ bl_0_383 br_0_383 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c383
+ bl_0_383 br_0_383 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c383
+ bl_0_383 br_0_383 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c384
+ bl_0_384 br_0_384 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c384
+ bl_0_384 br_0_384 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c384
+ bl_0_384 br_0_384 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c384
+ bl_0_384 br_0_384 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c384
+ bl_0_384 br_0_384 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c384
+ bl_0_384 br_0_384 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c384
+ bl_0_384 br_0_384 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c384
+ bl_0_384 br_0_384 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c384
+ bl_0_384 br_0_384 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c384
+ bl_0_384 br_0_384 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c384
+ bl_0_384 br_0_384 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c384
+ bl_0_384 br_0_384 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c384
+ bl_0_384 br_0_384 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c384
+ bl_0_384 br_0_384 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c384
+ bl_0_384 br_0_384 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c384
+ bl_0_384 br_0_384 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c384
+ bl_0_384 br_0_384 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c384
+ bl_0_384 br_0_384 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c384
+ bl_0_384 br_0_384 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c384
+ bl_0_384 br_0_384 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c384
+ bl_0_384 br_0_384 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c384
+ bl_0_384 br_0_384 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c384
+ bl_0_384 br_0_384 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c384
+ bl_0_384 br_0_384 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c384
+ bl_0_384 br_0_384 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c384
+ bl_0_384 br_0_384 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c384
+ bl_0_384 br_0_384 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c384
+ bl_0_384 br_0_384 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c384
+ bl_0_384 br_0_384 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c384
+ bl_0_384 br_0_384 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c384
+ bl_0_384 br_0_384 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c384
+ bl_0_384 br_0_384 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c384
+ bl_0_384 br_0_384 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c384
+ bl_0_384 br_0_384 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c384
+ bl_0_384 br_0_384 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c384
+ bl_0_384 br_0_384 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c384
+ bl_0_384 br_0_384 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c384
+ bl_0_384 br_0_384 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c384
+ bl_0_384 br_0_384 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c384
+ bl_0_384 br_0_384 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c384
+ bl_0_384 br_0_384 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c384
+ bl_0_384 br_0_384 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c384
+ bl_0_384 br_0_384 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c384
+ bl_0_384 br_0_384 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c384
+ bl_0_384 br_0_384 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c385
+ bl_0_385 br_0_385 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c385
+ bl_0_385 br_0_385 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c385
+ bl_0_385 br_0_385 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c385
+ bl_0_385 br_0_385 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c385
+ bl_0_385 br_0_385 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c385
+ bl_0_385 br_0_385 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c385
+ bl_0_385 br_0_385 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c385
+ bl_0_385 br_0_385 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c385
+ bl_0_385 br_0_385 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c385
+ bl_0_385 br_0_385 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c385
+ bl_0_385 br_0_385 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c385
+ bl_0_385 br_0_385 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c385
+ bl_0_385 br_0_385 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c385
+ bl_0_385 br_0_385 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c385
+ bl_0_385 br_0_385 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c385
+ bl_0_385 br_0_385 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c385
+ bl_0_385 br_0_385 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c385
+ bl_0_385 br_0_385 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c385
+ bl_0_385 br_0_385 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c385
+ bl_0_385 br_0_385 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c385
+ bl_0_385 br_0_385 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c385
+ bl_0_385 br_0_385 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c385
+ bl_0_385 br_0_385 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c385
+ bl_0_385 br_0_385 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c385
+ bl_0_385 br_0_385 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c385
+ bl_0_385 br_0_385 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c385
+ bl_0_385 br_0_385 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c385
+ bl_0_385 br_0_385 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c385
+ bl_0_385 br_0_385 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c385
+ bl_0_385 br_0_385 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c385
+ bl_0_385 br_0_385 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c385
+ bl_0_385 br_0_385 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c385
+ bl_0_385 br_0_385 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c385
+ bl_0_385 br_0_385 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c385
+ bl_0_385 br_0_385 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c385
+ bl_0_385 br_0_385 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c385
+ bl_0_385 br_0_385 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c385
+ bl_0_385 br_0_385 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c385
+ bl_0_385 br_0_385 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c385
+ bl_0_385 br_0_385 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c385
+ bl_0_385 br_0_385 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c385
+ bl_0_385 br_0_385 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c385
+ bl_0_385 br_0_385 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c385
+ bl_0_385 br_0_385 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c385
+ bl_0_385 br_0_385 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c386
+ bl_0_386 br_0_386 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c386
+ bl_0_386 br_0_386 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c386
+ bl_0_386 br_0_386 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c386
+ bl_0_386 br_0_386 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c386
+ bl_0_386 br_0_386 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c386
+ bl_0_386 br_0_386 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c386
+ bl_0_386 br_0_386 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c386
+ bl_0_386 br_0_386 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c386
+ bl_0_386 br_0_386 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c386
+ bl_0_386 br_0_386 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c386
+ bl_0_386 br_0_386 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c386
+ bl_0_386 br_0_386 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c386
+ bl_0_386 br_0_386 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c386
+ bl_0_386 br_0_386 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c386
+ bl_0_386 br_0_386 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c386
+ bl_0_386 br_0_386 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c386
+ bl_0_386 br_0_386 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c386
+ bl_0_386 br_0_386 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c386
+ bl_0_386 br_0_386 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c386
+ bl_0_386 br_0_386 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c386
+ bl_0_386 br_0_386 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c386
+ bl_0_386 br_0_386 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c386
+ bl_0_386 br_0_386 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c386
+ bl_0_386 br_0_386 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c386
+ bl_0_386 br_0_386 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c386
+ bl_0_386 br_0_386 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c386
+ bl_0_386 br_0_386 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c386
+ bl_0_386 br_0_386 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c386
+ bl_0_386 br_0_386 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c386
+ bl_0_386 br_0_386 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c386
+ bl_0_386 br_0_386 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c386
+ bl_0_386 br_0_386 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c386
+ bl_0_386 br_0_386 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c386
+ bl_0_386 br_0_386 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c386
+ bl_0_386 br_0_386 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c386
+ bl_0_386 br_0_386 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c386
+ bl_0_386 br_0_386 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c386
+ bl_0_386 br_0_386 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c386
+ bl_0_386 br_0_386 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c386
+ bl_0_386 br_0_386 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c386
+ bl_0_386 br_0_386 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c386
+ bl_0_386 br_0_386 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c386
+ bl_0_386 br_0_386 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c386
+ bl_0_386 br_0_386 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c386
+ bl_0_386 br_0_386 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c387
+ bl_0_387 br_0_387 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c387
+ bl_0_387 br_0_387 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c387
+ bl_0_387 br_0_387 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c387
+ bl_0_387 br_0_387 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c387
+ bl_0_387 br_0_387 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c387
+ bl_0_387 br_0_387 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c387
+ bl_0_387 br_0_387 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c387
+ bl_0_387 br_0_387 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c387
+ bl_0_387 br_0_387 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c387
+ bl_0_387 br_0_387 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c387
+ bl_0_387 br_0_387 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c387
+ bl_0_387 br_0_387 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c387
+ bl_0_387 br_0_387 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c387
+ bl_0_387 br_0_387 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c387
+ bl_0_387 br_0_387 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c387
+ bl_0_387 br_0_387 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c387
+ bl_0_387 br_0_387 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c387
+ bl_0_387 br_0_387 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c387
+ bl_0_387 br_0_387 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c387
+ bl_0_387 br_0_387 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c387
+ bl_0_387 br_0_387 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c387
+ bl_0_387 br_0_387 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c387
+ bl_0_387 br_0_387 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c387
+ bl_0_387 br_0_387 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c387
+ bl_0_387 br_0_387 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c387
+ bl_0_387 br_0_387 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c387
+ bl_0_387 br_0_387 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c387
+ bl_0_387 br_0_387 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c387
+ bl_0_387 br_0_387 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c387
+ bl_0_387 br_0_387 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c387
+ bl_0_387 br_0_387 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c387
+ bl_0_387 br_0_387 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c387
+ bl_0_387 br_0_387 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c387
+ bl_0_387 br_0_387 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c387
+ bl_0_387 br_0_387 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c387
+ bl_0_387 br_0_387 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c387
+ bl_0_387 br_0_387 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c387
+ bl_0_387 br_0_387 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c387
+ bl_0_387 br_0_387 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c387
+ bl_0_387 br_0_387 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c387
+ bl_0_387 br_0_387 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c387
+ bl_0_387 br_0_387 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c387
+ bl_0_387 br_0_387 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c387
+ bl_0_387 br_0_387 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c387
+ bl_0_387 br_0_387 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c388
+ bl_0_388 br_0_388 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c388
+ bl_0_388 br_0_388 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c388
+ bl_0_388 br_0_388 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c388
+ bl_0_388 br_0_388 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c388
+ bl_0_388 br_0_388 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c388
+ bl_0_388 br_0_388 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c388
+ bl_0_388 br_0_388 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c388
+ bl_0_388 br_0_388 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c388
+ bl_0_388 br_0_388 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c388
+ bl_0_388 br_0_388 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c388
+ bl_0_388 br_0_388 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c388
+ bl_0_388 br_0_388 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c388
+ bl_0_388 br_0_388 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c388
+ bl_0_388 br_0_388 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c388
+ bl_0_388 br_0_388 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c388
+ bl_0_388 br_0_388 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c388
+ bl_0_388 br_0_388 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c388
+ bl_0_388 br_0_388 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c388
+ bl_0_388 br_0_388 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c388
+ bl_0_388 br_0_388 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c388
+ bl_0_388 br_0_388 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c388
+ bl_0_388 br_0_388 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c388
+ bl_0_388 br_0_388 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c388
+ bl_0_388 br_0_388 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c388
+ bl_0_388 br_0_388 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c388
+ bl_0_388 br_0_388 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c388
+ bl_0_388 br_0_388 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c388
+ bl_0_388 br_0_388 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c388
+ bl_0_388 br_0_388 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c388
+ bl_0_388 br_0_388 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c388
+ bl_0_388 br_0_388 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c388
+ bl_0_388 br_0_388 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c388
+ bl_0_388 br_0_388 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c388
+ bl_0_388 br_0_388 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c388
+ bl_0_388 br_0_388 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c388
+ bl_0_388 br_0_388 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c388
+ bl_0_388 br_0_388 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c388
+ bl_0_388 br_0_388 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c388
+ bl_0_388 br_0_388 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c388
+ bl_0_388 br_0_388 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c388
+ bl_0_388 br_0_388 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c388
+ bl_0_388 br_0_388 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c388
+ bl_0_388 br_0_388 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c388
+ bl_0_388 br_0_388 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c388
+ bl_0_388 br_0_388 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c389
+ bl_0_389 br_0_389 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c389
+ bl_0_389 br_0_389 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c389
+ bl_0_389 br_0_389 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c389
+ bl_0_389 br_0_389 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c389
+ bl_0_389 br_0_389 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c389
+ bl_0_389 br_0_389 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c389
+ bl_0_389 br_0_389 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c389
+ bl_0_389 br_0_389 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c389
+ bl_0_389 br_0_389 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c389
+ bl_0_389 br_0_389 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c389
+ bl_0_389 br_0_389 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c389
+ bl_0_389 br_0_389 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c389
+ bl_0_389 br_0_389 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c389
+ bl_0_389 br_0_389 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c389
+ bl_0_389 br_0_389 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c389
+ bl_0_389 br_0_389 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c389
+ bl_0_389 br_0_389 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c389
+ bl_0_389 br_0_389 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c389
+ bl_0_389 br_0_389 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c389
+ bl_0_389 br_0_389 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c389
+ bl_0_389 br_0_389 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c389
+ bl_0_389 br_0_389 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c389
+ bl_0_389 br_0_389 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c389
+ bl_0_389 br_0_389 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c389
+ bl_0_389 br_0_389 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c389
+ bl_0_389 br_0_389 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c389
+ bl_0_389 br_0_389 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c389
+ bl_0_389 br_0_389 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c389
+ bl_0_389 br_0_389 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c389
+ bl_0_389 br_0_389 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c389
+ bl_0_389 br_0_389 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c389
+ bl_0_389 br_0_389 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c389
+ bl_0_389 br_0_389 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c389
+ bl_0_389 br_0_389 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c389
+ bl_0_389 br_0_389 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c389
+ bl_0_389 br_0_389 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c389
+ bl_0_389 br_0_389 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c389
+ bl_0_389 br_0_389 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c389
+ bl_0_389 br_0_389 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c389
+ bl_0_389 br_0_389 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c389
+ bl_0_389 br_0_389 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c389
+ bl_0_389 br_0_389 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c389
+ bl_0_389 br_0_389 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c389
+ bl_0_389 br_0_389 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c389
+ bl_0_389 br_0_389 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c390
+ bl_0_390 br_0_390 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c390
+ bl_0_390 br_0_390 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c390
+ bl_0_390 br_0_390 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c390
+ bl_0_390 br_0_390 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c390
+ bl_0_390 br_0_390 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c390
+ bl_0_390 br_0_390 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c390
+ bl_0_390 br_0_390 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c390
+ bl_0_390 br_0_390 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c390
+ bl_0_390 br_0_390 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c390
+ bl_0_390 br_0_390 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c390
+ bl_0_390 br_0_390 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c390
+ bl_0_390 br_0_390 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c390
+ bl_0_390 br_0_390 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c390
+ bl_0_390 br_0_390 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c390
+ bl_0_390 br_0_390 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c390
+ bl_0_390 br_0_390 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c390
+ bl_0_390 br_0_390 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c390
+ bl_0_390 br_0_390 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c390
+ bl_0_390 br_0_390 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c390
+ bl_0_390 br_0_390 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c390
+ bl_0_390 br_0_390 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c390
+ bl_0_390 br_0_390 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c390
+ bl_0_390 br_0_390 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c390
+ bl_0_390 br_0_390 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c390
+ bl_0_390 br_0_390 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c390
+ bl_0_390 br_0_390 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c390
+ bl_0_390 br_0_390 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c390
+ bl_0_390 br_0_390 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c390
+ bl_0_390 br_0_390 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c390
+ bl_0_390 br_0_390 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c390
+ bl_0_390 br_0_390 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c390
+ bl_0_390 br_0_390 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c390
+ bl_0_390 br_0_390 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c390
+ bl_0_390 br_0_390 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c390
+ bl_0_390 br_0_390 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c390
+ bl_0_390 br_0_390 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c390
+ bl_0_390 br_0_390 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c390
+ bl_0_390 br_0_390 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c390
+ bl_0_390 br_0_390 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c390
+ bl_0_390 br_0_390 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c390
+ bl_0_390 br_0_390 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c390
+ bl_0_390 br_0_390 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c390
+ bl_0_390 br_0_390 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c390
+ bl_0_390 br_0_390 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c390
+ bl_0_390 br_0_390 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c391
+ bl_0_391 br_0_391 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c391
+ bl_0_391 br_0_391 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c391
+ bl_0_391 br_0_391 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c391
+ bl_0_391 br_0_391 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c391
+ bl_0_391 br_0_391 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c391
+ bl_0_391 br_0_391 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c391
+ bl_0_391 br_0_391 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c391
+ bl_0_391 br_0_391 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c391
+ bl_0_391 br_0_391 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c391
+ bl_0_391 br_0_391 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c391
+ bl_0_391 br_0_391 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c391
+ bl_0_391 br_0_391 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c391
+ bl_0_391 br_0_391 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c391
+ bl_0_391 br_0_391 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c391
+ bl_0_391 br_0_391 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c391
+ bl_0_391 br_0_391 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c391
+ bl_0_391 br_0_391 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c391
+ bl_0_391 br_0_391 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c391
+ bl_0_391 br_0_391 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c391
+ bl_0_391 br_0_391 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c391
+ bl_0_391 br_0_391 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c391
+ bl_0_391 br_0_391 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c391
+ bl_0_391 br_0_391 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c391
+ bl_0_391 br_0_391 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c391
+ bl_0_391 br_0_391 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c391
+ bl_0_391 br_0_391 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c391
+ bl_0_391 br_0_391 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c391
+ bl_0_391 br_0_391 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c391
+ bl_0_391 br_0_391 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c391
+ bl_0_391 br_0_391 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c391
+ bl_0_391 br_0_391 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c391
+ bl_0_391 br_0_391 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c391
+ bl_0_391 br_0_391 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c391
+ bl_0_391 br_0_391 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c391
+ bl_0_391 br_0_391 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c391
+ bl_0_391 br_0_391 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c391
+ bl_0_391 br_0_391 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c391
+ bl_0_391 br_0_391 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c391
+ bl_0_391 br_0_391 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c391
+ bl_0_391 br_0_391 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c391
+ bl_0_391 br_0_391 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c391
+ bl_0_391 br_0_391 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c391
+ bl_0_391 br_0_391 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c391
+ bl_0_391 br_0_391 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c391
+ bl_0_391 br_0_391 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c392
+ bl_0_392 br_0_392 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c392
+ bl_0_392 br_0_392 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c392
+ bl_0_392 br_0_392 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c392
+ bl_0_392 br_0_392 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c392
+ bl_0_392 br_0_392 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c392
+ bl_0_392 br_0_392 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c392
+ bl_0_392 br_0_392 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c392
+ bl_0_392 br_0_392 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c392
+ bl_0_392 br_0_392 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c392
+ bl_0_392 br_0_392 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c392
+ bl_0_392 br_0_392 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c392
+ bl_0_392 br_0_392 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c392
+ bl_0_392 br_0_392 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c392
+ bl_0_392 br_0_392 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c392
+ bl_0_392 br_0_392 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c392
+ bl_0_392 br_0_392 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c392
+ bl_0_392 br_0_392 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c392
+ bl_0_392 br_0_392 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c392
+ bl_0_392 br_0_392 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c392
+ bl_0_392 br_0_392 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c392
+ bl_0_392 br_0_392 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c392
+ bl_0_392 br_0_392 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c392
+ bl_0_392 br_0_392 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c392
+ bl_0_392 br_0_392 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c392
+ bl_0_392 br_0_392 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c392
+ bl_0_392 br_0_392 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c392
+ bl_0_392 br_0_392 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c392
+ bl_0_392 br_0_392 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c392
+ bl_0_392 br_0_392 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c392
+ bl_0_392 br_0_392 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c392
+ bl_0_392 br_0_392 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c392
+ bl_0_392 br_0_392 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c392
+ bl_0_392 br_0_392 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c392
+ bl_0_392 br_0_392 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c392
+ bl_0_392 br_0_392 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c392
+ bl_0_392 br_0_392 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c392
+ bl_0_392 br_0_392 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c392
+ bl_0_392 br_0_392 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c392
+ bl_0_392 br_0_392 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c392
+ bl_0_392 br_0_392 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c392
+ bl_0_392 br_0_392 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c392
+ bl_0_392 br_0_392 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c392
+ bl_0_392 br_0_392 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c392
+ bl_0_392 br_0_392 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c392
+ bl_0_392 br_0_392 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c393
+ bl_0_393 br_0_393 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c393
+ bl_0_393 br_0_393 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c393
+ bl_0_393 br_0_393 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c393
+ bl_0_393 br_0_393 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c393
+ bl_0_393 br_0_393 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c393
+ bl_0_393 br_0_393 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c393
+ bl_0_393 br_0_393 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c393
+ bl_0_393 br_0_393 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c393
+ bl_0_393 br_0_393 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c393
+ bl_0_393 br_0_393 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c393
+ bl_0_393 br_0_393 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c393
+ bl_0_393 br_0_393 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c393
+ bl_0_393 br_0_393 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c393
+ bl_0_393 br_0_393 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c393
+ bl_0_393 br_0_393 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c393
+ bl_0_393 br_0_393 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c393
+ bl_0_393 br_0_393 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c393
+ bl_0_393 br_0_393 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c393
+ bl_0_393 br_0_393 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c393
+ bl_0_393 br_0_393 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c393
+ bl_0_393 br_0_393 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c393
+ bl_0_393 br_0_393 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c393
+ bl_0_393 br_0_393 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c393
+ bl_0_393 br_0_393 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c393
+ bl_0_393 br_0_393 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c393
+ bl_0_393 br_0_393 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c393
+ bl_0_393 br_0_393 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c393
+ bl_0_393 br_0_393 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c393
+ bl_0_393 br_0_393 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c393
+ bl_0_393 br_0_393 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c393
+ bl_0_393 br_0_393 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c393
+ bl_0_393 br_0_393 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c393
+ bl_0_393 br_0_393 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c393
+ bl_0_393 br_0_393 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c393
+ bl_0_393 br_0_393 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c393
+ bl_0_393 br_0_393 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c393
+ bl_0_393 br_0_393 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c393
+ bl_0_393 br_0_393 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c393
+ bl_0_393 br_0_393 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c393
+ bl_0_393 br_0_393 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c393
+ bl_0_393 br_0_393 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c393
+ bl_0_393 br_0_393 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c393
+ bl_0_393 br_0_393 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c393
+ bl_0_393 br_0_393 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c393
+ bl_0_393 br_0_393 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c394
+ bl_0_394 br_0_394 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c394
+ bl_0_394 br_0_394 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c394
+ bl_0_394 br_0_394 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c394
+ bl_0_394 br_0_394 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c394
+ bl_0_394 br_0_394 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c394
+ bl_0_394 br_0_394 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c394
+ bl_0_394 br_0_394 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c394
+ bl_0_394 br_0_394 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c394
+ bl_0_394 br_0_394 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c394
+ bl_0_394 br_0_394 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c394
+ bl_0_394 br_0_394 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c394
+ bl_0_394 br_0_394 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c394
+ bl_0_394 br_0_394 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c394
+ bl_0_394 br_0_394 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c394
+ bl_0_394 br_0_394 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c394
+ bl_0_394 br_0_394 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c394
+ bl_0_394 br_0_394 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c394
+ bl_0_394 br_0_394 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c394
+ bl_0_394 br_0_394 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c394
+ bl_0_394 br_0_394 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c394
+ bl_0_394 br_0_394 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c394
+ bl_0_394 br_0_394 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c394
+ bl_0_394 br_0_394 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c394
+ bl_0_394 br_0_394 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c394
+ bl_0_394 br_0_394 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c394
+ bl_0_394 br_0_394 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c394
+ bl_0_394 br_0_394 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c394
+ bl_0_394 br_0_394 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c394
+ bl_0_394 br_0_394 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c394
+ bl_0_394 br_0_394 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c394
+ bl_0_394 br_0_394 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c394
+ bl_0_394 br_0_394 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c394
+ bl_0_394 br_0_394 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c394
+ bl_0_394 br_0_394 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c394
+ bl_0_394 br_0_394 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c394
+ bl_0_394 br_0_394 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c394
+ bl_0_394 br_0_394 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c394
+ bl_0_394 br_0_394 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c394
+ bl_0_394 br_0_394 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c394
+ bl_0_394 br_0_394 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c394
+ bl_0_394 br_0_394 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c394
+ bl_0_394 br_0_394 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c394
+ bl_0_394 br_0_394 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c394
+ bl_0_394 br_0_394 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c394
+ bl_0_394 br_0_394 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c395
+ bl_0_395 br_0_395 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c395
+ bl_0_395 br_0_395 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c395
+ bl_0_395 br_0_395 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c395
+ bl_0_395 br_0_395 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c395
+ bl_0_395 br_0_395 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c395
+ bl_0_395 br_0_395 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c395
+ bl_0_395 br_0_395 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c395
+ bl_0_395 br_0_395 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c395
+ bl_0_395 br_0_395 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c395
+ bl_0_395 br_0_395 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c395
+ bl_0_395 br_0_395 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c395
+ bl_0_395 br_0_395 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c395
+ bl_0_395 br_0_395 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c395
+ bl_0_395 br_0_395 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c395
+ bl_0_395 br_0_395 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c395
+ bl_0_395 br_0_395 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c395
+ bl_0_395 br_0_395 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c395
+ bl_0_395 br_0_395 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c395
+ bl_0_395 br_0_395 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c395
+ bl_0_395 br_0_395 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c395
+ bl_0_395 br_0_395 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c395
+ bl_0_395 br_0_395 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c395
+ bl_0_395 br_0_395 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c395
+ bl_0_395 br_0_395 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c395
+ bl_0_395 br_0_395 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c395
+ bl_0_395 br_0_395 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c395
+ bl_0_395 br_0_395 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c395
+ bl_0_395 br_0_395 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c395
+ bl_0_395 br_0_395 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c395
+ bl_0_395 br_0_395 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c395
+ bl_0_395 br_0_395 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c395
+ bl_0_395 br_0_395 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c395
+ bl_0_395 br_0_395 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c395
+ bl_0_395 br_0_395 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c395
+ bl_0_395 br_0_395 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c395
+ bl_0_395 br_0_395 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c395
+ bl_0_395 br_0_395 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c395
+ bl_0_395 br_0_395 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c395
+ bl_0_395 br_0_395 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c395
+ bl_0_395 br_0_395 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c395
+ bl_0_395 br_0_395 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c395
+ bl_0_395 br_0_395 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c395
+ bl_0_395 br_0_395 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c395
+ bl_0_395 br_0_395 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c395
+ bl_0_395 br_0_395 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c396
+ bl_0_396 br_0_396 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c396
+ bl_0_396 br_0_396 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c396
+ bl_0_396 br_0_396 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c396
+ bl_0_396 br_0_396 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c396
+ bl_0_396 br_0_396 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c396
+ bl_0_396 br_0_396 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c396
+ bl_0_396 br_0_396 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c396
+ bl_0_396 br_0_396 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c396
+ bl_0_396 br_0_396 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c396
+ bl_0_396 br_0_396 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c396
+ bl_0_396 br_0_396 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c396
+ bl_0_396 br_0_396 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c396
+ bl_0_396 br_0_396 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c396
+ bl_0_396 br_0_396 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c396
+ bl_0_396 br_0_396 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c396
+ bl_0_396 br_0_396 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c396
+ bl_0_396 br_0_396 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c396
+ bl_0_396 br_0_396 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c396
+ bl_0_396 br_0_396 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c396
+ bl_0_396 br_0_396 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c396
+ bl_0_396 br_0_396 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c396
+ bl_0_396 br_0_396 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c396
+ bl_0_396 br_0_396 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c396
+ bl_0_396 br_0_396 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c396
+ bl_0_396 br_0_396 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c396
+ bl_0_396 br_0_396 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c396
+ bl_0_396 br_0_396 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c396
+ bl_0_396 br_0_396 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c396
+ bl_0_396 br_0_396 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c396
+ bl_0_396 br_0_396 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c396
+ bl_0_396 br_0_396 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c396
+ bl_0_396 br_0_396 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c396
+ bl_0_396 br_0_396 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c396
+ bl_0_396 br_0_396 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c396
+ bl_0_396 br_0_396 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c396
+ bl_0_396 br_0_396 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c396
+ bl_0_396 br_0_396 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c396
+ bl_0_396 br_0_396 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c396
+ bl_0_396 br_0_396 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c396
+ bl_0_396 br_0_396 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c396
+ bl_0_396 br_0_396 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c396
+ bl_0_396 br_0_396 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c396
+ bl_0_396 br_0_396 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c396
+ bl_0_396 br_0_396 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c396
+ bl_0_396 br_0_396 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c397
+ bl_0_397 br_0_397 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c397
+ bl_0_397 br_0_397 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c397
+ bl_0_397 br_0_397 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c397
+ bl_0_397 br_0_397 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c397
+ bl_0_397 br_0_397 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c397
+ bl_0_397 br_0_397 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c397
+ bl_0_397 br_0_397 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c397
+ bl_0_397 br_0_397 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c397
+ bl_0_397 br_0_397 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c397
+ bl_0_397 br_0_397 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c397
+ bl_0_397 br_0_397 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c397
+ bl_0_397 br_0_397 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c397
+ bl_0_397 br_0_397 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c397
+ bl_0_397 br_0_397 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c397
+ bl_0_397 br_0_397 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c397
+ bl_0_397 br_0_397 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c397
+ bl_0_397 br_0_397 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c397
+ bl_0_397 br_0_397 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c397
+ bl_0_397 br_0_397 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c397
+ bl_0_397 br_0_397 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c397
+ bl_0_397 br_0_397 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c397
+ bl_0_397 br_0_397 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c397
+ bl_0_397 br_0_397 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c397
+ bl_0_397 br_0_397 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c397
+ bl_0_397 br_0_397 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c397
+ bl_0_397 br_0_397 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c397
+ bl_0_397 br_0_397 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c397
+ bl_0_397 br_0_397 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c397
+ bl_0_397 br_0_397 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c397
+ bl_0_397 br_0_397 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c397
+ bl_0_397 br_0_397 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c397
+ bl_0_397 br_0_397 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c397
+ bl_0_397 br_0_397 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c397
+ bl_0_397 br_0_397 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c397
+ bl_0_397 br_0_397 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c397
+ bl_0_397 br_0_397 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c397
+ bl_0_397 br_0_397 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c397
+ bl_0_397 br_0_397 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c397
+ bl_0_397 br_0_397 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c397
+ bl_0_397 br_0_397 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c397
+ bl_0_397 br_0_397 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c397
+ bl_0_397 br_0_397 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c397
+ bl_0_397 br_0_397 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c397
+ bl_0_397 br_0_397 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c397
+ bl_0_397 br_0_397 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c398
+ bl_0_398 br_0_398 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c398
+ bl_0_398 br_0_398 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c398
+ bl_0_398 br_0_398 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c398
+ bl_0_398 br_0_398 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c398
+ bl_0_398 br_0_398 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c398
+ bl_0_398 br_0_398 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c398
+ bl_0_398 br_0_398 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c398
+ bl_0_398 br_0_398 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c398
+ bl_0_398 br_0_398 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c398
+ bl_0_398 br_0_398 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c398
+ bl_0_398 br_0_398 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c398
+ bl_0_398 br_0_398 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c398
+ bl_0_398 br_0_398 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c398
+ bl_0_398 br_0_398 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c398
+ bl_0_398 br_0_398 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c398
+ bl_0_398 br_0_398 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c398
+ bl_0_398 br_0_398 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c398
+ bl_0_398 br_0_398 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c398
+ bl_0_398 br_0_398 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c398
+ bl_0_398 br_0_398 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c398
+ bl_0_398 br_0_398 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c398
+ bl_0_398 br_0_398 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c398
+ bl_0_398 br_0_398 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c398
+ bl_0_398 br_0_398 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c398
+ bl_0_398 br_0_398 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c398
+ bl_0_398 br_0_398 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c398
+ bl_0_398 br_0_398 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c398
+ bl_0_398 br_0_398 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c398
+ bl_0_398 br_0_398 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c398
+ bl_0_398 br_0_398 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c398
+ bl_0_398 br_0_398 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c398
+ bl_0_398 br_0_398 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c398
+ bl_0_398 br_0_398 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c398
+ bl_0_398 br_0_398 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c398
+ bl_0_398 br_0_398 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c398
+ bl_0_398 br_0_398 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c398
+ bl_0_398 br_0_398 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c398
+ bl_0_398 br_0_398 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c398
+ bl_0_398 br_0_398 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c398
+ bl_0_398 br_0_398 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c398
+ bl_0_398 br_0_398 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c398
+ bl_0_398 br_0_398 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c398
+ bl_0_398 br_0_398 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c398
+ bl_0_398 br_0_398 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c398
+ bl_0_398 br_0_398 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c399
+ bl_0_399 br_0_399 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c399
+ bl_0_399 br_0_399 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c399
+ bl_0_399 br_0_399 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c399
+ bl_0_399 br_0_399 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c399
+ bl_0_399 br_0_399 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c399
+ bl_0_399 br_0_399 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c399
+ bl_0_399 br_0_399 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c399
+ bl_0_399 br_0_399 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c399
+ bl_0_399 br_0_399 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c399
+ bl_0_399 br_0_399 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c399
+ bl_0_399 br_0_399 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c399
+ bl_0_399 br_0_399 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c399
+ bl_0_399 br_0_399 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c399
+ bl_0_399 br_0_399 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c399
+ bl_0_399 br_0_399 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c399
+ bl_0_399 br_0_399 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c399
+ bl_0_399 br_0_399 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c399
+ bl_0_399 br_0_399 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c399
+ bl_0_399 br_0_399 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c399
+ bl_0_399 br_0_399 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c399
+ bl_0_399 br_0_399 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c399
+ bl_0_399 br_0_399 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c399
+ bl_0_399 br_0_399 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c399
+ bl_0_399 br_0_399 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c399
+ bl_0_399 br_0_399 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c399
+ bl_0_399 br_0_399 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c399
+ bl_0_399 br_0_399 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c399
+ bl_0_399 br_0_399 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c399
+ bl_0_399 br_0_399 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c399
+ bl_0_399 br_0_399 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c399
+ bl_0_399 br_0_399 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c399
+ bl_0_399 br_0_399 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c399
+ bl_0_399 br_0_399 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c399
+ bl_0_399 br_0_399 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c399
+ bl_0_399 br_0_399 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c399
+ bl_0_399 br_0_399 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c399
+ bl_0_399 br_0_399 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c399
+ bl_0_399 br_0_399 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c399
+ bl_0_399 br_0_399 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c399
+ bl_0_399 br_0_399 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c399
+ bl_0_399 br_0_399 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c399
+ bl_0_399 br_0_399 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c399
+ bl_0_399 br_0_399 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c399
+ bl_0_399 br_0_399 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c399
+ bl_0_399 br_0_399 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c400
+ bl_0_400 br_0_400 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c400
+ bl_0_400 br_0_400 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c400
+ bl_0_400 br_0_400 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c400
+ bl_0_400 br_0_400 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c400
+ bl_0_400 br_0_400 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c400
+ bl_0_400 br_0_400 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c400
+ bl_0_400 br_0_400 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c400
+ bl_0_400 br_0_400 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c400
+ bl_0_400 br_0_400 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c400
+ bl_0_400 br_0_400 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c400
+ bl_0_400 br_0_400 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c400
+ bl_0_400 br_0_400 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c400
+ bl_0_400 br_0_400 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c400
+ bl_0_400 br_0_400 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c400
+ bl_0_400 br_0_400 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c400
+ bl_0_400 br_0_400 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c400
+ bl_0_400 br_0_400 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c400
+ bl_0_400 br_0_400 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c400
+ bl_0_400 br_0_400 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c400
+ bl_0_400 br_0_400 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c400
+ bl_0_400 br_0_400 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c400
+ bl_0_400 br_0_400 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c400
+ bl_0_400 br_0_400 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c400
+ bl_0_400 br_0_400 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c400
+ bl_0_400 br_0_400 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c400
+ bl_0_400 br_0_400 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c400
+ bl_0_400 br_0_400 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c400
+ bl_0_400 br_0_400 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c400
+ bl_0_400 br_0_400 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c400
+ bl_0_400 br_0_400 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c400
+ bl_0_400 br_0_400 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c400
+ bl_0_400 br_0_400 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c400
+ bl_0_400 br_0_400 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c400
+ bl_0_400 br_0_400 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c400
+ bl_0_400 br_0_400 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c400
+ bl_0_400 br_0_400 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c400
+ bl_0_400 br_0_400 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c400
+ bl_0_400 br_0_400 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c400
+ bl_0_400 br_0_400 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c400
+ bl_0_400 br_0_400 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c400
+ bl_0_400 br_0_400 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c400
+ bl_0_400 br_0_400 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c400
+ bl_0_400 br_0_400 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c400
+ bl_0_400 br_0_400 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c400
+ bl_0_400 br_0_400 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c401
+ bl_0_401 br_0_401 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c401
+ bl_0_401 br_0_401 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c401
+ bl_0_401 br_0_401 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c401
+ bl_0_401 br_0_401 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c401
+ bl_0_401 br_0_401 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c401
+ bl_0_401 br_0_401 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c401
+ bl_0_401 br_0_401 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c401
+ bl_0_401 br_0_401 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c401
+ bl_0_401 br_0_401 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c401
+ bl_0_401 br_0_401 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c401
+ bl_0_401 br_0_401 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c401
+ bl_0_401 br_0_401 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c401
+ bl_0_401 br_0_401 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c401
+ bl_0_401 br_0_401 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c401
+ bl_0_401 br_0_401 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c401
+ bl_0_401 br_0_401 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c401
+ bl_0_401 br_0_401 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c401
+ bl_0_401 br_0_401 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c401
+ bl_0_401 br_0_401 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c401
+ bl_0_401 br_0_401 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c401
+ bl_0_401 br_0_401 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c401
+ bl_0_401 br_0_401 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c401
+ bl_0_401 br_0_401 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c401
+ bl_0_401 br_0_401 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c401
+ bl_0_401 br_0_401 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c401
+ bl_0_401 br_0_401 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c401
+ bl_0_401 br_0_401 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c401
+ bl_0_401 br_0_401 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c401
+ bl_0_401 br_0_401 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c401
+ bl_0_401 br_0_401 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c401
+ bl_0_401 br_0_401 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c401
+ bl_0_401 br_0_401 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c401
+ bl_0_401 br_0_401 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c401
+ bl_0_401 br_0_401 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c401
+ bl_0_401 br_0_401 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c401
+ bl_0_401 br_0_401 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c401
+ bl_0_401 br_0_401 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c401
+ bl_0_401 br_0_401 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c401
+ bl_0_401 br_0_401 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c401
+ bl_0_401 br_0_401 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c401
+ bl_0_401 br_0_401 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c401
+ bl_0_401 br_0_401 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c401
+ bl_0_401 br_0_401 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c401
+ bl_0_401 br_0_401 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c401
+ bl_0_401 br_0_401 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c402
+ bl_0_402 br_0_402 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c402
+ bl_0_402 br_0_402 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c402
+ bl_0_402 br_0_402 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c402
+ bl_0_402 br_0_402 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c402
+ bl_0_402 br_0_402 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c402
+ bl_0_402 br_0_402 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c402
+ bl_0_402 br_0_402 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c402
+ bl_0_402 br_0_402 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c402
+ bl_0_402 br_0_402 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c402
+ bl_0_402 br_0_402 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c402
+ bl_0_402 br_0_402 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c402
+ bl_0_402 br_0_402 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c402
+ bl_0_402 br_0_402 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c402
+ bl_0_402 br_0_402 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c402
+ bl_0_402 br_0_402 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c402
+ bl_0_402 br_0_402 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c402
+ bl_0_402 br_0_402 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c402
+ bl_0_402 br_0_402 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c402
+ bl_0_402 br_0_402 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c402
+ bl_0_402 br_0_402 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c402
+ bl_0_402 br_0_402 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c402
+ bl_0_402 br_0_402 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c402
+ bl_0_402 br_0_402 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c402
+ bl_0_402 br_0_402 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c402
+ bl_0_402 br_0_402 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c402
+ bl_0_402 br_0_402 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c402
+ bl_0_402 br_0_402 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c402
+ bl_0_402 br_0_402 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c402
+ bl_0_402 br_0_402 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c402
+ bl_0_402 br_0_402 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c402
+ bl_0_402 br_0_402 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c402
+ bl_0_402 br_0_402 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c402
+ bl_0_402 br_0_402 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c402
+ bl_0_402 br_0_402 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c402
+ bl_0_402 br_0_402 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c402
+ bl_0_402 br_0_402 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c402
+ bl_0_402 br_0_402 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c402
+ bl_0_402 br_0_402 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c402
+ bl_0_402 br_0_402 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c402
+ bl_0_402 br_0_402 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c402
+ bl_0_402 br_0_402 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c402
+ bl_0_402 br_0_402 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c402
+ bl_0_402 br_0_402 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c402
+ bl_0_402 br_0_402 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c402
+ bl_0_402 br_0_402 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c403
+ bl_0_403 br_0_403 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c403
+ bl_0_403 br_0_403 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c403
+ bl_0_403 br_0_403 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c403
+ bl_0_403 br_0_403 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c403
+ bl_0_403 br_0_403 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c403
+ bl_0_403 br_0_403 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c403
+ bl_0_403 br_0_403 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c403
+ bl_0_403 br_0_403 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c403
+ bl_0_403 br_0_403 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c403
+ bl_0_403 br_0_403 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c403
+ bl_0_403 br_0_403 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c403
+ bl_0_403 br_0_403 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c403
+ bl_0_403 br_0_403 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c403
+ bl_0_403 br_0_403 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c403
+ bl_0_403 br_0_403 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c403
+ bl_0_403 br_0_403 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c403
+ bl_0_403 br_0_403 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c403
+ bl_0_403 br_0_403 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c403
+ bl_0_403 br_0_403 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c403
+ bl_0_403 br_0_403 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c403
+ bl_0_403 br_0_403 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c403
+ bl_0_403 br_0_403 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c403
+ bl_0_403 br_0_403 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c403
+ bl_0_403 br_0_403 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c403
+ bl_0_403 br_0_403 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c403
+ bl_0_403 br_0_403 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c403
+ bl_0_403 br_0_403 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c403
+ bl_0_403 br_0_403 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c403
+ bl_0_403 br_0_403 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c403
+ bl_0_403 br_0_403 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c403
+ bl_0_403 br_0_403 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c403
+ bl_0_403 br_0_403 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c403
+ bl_0_403 br_0_403 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c403
+ bl_0_403 br_0_403 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c403
+ bl_0_403 br_0_403 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c403
+ bl_0_403 br_0_403 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c403
+ bl_0_403 br_0_403 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c403
+ bl_0_403 br_0_403 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c403
+ bl_0_403 br_0_403 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c403
+ bl_0_403 br_0_403 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c403
+ bl_0_403 br_0_403 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c403
+ bl_0_403 br_0_403 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c403
+ bl_0_403 br_0_403 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c403
+ bl_0_403 br_0_403 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c403
+ bl_0_403 br_0_403 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c404
+ bl_0_404 br_0_404 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c404
+ bl_0_404 br_0_404 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c404
+ bl_0_404 br_0_404 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c404
+ bl_0_404 br_0_404 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c404
+ bl_0_404 br_0_404 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c404
+ bl_0_404 br_0_404 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c404
+ bl_0_404 br_0_404 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c404
+ bl_0_404 br_0_404 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c404
+ bl_0_404 br_0_404 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c404
+ bl_0_404 br_0_404 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c404
+ bl_0_404 br_0_404 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c404
+ bl_0_404 br_0_404 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c404
+ bl_0_404 br_0_404 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c404
+ bl_0_404 br_0_404 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c404
+ bl_0_404 br_0_404 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c404
+ bl_0_404 br_0_404 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c404
+ bl_0_404 br_0_404 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c404
+ bl_0_404 br_0_404 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c404
+ bl_0_404 br_0_404 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c404
+ bl_0_404 br_0_404 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c404
+ bl_0_404 br_0_404 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c404
+ bl_0_404 br_0_404 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c404
+ bl_0_404 br_0_404 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c404
+ bl_0_404 br_0_404 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c404
+ bl_0_404 br_0_404 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c404
+ bl_0_404 br_0_404 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c404
+ bl_0_404 br_0_404 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c404
+ bl_0_404 br_0_404 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c404
+ bl_0_404 br_0_404 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c404
+ bl_0_404 br_0_404 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c404
+ bl_0_404 br_0_404 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c404
+ bl_0_404 br_0_404 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c404
+ bl_0_404 br_0_404 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c404
+ bl_0_404 br_0_404 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c404
+ bl_0_404 br_0_404 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c404
+ bl_0_404 br_0_404 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c404
+ bl_0_404 br_0_404 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c404
+ bl_0_404 br_0_404 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c404
+ bl_0_404 br_0_404 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c404
+ bl_0_404 br_0_404 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c404
+ bl_0_404 br_0_404 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c404
+ bl_0_404 br_0_404 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c404
+ bl_0_404 br_0_404 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c404
+ bl_0_404 br_0_404 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c404
+ bl_0_404 br_0_404 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c405
+ bl_0_405 br_0_405 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c405
+ bl_0_405 br_0_405 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c405
+ bl_0_405 br_0_405 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c405
+ bl_0_405 br_0_405 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c405
+ bl_0_405 br_0_405 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c405
+ bl_0_405 br_0_405 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c405
+ bl_0_405 br_0_405 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c405
+ bl_0_405 br_0_405 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c405
+ bl_0_405 br_0_405 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c405
+ bl_0_405 br_0_405 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c405
+ bl_0_405 br_0_405 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c405
+ bl_0_405 br_0_405 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c405
+ bl_0_405 br_0_405 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c405
+ bl_0_405 br_0_405 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c405
+ bl_0_405 br_0_405 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c405
+ bl_0_405 br_0_405 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c405
+ bl_0_405 br_0_405 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c405
+ bl_0_405 br_0_405 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c405
+ bl_0_405 br_0_405 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c405
+ bl_0_405 br_0_405 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c405
+ bl_0_405 br_0_405 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c405
+ bl_0_405 br_0_405 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c405
+ bl_0_405 br_0_405 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c405
+ bl_0_405 br_0_405 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c405
+ bl_0_405 br_0_405 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c405
+ bl_0_405 br_0_405 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c405
+ bl_0_405 br_0_405 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c405
+ bl_0_405 br_0_405 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c405
+ bl_0_405 br_0_405 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c405
+ bl_0_405 br_0_405 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c405
+ bl_0_405 br_0_405 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c405
+ bl_0_405 br_0_405 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c405
+ bl_0_405 br_0_405 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c405
+ bl_0_405 br_0_405 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c405
+ bl_0_405 br_0_405 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c405
+ bl_0_405 br_0_405 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c405
+ bl_0_405 br_0_405 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c405
+ bl_0_405 br_0_405 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c405
+ bl_0_405 br_0_405 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c405
+ bl_0_405 br_0_405 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c405
+ bl_0_405 br_0_405 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c405
+ bl_0_405 br_0_405 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c405
+ bl_0_405 br_0_405 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c405
+ bl_0_405 br_0_405 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c405
+ bl_0_405 br_0_405 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c406
+ bl_0_406 br_0_406 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c406
+ bl_0_406 br_0_406 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c406
+ bl_0_406 br_0_406 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c406
+ bl_0_406 br_0_406 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c406
+ bl_0_406 br_0_406 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c406
+ bl_0_406 br_0_406 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c406
+ bl_0_406 br_0_406 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c406
+ bl_0_406 br_0_406 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c406
+ bl_0_406 br_0_406 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c406
+ bl_0_406 br_0_406 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c406
+ bl_0_406 br_0_406 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c406
+ bl_0_406 br_0_406 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c406
+ bl_0_406 br_0_406 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c406
+ bl_0_406 br_0_406 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c406
+ bl_0_406 br_0_406 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c406
+ bl_0_406 br_0_406 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c406
+ bl_0_406 br_0_406 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c406
+ bl_0_406 br_0_406 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c406
+ bl_0_406 br_0_406 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c406
+ bl_0_406 br_0_406 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c406
+ bl_0_406 br_0_406 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c406
+ bl_0_406 br_0_406 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c406
+ bl_0_406 br_0_406 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c406
+ bl_0_406 br_0_406 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c406
+ bl_0_406 br_0_406 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c406
+ bl_0_406 br_0_406 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c406
+ bl_0_406 br_0_406 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c406
+ bl_0_406 br_0_406 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c406
+ bl_0_406 br_0_406 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c406
+ bl_0_406 br_0_406 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c406
+ bl_0_406 br_0_406 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c406
+ bl_0_406 br_0_406 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c406
+ bl_0_406 br_0_406 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c406
+ bl_0_406 br_0_406 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c406
+ bl_0_406 br_0_406 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c406
+ bl_0_406 br_0_406 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c406
+ bl_0_406 br_0_406 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c406
+ bl_0_406 br_0_406 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c406
+ bl_0_406 br_0_406 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c406
+ bl_0_406 br_0_406 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c406
+ bl_0_406 br_0_406 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c406
+ bl_0_406 br_0_406 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c406
+ bl_0_406 br_0_406 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c406
+ bl_0_406 br_0_406 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c406
+ bl_0_406 br_0_406 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c407
+ bl_0_407 br_0_407 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c407
+ bl_0_407 br_0_407 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c407
+ bl_0_407 br_0_407 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c407
+ bl_0_407 br_0_407 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c407
+ bl_0_407 br_0_407 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c407
+ bl_0_407 br_0_407 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c407
+ bl_0_407 br_0_407 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c407
+ bl_0_407 br_0_407 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c407
+ bl_0_407 br_0_407 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c407
+ bl_0_407 br_0_407 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c407
+ bl_0_407 br_0_407 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c407
+ bl_0_407 br_0_407 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c407
+ bl_0_407 br_0_407 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c407
+ bl_0_407 br_0_407 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c407
+ bl_0_407 br_0_407 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c407
+ bl_0_407 br_0_407 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c407
+ bl_0_407 br_0_407 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c407
+ bl_0_407 br_0_407 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c407
+ bl_0_407 br_0_407 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c407
+ bl_0_407 br_0_407 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c407
+ bl_0_407 br_0_407 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c407
+ bl_0_407 br_0_407 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c407
+ bl_0_407 br_0_407 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c407
+ bl_0_407 br_0_407 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c407
+ bl_0_407 br_0_407 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c407
+ bl_0_407 br_0_407 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c407
+ bl_0_407 br_0_407 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c407
+ bl_0_407 br_0_407 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c407
+ bl_0_407 br_0_407 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c407
+ bl_0_407 br_0_407 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c407
+ bl_0_407 br_0_407 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c407
+ bl_0_407 br_0_407 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c407
+ bl_0_407 br_0_407 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c407
+ bl_0_407 br_0_407 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c407
+ bl_0_407 br_0_407 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c407
+ bl_0_407 br_0_407 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c407
+ bl_0_407 br_0_407 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c407
+ bl_0_407 br_0_407 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c407
+ bl_0_407 br_0_407 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c407
+ bl_0_407 br_0_407 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c407
+ bl_0_407 br_0_407 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c407
+ bl_0_407 br_0_407 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c407
+ bl_0_407 br_0_407 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c407
+ bl_0_407 br_0_407 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c407
+ bl_0_407 br_0_407 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c408
+ bl_0_408 br_0_408 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c408
+ bl_0_408 br_0_408 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c408
+ bl_0_408 br_0_408 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c408
+ bl_0_408 br_0_408 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c408
+ bl_0_408 br_0_408 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c408
+ bl_0_408 br_0_408 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c408
+ bl_0_408 br_0_408 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c408
+ bl_0_408 br_0_408 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c408
+ bl_0_408 br_0_408 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c408
+ bl_0_408 br_0_408 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c408
+ bl_0_408 br_0_408 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c408
+ bl_0_408 br_0_408 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c408
+ bl_0_408 br_0_408 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c408
+ bl_0_408 br_0_408 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c408
+ bl_0_408 br_0_408 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c408
+ bl_0_408 br_0_408 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c408
+ bl_0_408 br_0_408 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c408
+ bl_0_408 br_0_408 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c408
+ bl_0_408 br_0_408 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c408
+ bl_0_408 br_0_408 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c408
+ bl_0_408 br_0_408 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c408
+ bl_0_408 br_0_408 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c408
+ bl_0_408 br_0_408 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c408
+ bl_0_408 br_0_408 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c408
+ bl_0_408 br_0_408 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c408
+ bl_0_408 br_0_408 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c408
+ bl_0_408 br_0_408 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c408
+ bl_0_408 br_0_408 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c408
+ bl_0_408 br_0_408 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c408
+ bl_0_408 br_0_408 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c408
+ bl_0_408 br_0_408 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c408
+ bl_0_408 br_0_408 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c408
+ bl_0_408 br_0_408 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c408
+ bl_0_408 br_0_408 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c408
+ bl_0_408 br_0_408 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c408
+ bl_0_408 br_0_408 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c408
+ bl_0_408 br_0_408 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c408
+ bl_0_408 br_0_408 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c408
+ bl_0_408 br_0_408 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c408
+ bl_0_408 br_0_408 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c408
+ bl_0_408 br_0_408 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c408
+ bl_0_408 br_0_408 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c408
+ bl_0_408 br_0_408 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c408
+ bl_0_408 br_0_408 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c408
+ bl_0_408 br_0_408 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c409
+ bl_0_409 br_0_409 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c409
+ bl_0_409 br_0_409 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c409
+ bl_0_409 br_0_409 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c409
+ bl_0_409 br_0_409 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c409
+ bl_0_409 br_0_409 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c409
+ bl_0_409 br_0_409 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c409
+ bl_0_409 br_0_409 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c409
+ bl_0_409 br_0_409 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c409
+ bl_0_409 br_0_409 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c409
+ bl_0_409 br_0_409 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c409
+ bl_0_409 br_0_409 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c409
+ bl_0_409 br_0_409 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c409
+ bl_0_409 br_0_409 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c409
+ bl_0_409 br_0_409 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c409
+ bl_0_409 br_0_409 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c409
+ bl_0_409 br_0_409 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c409
+ bl_0_409 br_0_409 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c409
+ bl_0_409 br_0_409 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c409
+ bl_0_409 br_0_409 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c409
+ bl_0_409 br_0_409 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c409
+ bl_0_409 br_0_409 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c409
+ bl_0_409 br_0_409 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c409
+ bl_0_409 br_0_409 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c409
+ bl_0_409 br_0_409 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c409
+ bl_0_409 br_0_409 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c409
+ bl_0_409 br_0_409 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c409
+ bl_0_409 br_0_409 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c409
+ bl_0_409 br_0_409 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c409
+ bl_0_409 br_0_409 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c409
+ bl_0_409 br_0_409 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c409
+ bl_0_409 br_0_409 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c409
+ bl_0_409 br_0_409 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c409
+ bl_0_409 br_0_409 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c409
+ bl_0_409 br_0_409 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c409
+ bl_0_409 br_0_409 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c409
+ bl_0_409 br_0_409 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c409
+ bl_0_409 br_0_409 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c409
+ bl_0_409 br_0_409 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c409
+ bl_0_409 br_0_409 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c409
+ bl_0_409 br_0_409 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c409
+ bl_0_409 br_0_409 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c409
+ bl_0_409 br_0_409 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c409
+ bl_0_409 br_0_409 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c409
+ bl_0_409 br_0_409 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c409
+ bl_0_409 br_0_409 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c410
+ bl_0_410 br_0_410 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c410
+ bl_0_410 br_0_410 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c410
+ bl_0_410 br_0_410 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c410
+ bl_0_410 br_0_410 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c410
+ bl_0_410 br_0_410 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c410
+ bl_0_410 br_0_410 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c410
+ bl_0_410 br_0_410 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c410
+ bl_0_410 br_0_410 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c410
+ bl_0_410 br_0_410 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c410
+ bl_0_410 br_0_410 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c410
+ bl_0_410 br_0_410 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c410
+ bl_0_410 br_0_410 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c410
+ bl_0_410 br_0_410 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c410
+ bl_0_410 br_0_410 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c410
+ bl_0_410 br_0_410 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c410
+ bl_0_410 br_0_410 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c410
+ bl_0_410 br_0_410 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c410
+ bl_0_410 br_0_410 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c410
+ bl_0_410 br_0_410 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c410
+ bl_0_410 br_0_410 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c410
+ bl_0_410 br_0_410 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c410
+ bl_0_410 br_0_410 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c410
+ bl_0_410 br_0_410 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c410
+ bl_0_410 br_0_410 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c410
+ bl_0_410 br_0_410 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c410
+ bl_0_410 br_0_410 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c410
+ bl_0_410 br_0_410 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c410
+ bl_0_410 br_0_410 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c410
+ bl_0_410 br_0_410 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c410
+ bl_0_410 br_0_410 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c410
+ bl_0_410 br_0_410 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c410
+ bl_0_410 br_0_410 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c410
+ bl_0_410 br_0_410 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c410
+ bl_0_410 br_0_410 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c410
+ bl_0_410 br_0_410 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c410
+ bl_0_410 br_0_410 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c410
+ bl_0_410 br_0_410 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c410
+ bl_0_410 br_0_410 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c410
+ bl_0_410 br_0_410 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c410
+ bl_0_410 br_0_410 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c410
+ bl_0_410 br_0_410 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c410
+ bl_0_410 br_0_410 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c410
+ bl_0_410 br_0_410 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c410
+ bl_0_410 br_0_410 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c410
+ bl_0_410 br_0_410 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c411
+ bl_0_411 br_0_411 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c411
+ bl_0_411 br_0_411 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c411
+ bl_0_411 br_0_411 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c411
+ bl_0_411 br_0_411 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c411
+ bl_0_411 br_0_411 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c411
+ bl_0_411 br_0_411 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c411
+ bl_0_411 br_0_411 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c411
+ bl_0_411 br_0_411 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c411
+ bl_0_411 br_0_411 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c411
+ bl_0_411 br_0_411 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c411
+ bl_0_411 br_0_411 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c411
+ bl_0_411 br_0_411 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c411
+ bl_0_411 br_0_411 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c411
+ bl_0_411 br_0_411 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c411
+ bl_0_411 br_0_411 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c411
+ bl_0_411 br_0_411 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c411
+ bl_0_411 br_0_411 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c411
+ bl_0_411 br_0_411 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c411
+ bl_0_411 br_0_411 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c411
+ bl_0_411 br_0_411 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c411
+ bl_0_411 br_0_411 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c411
+ bl_0_411 br_0_411 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c411
+ bl_0_411 br_0_411 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c411
+ bl_0_411 br_0_411 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c411
+ bl_0_411 br_0_411 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c411
+ bl_0_411 br_0_411 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c411
+ bl_0_411 br_0_411 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c411
+ bl_0_411 br_0_411 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c411
+ bl_0_411 br_0_411 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c411
+ bl_0_411 br_0_411 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c411
+ bl_0_411 br_0_411 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c411
+ bl_0_411 br_0_411 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c411
+ bl_0_411 br_0_411 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c411
+ bl_0_411 br_0_411 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c411
+ bl_0_411 br_0_411 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c411
+ bl_0_411 br_0_411 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c411
+ bl_0_411 br_0_411 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c411
+ bl_0_411 br_0_411 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c411
+ bl_0_411 br_0_411 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c411
+ bl_0_411 br_0_411 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c411
+ bl_0_411 br_0_411 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c411
+ bl_0_411 br_0_411 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c411
+ bl_0_411 br_0_411 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c411
+ bl_0_411 br_0_411 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c411
+ bl_0_411 br_0_411 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c412
+ bl_0_412 br_0_412 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c412
+ bl_0_412 br_0_412 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c412
+ bl_0_412 br_0_412 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c412
+ bl_0_412 br_0_412 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c412
+ bl_0_412 br_0_412 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c412
+ bl_0_412 br_0_412 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c412
+ bl_0_412 br_0_412 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c412
+ bl_0_412 br_0_412 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c412
+ bl_0_412 br_0_412 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c412
+ bl_0_412 br_0_412 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c412
+ bl_0_412 br_0_412 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c412
+ bl_0_412 br_0_412 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c412
+ bl_0_412 br_0_412 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c412
+ bl_0_412 br_0_412 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c412
+ bl_0_412 br_0_412 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c412
+ bl_0_412 br_0_412 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c412
+ bl_0_412 br_0_412 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c412
+ bl_0_412 br_0_412 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c412
+ bl_0_412 br_0_412 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c412
+ bl_0_412 br_0_412 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c412
+ bl_0_412 br_0_412 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c412
+ bl_0_412 br_0_412 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c412
+ bl_0_412 br_0_412 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c412
+ bl_0_412 br_0_412 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c412
+ bl_0_412 br_0_412 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c412
+ bl_0_412 br_0_412 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c412
+ bl_0_412 br_0_412 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c412
+ bl_0_412 br_0_412 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c412
+ bl_0_412 br_0_412 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c412
+ bl_0_412 br_0_412 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c412
+ bl_0_412 br_0_412 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c412
+ bl_0_412 br_0_412 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c412
+ bl_0_412 br_0_412 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c412
+ bl_0_412 br_0_412 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c412
+ bl_0_412 br_0_412 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c412
+ bl_0_412 br_0_412 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c412
+ bl_0_412 br_0_412 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c412
+ bl_0_412 br_0_412 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c412
+ bl_0_412 br_0_412 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c412
+ bl_0_412 br_0_412 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c412
+ bl_0_412 br_0_412 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c412
+ bl_0_412 br_0_412 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c412
+ bl_0_412 br_0_412 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c412
+ bl_0_412 br_0_412 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c412
+ bl_0_412 br_0_412 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c413
+ bl_0_413 br_0_413 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c413
+ bl_0_413 br_0_413 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c413
+ bl_0_413 br_0_413 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c413
+ bl_0_413 br_0_413 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c413
+ bl_0_413 br_0_413 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c413
+ bl_0_413 br_0_413 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c413
+ bl_0_413 br_0_413 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c413
+ bl_0_413 br_0_413 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c413
+ bl_0_413 br_0_413 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c413
+ bl_0_413 br_0_413 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c413
+ bl_0_413 br_0_413 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c413
+ bl_0_413 br_0_413 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c413
+ bl_0_413 br_0_413 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c413
+ bl_0_413 br_0_413 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c413
+ bl_0_413 br_0_413 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c413
+ bl_0_413 br_0_413 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c413
+ bl_0_413 br_0_413 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c413
+ bl_0_413 br_0_413 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c413
+ bl_0_413 br_0_413 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c413
+ bl_0_413 br_0_413 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c413
+ bl_0_413 br_0_413 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c413
+ bl_0_413 br_0_413 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c413
+ bl_0_413 br_0_413 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c413
+ bl_0_413 br_0_413 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c413
+ bl_0_413 br_0_413 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c413
+ bl_0_413 br_0_413 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c413
+ bl_0_413 br_0_413 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c413
+ bl_0_413 br_0_413 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c413
+ bl_0_413 br_0_413 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c413
+ bl_0_413 br_0_413 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c413
+ bl_0_413 br_0_413 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c413
+ bl_0_413 br_0_413 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c413
+ bl_0_413 br_0_413 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c413
+ bl_0_413 br_0_413 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c413
+ bl_0_413 br_0_413 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c413
+ bl_0_413 br_0_413 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c413
+ bl_0_413 br_0_413 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c413
+ bl_0_413 br_0_413 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c413
+ bl_0_413 br_0_413 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c413
+ bl_0_413 br_0_413 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c413
+ bl_0_413 br_0_413 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c413
+ bl_0_413 br_0_413 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c413
+ bl_0_413 br_0_413 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c413
+ bl_0_413 br_0_413 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c413
+ bl_0_413 br_0_413 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c414
+ bl_0_414 br_0_414 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c414
+ bl_0_414 br_0_414 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c414
+ bl_0_414 br_0_414 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c414
+ bl_0_414 br_0_414 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c414
+ bl_0_414 br_0_414 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c414
+ bl_0_414 br_0_414 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c414
+ bl_0_414 br_0_414 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c414
+ bl_0_414 br_0_414 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c414
+ bl_0_414 br_0_414 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c414
+ bl_0_414 br_0_414 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c414
+ bl_0_414 br_0_414 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c414
+ bl_0_414 br_0_414 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c414
+ bl_0_414 br_0_414 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c414
+ bl_0_414 br_0_414 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c414
+ bl_0_414 br_0_414 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c414
+ bl_0_414 br_0_414 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c414
+ bl_0_414 br_0_414 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c414
+ bl_0_414 br_0_414 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c414
+ bl_0_414 br_0_414 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c414
+ bl_0_414 br_0_414 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c414
+ bl_0_414 br_0_414 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c414
+ bl_0_414 br_0_414 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c414
+ bl_0_414 br_0_414 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c414
+ bl_0_414 br_0_414 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c414
+ bl_0_414 br_0_414 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c414
+ bl_0_414 br_0_414 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c414
+ bl_0_414 br_0_414 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c414
+ bl_0_414 br_0_414 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c414
+ bl_0_414 br_0_414 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c414
+ bl_0_414 br_0_414 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c414
+ bl_0_414 br_0_414 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c414
+ bl_0_414 br_0_414 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c414
+ bl_0_414 br_0_414 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c414
+ bl_0_414 br_0_414 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c414
+ bl_0_414 br_0_414 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c414
+ bl_0_414 br_0_414 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c414
+ bl_0_414 br_0_414 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c414
+ bl_0_414 br_0_414 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c414
+ bl_0_414 br_0_414 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c414
+ bl_0_414 br_0_414 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c414
+ bl_0_414 br_0_414 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c414
+ bl_0_414 br_0_414 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c414
+ bl_0_414 br_0_414 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c414
+ bl_0_414 br_0_414 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c414
+ bl_0_414 br_0_414 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c415
+ bl_0_415 br_0_415 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c415
+ bl_0_415 br_0_415 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c415
+ bl_0_415 br_0_415 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c415
+ bl_0_415 br_0_415 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c415
+ bl_0_415 br_0_415 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c415
+ bl_0_415 br_0_415 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c415
+ bl_0_415 br_0_415 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c415
+ bl_0_415 br_0_415 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c415
+ bl_0_415 br_0_415 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c415
+ bl_0_415 br_0_415 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c415
+ bl_0_415 br_0_415 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c415
+ bl_0_415 br_0_415 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c415
+ bl_0_415 br_0_415 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c415
+ bl_0_415 br_0_415 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c415
+ bl_0_415 br_0_415 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c415
+ bl_0_415 br_0_415 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c415
+ bl_0_415 br_0_415 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c415
+ bl_0_415 br_0_415 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c415
+ bl_0_415 br_0_415 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c415
+ bl_0_415 br_0_415 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c415
+ bl_0_415 br_0_415 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c415
+ bl_0_415 br_0_415 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c415
+ bl_0_415 br_0_415 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c415
+ bl_0_415 br_0_415 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c415
+ bl_0_415 br_0_415 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c415
+ bl_0_415 br_0_415 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c415
+ bl_0_415 br_0_415 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c415
+ bl_0_415 br_0_415 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c415
+ bl_0_415 br_0_415 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c415
+ bl_0_415 br_0_415 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c415
+ bl_0_415 br_0_415 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c415
+ bl_0_415 br_0_415 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c415
+ bl_0_415 br_0_415 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c415
+ bl_0_415 br_0_415 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c415
+ bl_0_415 br_0_415 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c415
+ bl_0_415 br_0_415 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c415
+ bl_0_415 br_0_415 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c415
+ bl_0_415 br_0_415 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c415
+ bl_0_415 br_0_415 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c415
+ bl_0_415 br_0_415 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c415
+ bl_0_415 br_0_415 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c415
+ bl_0_415 br_0_415 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c415
+ bl_0_415 br_0_415 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c415
+ bl_0_415 br_0_415 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c415
+ bl_0_415 br_0_415 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c416
+ bl_0_416 br_0_416 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c416
+ bl_0_416 br_0_416 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c416
+ bl_0_416 br_0_416 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c416
+ bl_0_416 br_0_416 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c416
+ bl_0_416 br_0_416 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c416
+ bl_0_416 br_0_416 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c416
+ bl_0_416 br_0_416 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c416
+ bl_0_416 br_0_416 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c416
+ bl_0_416 br_0_416 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c416
+ bl_0_416 br_0_416 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c416
+ bl_0_416 br_0_416 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c416
+ bl_0_416 br_0_416 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c416
+ bl_0_416 br_0_416 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c416
+ bl_0_416 br_0_416 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c416
+ bl_0_416 br_0_416 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c416
+ bl_0_416 br_0_416 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c416
+ bl_0_416 br_0_416 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c416
+ bl_0_416 br_0_416 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c416
+ bl_0_416 br_0_416 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c416
+ bl_0_416 br_0_416 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c416
+ bl_0_416 br_0_416 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c416
+ bl_0_416 br_0_416 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c416
+ bl_0_416 br_0_416 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c416
+ bl_0_416 br_0_416 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c416
+ bl_0_416 br_0_416 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c416
+ bl_0_416 br_0_416 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c416
+ bl_0_416 br_0_416 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c416
+ bl_0_416 br_0_416 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c416
+ bl_0_416 br_0_416 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c416
+ bl_0_416 br_0_416 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c416
+ bl_0_416 br_0_416 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c416
+ bl_0_416 br_0_416 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c416
+ bl_0_416 br_0_416 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c416
+ bl_0_416 br_0_416 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c416
+ bl_0_416 br_0_416 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c416
+ bl_0_416 br_0_416 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c416
+ bl_0_416 br_0_416 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c416
+ bl_0_416 br_0_416 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c416
+ bl_0_416 br_0_416 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c416
+ bl_0_416 br_0_416 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c416
+ bl_0_416 br_0_416 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c416
+ bl_0_416 br_0_416 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c416
+ bl_0_416 br_0_416 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c416
+ bl_0_416 br_0_416 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c416
+ bl_0_416 br_0_416 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c417
+ bl_0_417 br_0_417 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c417
+ bl_0_417 br_0_417 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c417
+ bl_0_417 br_0_417 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c417
+ bl_0_417 br_0_417 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c417
+ bl_0_417 br_0_417 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c417
+ bl_0_417 br_0_417 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c417
+ bl_0_417 br_0_417 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c417
+ bl_0_417 br_0_417 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c417
+ bl_0_417 br_0_417 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c417
+ bl_0_417 br_0_417 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c417
+ bl_0_417 br_0_417 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c417
+ bl_0_417 br_0_417 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c417
+ bl_0_417 br_0_417 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c417
+ bl_0_417 br_0_417 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c417
+ bl_0_417 br_0_417 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c417
+ bl_0_417 br_0_417 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c417
+ bl_0_417 br_0_417 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c417
+ bl_0_417 br_0_417 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c417
+ bl_0_417 br_0_417 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c417
+ bl_0_417 br_0_417 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c417
+ bl_0_417 br_0_417 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c417
+ bl_0_417 br_0_417 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c417
+ bl_0_417 br_0_417 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c417
+ bl_0_417 br_0_417 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c417
+ bl_0_417 br_0_417 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c417
+ bl_0_417 br_0_417 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c417
+ bl_0_417 br_0_417 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c417
+ bl_0_417 br_0_417 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c417
+ bl_0_417 br_0_417 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c417
+ bl_0_417 br_0_417 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c417
+ bl_0_417 br_0_417 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c417
+ bl_0_417 br_0_417 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c417
+ bl_0_417 br_0_417 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c417
+ bl_0_417 br_0_417 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c417
+ bl_0_417 br_0_417 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c417
+ bl_0_417 br_0_417 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c417
+ bl_0_417 br_0_417 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c417
+ bl_0_417 br_0_417 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c417
+ bl_0_417 br_0_417 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c417
+ bl_0_417 br_0_417 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c417
+ bl_0_417 br_0_417 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c417
+ bl_0_417 br_0_417 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c417
+ bl_0_417 br_0_417 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c417
+ bl_0_417 br_0_417 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c417
+ bl_0_417 br_0_417 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c418
+ bl_0_418 br_0_418 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c418
+ bl_0_418 br_0_418 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c418
+ bl_0_418 br_0_418 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c418
+ bl_0_418 br_0_418 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c418
+ bl_0_418 br_0_418 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c418
+ bl_0_418 br_0_418 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c418
+ bl_0_418 br_0_418 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c418
+ bl_0_418 br_0_418 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c418
+ bl_0_418 br_0_418 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c418
+ bl_0_418 br_0_418 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c418
+ bl_0_418 br_0_418 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c418
+ bl_0_418 br_0_418 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c418
+ bl_0_418 br_0_418 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c418
+ bl_0_418 br_0_418 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c418
+ bl_0_418 br_0_418 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c418
+ bl_0_418 br_0_418 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c418
+ bl_0_418 br_0_418 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c418
+ bl_0_418 br_0_418 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c418
+ bl_0_418 br_0_418 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c418
+ bl_0_418 br_0_418 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c418
+ bl_0_418 br_0_418 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c418
+ bl_0_418 br_0_418 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c418
+ bl_0_418 br_0_418 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c418
+ bl_0_418 br_0_418 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c418
+ bl_0_418 br_0_418 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c418
+ bl_0_418 br_0_418 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c418
+ bl_0_418 br_0_418 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c418
+ bl_0_418 br_0_418 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c418
+ bl_0_418 br_0_418 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c418
+ bl_0_418 br_0_418 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c418
+ bl_0_418 br_0_418 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c418
+ bl_0_418 br_0_418 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c418
+ bl_0_418 br_0_418 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c418
+ bl_0_418 br_0_418 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c418
+ bl_0_418 br_0_418 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c418
+ bl_0_418 br_0_418 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c418
+ bl_0_418 br_0_418 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c418
+ bl_0_418 br_0_418 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c418
+ bl_0_418 br_0_418 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c418
+ bl_0_418 br_0_418 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c418
+ bl_0_418 br_0_418 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c418
+ bl_0_418 br_0_418 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c418
+ bl_0_418 br_0_418 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c418
+ bl_0_418 br_0_418 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c418
+ bl_0_418 br_0_418 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c419
+ bl_0_419 br_0_419 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c419
+ bl_0_419 br_0_419 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c419
+ bl_0_419 br_0_419 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c419
+ bl_0_419 br_0_419 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c419
+ bl_0_419 br_0_419 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c419
+ bl_0_419 br_0_419 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c419
+ bl_0_419 br_0_419 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c419
+ bl_0_419 br_0_419 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c419
+ bl_0_419 br_0_419 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c419
+ bl_0_419 br_0_419 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c419
+ bl_0_419 br_0_419 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c419
+ bl_0_419 br_0_419 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c419
+ bl_0_419 br_0_419 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c419
+ bl_0_419 br_0_419 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c419
+ bl_0_419 br_0_419 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c419
+ bl_0_419 br_0_419 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c419
+ bl_0_419 br_0_419 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c419
+ bl_0_419 br_0_419 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c419
+ bl_0_419 br_0_419 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c419
+ bl_0_419 br_0_419 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c419
+ bl_0_419 br_0_419 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c419
+ bl_0_419 br_0_419 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c419
+ bl_0_419 br_0_419 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c419
+ bl_0_419 br_0_419 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c419
+ bl_0_419 br_0_419 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c419
+ bl_0_419 br_0_419 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c419
+ bl_0_419 br_0_419 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c419
+ bl_0_419 br_0_419 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c419
+ bl_0_419 br_0_419 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c419
+ bl_0_419 br_0_419 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c419
+ bl_0_419 br_0_419 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c419
+ bl_0_419 br_0_419 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c419
+ bl_0_419 br_0_419 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c419
+ bl_0_419 br_0_419 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c419
+ bl_0_419 br_0_419 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c419
+ bl_0_419 br_0_419 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c419
+ bl_0_419 br_0_419 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c419
+ bl_0_419 br_0_419 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c419
+ bl_0_419 br_0_419 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c419
+ bl_0_419 br_0_419 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c419
+ bl_0_419 br_0_419 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c419
+ bl_0_419 br_0_419 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c419
+ bl_0_419 br_0_419 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c419
+ bl_0_419 br_0_419 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c419
+ bl_0_419 br_0_419 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c420
+ bl_0_420 br_0_420 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c420
+ bl_0_420 br_0_420 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c420
+ bl_0_420 br_0_420 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c420
+ bl_0_420 br_0_420 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c420
+ bl_0_420 br_0_420 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c420
+ bl_0_420 br_0_420 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c420
+ bl_0_420 br_0_420 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c420
+ bl_0_420 br_0_420 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c420
+ bl_0_420 br_0_420 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c420
+ bl_0_420 br_0_420 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c420
+ bl_0_420 br_0_420 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c420
+ bl_0_420 br_0_420 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c420
+ bl_0_420 br_0_420 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c420
+ bl_0_420 br_0_420 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c420
+ bl_0_420 br_0_420 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c420
+ bl_0_420 br_0_420 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c420
+ bl_0_420 br_0_420 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c420
+ bl_0_420 br_0_420 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c420
+ bl_0_420 br_0_420 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c420
+ bl_0_420 br_0_420 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c420
+ bl_0_420 br_0_420 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c420
+ bl_0_420 br_0_420 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c420
+ bl_0_420 br_0_420 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c420
+ bl_0_420 br_0_420 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c420
+ bl_0_420 br_0_420 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c420
+ bl_0_420 br_0_420 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c420
+ bl_0_420 br_0_420 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c420
+ bl_0_420 br_0_420 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c420
+ bl_0_420 br_0_420 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c420
+ bl_0_420 br_0_420 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c420
+ bl_0_420 br_0_420 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c420
+ bl_0_420 br_0_420 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c420
+ bl_0_420 br_0_420 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c420
+ bl_0_420 br_0_420 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c420
+ bl_0_420 br_0_420 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c420
+ bl_0_420 br_0_420 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c420
+ bl_0_420 br_0_420 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c420
+ bl_0_420 br_0_420 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c420
+ bl_0_420 br_0_420 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c420
+ bl_0_420 br_0_420 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c420
+ bl_0_420 br_0_420 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c420
+ bl_0_420 br_0_420 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c420
+ bl_0_420 br_0_420 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c420
+ bl_0_420 br_0_420 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c420
+ bl_0_420 br_0_420 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c421
+ bl_0_421 br_0_421 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c421
+ bl_0_421 br_0_421 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c421
+ bl_0_421 br_0_421 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c421
+ bl_0_421 br_0_421 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c421
+ bl_0_421 br_0_421 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c421
+ bl_0_421 br_0_421 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c421
+ bl_0_421 br_0_421 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c421
+ bl_0_421 br_0_421 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c421
+ bl_0_421 br_0_421 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c421
+ bl_0_421 br_0_421 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c421
+ bl_0_421 br_0_421 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c421
+ bl_0_421 br_0_421 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c421
+ bl_0_421 br_0_421 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c421
+ bl_0_421 br_0_421 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c421
+ bl_0_421 br_0_421 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c421
+ bl_0_421 br_0_421 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c421
+ bl_0_421 br_0_421 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c421
+ bl_0_421 br_0_421 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c421
+ bl_0_421 br_0_421 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c421
+ bl_0_421 br_0_421 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c421
+ bl_0_421 br_0_421 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c421
+ bl_0_421 br_0_421 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c421
+ bl_0_421 br_0_421 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c421
+ bl_0_421 br_0_421 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c421
+ bl_0_421 br_0_421 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c421
+ bl_0_421 br_0_421 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c421
+ bl_0_421 br_0_421 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c421
+ bl_0_421 br_0_421 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c421
+ bl_0_421 br_0_421 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c421
+ bl_0_421 br_0_421 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c421
+ bl_0_421 br_0_421 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c421
+ bl_0_421 br_0_421 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c421
+ bl_0_421 br_0_421 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c421
+ bl_0_421 br_0_421 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c421
+ bl_0_421 br_0_421 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c421
+ bl_0_421 br_0_421 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c421
+ bl_0_421 br_0_421 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c421
+ bl_0_421 br_0_421 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c421
+ bl_0_421 br_0_421 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c421
+ bl_0_421 br_0_421 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c421
+ bl_0_421 br_0_421 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c421
+ bl_0_421 br_0_421 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c421
+ bl_0_421 br_0_421 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c421
+ bl_0_421 br_0_421 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c421
+ bl_0_421 br_0_421 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c422
+ bl_0_422 br_0_422 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c422
+ bl_0_422 br_0_422 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c422
+ bl_0_422 br_0_422 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c422
+ bl_0_422 br_0_422 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c422
+ bl_0_422 br_0_422 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c422
+ bl_0_422 br_0_422 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c422
+ bl_0_422 br_0_422 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c422
+ bl_0_422 br_0_422 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c422
+ bl_0_422 br_0_422 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c422
+ bl_0_422 br_0_422 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c422
+ bl_0_422 br_0_422 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c422
+ bl_0_422 br_0_422 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c422
+ bl_0_422 br_0_422 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c422
+ bl_0_422 br_0_422 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c422
+ bl_0_422 br_0_422 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c422
+ bl_0_422 br_0_422 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c422
+ bl_0_422 br_0_422 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c422
+ bl_0_422 br_0_422 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c422
+ bl_0_422 br_0_422 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c422
+ bl_0_422 br_0_422 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c422
+ bl_0_422 br_0_422 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c422
+ bl_0_422 br_0_422 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c422
+ bl_0_422 br_0_422 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c422
+ bl_0_422 br_0_422 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c422
+ bl_0_422 br_0_422 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c422
+ bl_0_422 br_0_422 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c422
+ bl_0_422 br_0_422 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c422
+ bl_0_422 br_0_422 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c422
+ bl_0_422 br_0_422 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c422
+ bl_0_422 br_0_422 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c422
+ bl_0_422 br_0_422 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c422
+ bl_0_422 br_0_422 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c422
+ bl_0_422 br_0_422 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c422
+ bl_0_422 br_0_422 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c422
+ bl_0_422 br_0_422 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c422
+ bl_0_422 br_0_422 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c422
+ bl_0_422 br_0_422 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c422
+ bl_0_422 br_0_422 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c422
+ bl_0_422 br_0_422 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c422
+ bl_0_422 br_0_422 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c422
+ bl_0_422 br_0_422 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c422
+ bl_0_422 br_0_422 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c422
+ bl_0_422 br_0_422 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c422
+ bl_0_422 br_0_422 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c422
+ bl_0_422 br_0_422 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c423
+ bl_0_423 br_0_423 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c423
+ bl_0_423 br_0_423 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c423
+ bl_0_423 br_0_423 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c423
+ bl_0_423 br_0_423 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c423
+ bl_0_423 br_0_423 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c423
+ bl_0_423 br_0_423 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c423
+ bl_0_423 br_0_423 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c423
+ bl_0_423 br_0_423 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c423
+ bl_0_423 br_0_423 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c423
+ bl_0_423 br_0_423 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c423
+ bl_0_423 br_0_423 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c423
+ bl_0_423 br_0_423 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c423
+ bl_0_423 br_0_423 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c423
+ bl_0_423 br_0_423 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c423
+ bl_0_423 br_0_423 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c423
+ bl_0_423 br_0_423 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c423
+ bl_0_423 br_0_423 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c423
+ bl_0_423 br_0_423 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c423
+ bl_0_423 br_0_423 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c423
+ bl_0_423 br_0_423 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c423
+ bl_0_423 br_0_423 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c423
+ bl_0_423 br_0_423 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c423
+ bl_0_423 br_0_423 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c423
+ bl_0_423 br_0_423 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c423
+ bl_0_423 br_0_423 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c423
+ bl_0_423 br_0_423 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c423
+ bl_0_423 br_0_423 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c423
+ bl_0_423 br_0_423 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c423
+ bl_0_423 br_0_423 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c423
+ bl_0_423 br_0_423 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c423
+ bl_0_423 br_0_423 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c423
+ bl_0_423 br_0_423 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c423
+ bl_0_423 br_0_423 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c423
+ bl_0_423 br_0_423 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c423
+ bl_0_423 br_0_423 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c423
+ bl_0_423 br_0_423 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c423
+ bl_0_423 br_0_423 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c423
+ bl_0_423 br_0_423 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c423
+ bl_0_423 br_0_423 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c423
+ bl_0_423 br_0_423 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c423
+ bl_0_423 br_0_423 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c423
+ bl_0_423 br_0_423 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c423
+ bl_0_423 br_0_423 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c423
+ bl_0_423 br_0_423 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c423
+ bl_0_423 br_0_423 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c424
+ bl_0_424 br_0_424 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c424
+ bl_0_424 br_0_424 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c424
+ bl_0_424 br_0_424 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c424
+ bl_0_424 br_0_424 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c424
+ bl_0_424 br_0_424 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c424
+ bl_0_424 br_0_424 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c424
+ bl_0_424 br_0_424 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c424
+ bl_0_424 br_0_424 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c424
+ bl_0_424 br_0_424 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c424
+ bl_0_424 br_0_424 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c424
+ bl_0_424 br_0_424 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c424
+ bl_0_424 br_0_424 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c424
+ bl_0_424 br_0_424 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c424
+ bl_0_424 br_0_424 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c424
+ bl_0_424 br_0_424 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c424
+ bl_0_424 br_0_424 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c424
+ bl_0_424 br_0_424 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c424
+ bl_0_424 br_0_424 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c424
+ bl_0_424 br_0_424 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c424
+ bl_0_424 br_0_424 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c424
+ bl_0_424 br_0_424 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c424
+ bl_0_424 br_0_424 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c424
+ bl_0_424 br_0_424 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c424
+ bl_0_424 br_0_424 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c424
+ bl_0_424 br_0_424 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c424
+ bl_0_424 br_0_424 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c424
+ bl_0_424 br_0_424 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c424
+ bl_0_424 br_0_424 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c424
+ bl_0_424 br_0_424 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c424
+ bl_0_424 br_0_424 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c424
+ bl_0_424 br_0_424 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c424
+ bl_0_424 br_0_424 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c424
+ bl_0_424 br_0_424 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c424
+ bl_0_424 br_0_424 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c424
+ bl_0_424 br_0_424 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c424
+ bl_0_424 br_0_424 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c424
+ bl_0_424 br_0_424 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c424
+ bl_0_424 br_0_424 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c424
+ bl_0_424 br_0_424 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c424
+ bl_0_424 br_0_424 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c424
+ bl_0_424 br_0_424 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c424
+ bl_0_424 br_0_424 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c424
+ bl_0_424 br_0_424 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c424
+ bl_0_424 br_0_424 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c424
+ bl_0_424 br_0_424 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c425
+ bl_0_425 br_0_425 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c425
+ bl_0_425 br_0_425 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c425
+ bl_0_425 br_0_425 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c425
+ bl_0_425 br_0_425 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c425
+ bl_0_425 br_0_425 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c425
+ bl_0_425 br_0_425 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c425
+ bl_0_425 br_0_425 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c425
+ bl_0_425 br_0_425 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c425
+ bl_0_425 br_0_425 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c425
+ bl_0_425 br_0_425 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c425
+ bl_0_425 br_0_425 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c425
+ bl_0_425 br_0_425 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c425
+ bl_0_425 br_0_425 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c425
+ bl_0_425 br_0_425 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c425
+ bl_0_425 br_0_425 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c425
+ bl_0_425 br_0_425 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c425
+ bl_0_425 br_0_425 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c425
+ bl_0_425 br_0_425 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c425
+ bl_0_425 br_0_425 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c425
+ bl_0_425 br_0_425 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c425
+ bl_0_425 br_0_425 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c425
+ bl_0_425 br_0_425 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c425
+ bl_0_425 br_0_425 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c425
+ bl_0_425 br_0_425 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c425
+ bl_0_425 br_0_425 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c425
+ bl_0_425 br_0_425 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c425
+ bl_0_425 br_0_425 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c425
+ bl_0_425 br_0_425 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c425
+ bl_0_425 br_0_425 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c425
+ bl_0_425 br_0_425 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c425
+ bl_0_425 br_0_425 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c425
+ bl_0_425 br_0_425 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c425
+ bl_0_425 br_0_425 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c425
+ bl_0_425 br_0_425 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c425
+ bl_0_425 br_0_425 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c425
+ bl_0_425 br_0_425 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c425
+ bl_0_425 br_0_425 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c425
+ bl_0_425 br_0_425 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c425
+ bl_0_425 br_0_425 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c425
+ bl_0_425 br_0_425 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c425
+ bl_0_425 br_0_425 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c425
+ bl_0_425 br_0_425 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c425
+ bl_0_425 br_0_425 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c425
+ bl_0_425 br_0_425 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c425
+ bl_0_425 br_0_425 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c426
+ bl_0_426 br_0_426 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c426
+ bl_0_426 br_0_426 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c426
+ bl_0_426 br_0_426 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c426
+ bl_0_426 br_0_426 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c426
+ bl_0_426 br_0_426 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c426
+ bl_0_426 br_0_426 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c426
+ bl_0_426 br_0_426 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c426
+ bl_0_426 br_0_426 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c426
+ bl_0_426 br_0_426 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c426
+ bl_0_426 br_0_426 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c426
+ bl_0_426 br_0_426 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c426
+ bl_0_426 br_0_426 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c426
+ bl_0_426 br_0_426 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c426
+ bl_0_426 br_0_426 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c426
+ bl_0_426 br_0_426 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c426
+ bl_0_426 br_0_426 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c426
+ bl_0_426 br_0_426 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c426
+ bl_0_426 br_0_426 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c426
+ bl_0_426 br_0_426 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c426
+ bl_0_426 br_0_426 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c426
+ bl_0_426 br_0_426 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c426
+ bl_0_426 br_0_426 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c426
+ bl_0_426 br_0_426 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c426
+ bl_0_426 br_0_426 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c426
+ bl_0_426 br_0_426 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c426
+ bl_0_426 br_0_426 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c426
+ bl_0_426 br_0_426 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c426
+ bl_0_426 br_0_426 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c426
+ bl_0_426 br_0_426 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c426
+ bl_0_426 br_0_426 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c426
+ bl_0_426 br_0_426 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c426
+ bl_0_426 br_0_426 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c426
+ bl_0_426 br_0_426 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c426
+ bl_0_426 br_0_426 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c426
+ bl_0_426 br_0_426 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c426
+ bl_0_426 br_0_426 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c426
+ bl_0_426 br_0_426 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c426
+ bl_0_426 br_0_426 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c426
+ bl_0_426 br_0_426 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c426
+ bl_0_426 br_0_426 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c426
+ bl_0_426 br_0_426 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c426
+ bl_0_426 br_0_426 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c426
+ bl_0_426 br_0_426 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c426
+ bl_0_426 br_0_426 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c426
+ bl_0_426 br_0_426 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c427
+ bl_0_427 br_0_427 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c427
+ bl_0_427 br_0_427 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c427
+ bl_0_427 br_0_427 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c427
+ bl_0_427 br_0_427 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c427
+ bl_0_427 br_0_427 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c427
+ bl_0_427 br_0_427 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c427
+ bl_0_427 br_0_427 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c427
+ bl_0_427 br_0_427 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c427
+ bl_0_427 br_0_427 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c427
+ bl_0_427 br_0_427 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c427
+ bl_0_427 br_0_427 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c427
+ bl_0_427 br_0_427 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c427
+ bl_0_427 br_0_427 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c427
+ bl_0_427 br_0_427 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c427
+ bl_0_427 br_0_427 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c427
+ bl_0_427 br_0_427 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c427
+ bl_0_427 br_0_427 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c427
+ bl_0_427 br_0_427 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c427
+ bl_0_427 br_0_427 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c427
+ bl_0_427 br_0_427 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c427
+ bl_0_427 br_0_427 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c427
+ bl_0_427 br_0_427 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c427
+ bl_0_427 br_0_427 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c427
+ bl_0_427 br_0_427 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c427
+ bl_0_427 br_0_427 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c427
+ bl_0_427 br_0_427 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c427
+ bl_0_427 br_0_427 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c427
+ bl_0_427 br_0_427 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c427
+ bl_0_427 br_0_427 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c427
+ bl_0_427 br_0_427 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c427
+ bl_0_427 br_0_427 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c427
+ bl_0_427 br_0_427 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c427
+ bl_0_427 br_0_427 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c427
+ bl_0_427 br_0_427 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c427
+ bl_0_427 br_0_427 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c427
+ bl_0_427 br_0_427 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c427
+ bl_0_427 br_0_427 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c427
+ bl_0_427 br_0_427 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c427
+ bl_0_427 br_0_427 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c427
+ bl_0_427 br_0_427 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c427
+ bl_0_427 br_0_427 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c427
+ bl_0_427 br_0_427 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c427
+ bl_0_427 br_0_427 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c427
+ bl_0_427 br_0_427 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c427
+ bl_0_427 br_0_427 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c428
+ bl_0_428 br_0_428 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c428
+ bl_0_428 br_0_428 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c428
+ bl_0_428 br_0_428 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c428
+ bl_0_428 br_0_428 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c428
+ bl_0_428 br_0_428 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c428
+ bl_0_428 br_0_428 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c428
+ bl_0_428 br_0_428 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c428
+ bl_0_428 br_0_428 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c428
+ bl_0_428 br_0_428 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c428
+ bl_0_428 br_0_428 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c428
+ bl_0_428 br_0_428 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c428
+ bl_0_428 br_0_428 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c428
+ bl_0_428 br_0_428 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c428
+ bl_0_428 br_0_428 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c428
+ bl_0_428 br_0_428 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c428
+ bl_0_428 br_0_428 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c428
+ bl_0_428 br_0_428 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c428
+ bl_0_428 br_0_428 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c428
+ bl_0_428 br_0_428 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c428
+ bl_0_428 br_0_428 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c428
+ bl_0_428 br_0_428 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c428
+ bl_0_428 br_0_428 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c428
+ bl_0_428 br_0_428 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c428
+ bl_0_428 br_0_428 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c428
+ bl_0_428 br_0_428 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c428
+ bl_0_428 br_0_428 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c428
+ bl_0_428 br_0_428 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c428
+ bl_0_428 br_0_428 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c428
+ bl_0_428 br_0_428 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c428
+ bl_0_428 br_0_428 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c428
+ bl_0_428 br_0_428 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c428
+ bl_0_428 br_0_428 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c428
+ bl_0_428 br_0_428 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c428
+ bl_0_428 br_0_428 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c428
+ bl_0_428 br_0_428 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c428
+ bl_0_428 br_0_428 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c428
+ bl_0_428 br_0_428 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c428
+ bl_0_428 br_0_428 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c428
+ bl_0_428 br_0_428 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c428
+ bl_0_428 br_0_428 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c428
+ bl_0_428 br_0_428 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c428
+ bl_0_428 br_0_428 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c428
+ bl_0_428 br_0_428 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c428
+ bl_0_428 br_0_428 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c428
+ bl_0_428 br_0_428 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c429
+ bl_0_429 br_0_429 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c429
+ bl_0_429 br_0_429 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c429
+ bl_0_429 br_0_429 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c429
+ bl_0_429 br_0_429 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c429
+ bl_0_429 br_0_429 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c429
+ bl_0_429 br_0_429 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c429
+ bl_0_429 br_0_429 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c429
+ bl_0_429 br_0_429 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c429
+ bl_0_429 br_0_429 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c429
+ bl_0_429 br_0_429 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c429
+ bl_0_429 br_0_429 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c429
+ bl_0_429 br_0_429 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c429
+ bl_0_429 br_0_429 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c429
+ bl_0_429 br_0_429 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c429
+ bl_0_429 br_0_429 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c429
+ bl_0_429 br_0_429 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c429
+ bl_0_429 br_0_429 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c429
+ bl_0_429 br_0_429 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c429
+ bl_0_429 br_0_429 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c429
+ bl_0_429 br_0_429 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c429
+ bl_0_429 br_0_429 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c429
+ bl_0_429 br_0_429 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c429
+ bl_0_429 br_0_429 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c429
+ bl_0_429 br_0_429 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c429
+ bl_0_429 br_0_429 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c429
+ bl_0_429 br_0_429 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c429
+ bl_0_429 br_0_429 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c429
+ bl_0_429 br_0_429 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c429
+ bl_0_429 br_0_429 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c429
+ bl_0_429 br_0_429 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c429
+ bl_0_429 br_0_429 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c429
+ bl_0_429 br_0_429 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c429
+ bl_0_429 br_0_429 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c429
+ bl_0_429 br_0_429 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c429
+ bl_0_429 br_0_429 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c429
+ bl_0_429 br_0_429 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c429
+ bl_0_429 br_0_429 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c429
+ bl_0_429 br_0_429 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c429
+ bl_0_429 br_0_429 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c429
+ bl_0_429 br_0_429 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c429
+ bl_0_429 br_0_429 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c429
+ bl_0_429 br_0_429 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c429
+ bl_0_429 br_0_429 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c429
+ bl_0_429 br_0_429 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c429
+ bl_0_429 br_0_429 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c430
+ bl_0_430 br_0_430 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c430
+ bl_0_430 br_0_430 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c430
+ bl_0_430 br_0_430 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c430
+ bl_0_430 br_0_430 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c430
+ bl_0_430 br_0_430 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c430
+ bl_0_430 br_0_430 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c430
+ bl_0_430 br_0_430 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c430
+ bl_0_430 br_0_430 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c430
+ bl_0_430 br_0_430 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c430
+ bl_0_430 br_0_430 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c430
+ bl_0_430 br_0_430 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c430
+ bl_0_430 br_0_430 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c430
+ bl_0_430 br_0_430 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c430
+ bl_0_430 br_0_430 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c430
+ bl_0_430 br_0_430 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c430
+ bl_0_430 br_0_430 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c430
+ bl_0_430 br_0_430 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c430
+ bl_0_430 br_0_430 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c430
+ bl_0_430 br_0_430 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c430
+ bl_0_430 br_0_430 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c430
+ bl_0_430 br_0_430 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c430
+ bl_0_430 br_0_430 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c430
+ bl_0_430 br_0_430 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c430
+ bl_0_430 br_0_430 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c430
+ bl_0_430 br_0_430 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c430
+ bl_0_430 br_0_430 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c430
+ bl_0_430 br_0_430 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c430
+ bl_0_430 br_0_430 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c430
+ bl_0_430 br_0_430 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c430
+ bl_0_430 br_0_430 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c430
+ bl_0_430 br_0_430 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c430
+ bl_0_430 br_0_430 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c430
+ bl_0_430 br_0_430 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c430
+ bl_0_430 br_0_430 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c430
+ bl_0_430 br_0_430 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c430
+ bl_0_430 br_0_430 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c430
+ bl_0_430 br_0_430 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c430
+ bl_0_430 br_0_430 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c430
+ bl_0_430 br_0_430 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c430
+ bl_0_430 br_0_430 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c430
+ bl_0_430 br_0_430 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c430
+ bl_0_430 br_0_430 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c430
+ bl_0_430 br_0_430 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c430
+ bl_0_430 br_0_430 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c430
+ bl_0_430 br_0_430 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c431
+ bl_0_431 br_0_431 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c431
+ bl_0_431 br_0_431 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c431
+ bl_0_431 br_0_431 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c431
+ bl_0_431 br_0_431 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c431
+ bl_0_431 br_0_431 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c431
+ bl_0_431 br_0_431 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c431
+ bl_0_431 br_0_431 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c431
+ bl_0_431 br_0_431 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c431
+ bl_0_431 br_0_431 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c431
+ bl_0_431 br_0_431 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c431
+ bl_0_431 br_0_431 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c431
+ bl_0_431 br_0_431 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c431
+ bl_0_431 br_0_431 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c431
+ bl_0_431 br_0_431 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c431
+ bl_0_431 br_0_431 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c431
+ bl_0_431 br_0_431 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c431
+ bl_0_431 br_0_431 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c431
+ bl_0_431 br_0_431 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c431
+ bl_0_431 br_0_431 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c431
+ bl_0_431 br_0_431 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c431
+ bl_0_431 br_0_431 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c431
+ bl_0_431 br_0_431 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c431
+ bl_0_431 br_0_431 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c431
+ bl_0_431 br_0_431 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c431
+ bl_0_431 br_0_431 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c431
+ bl_0_431 br_0_431 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c431
+ bl_0_431 br_0_431 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c431
+ bl_0_431 br_0_431 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c431
+ bl_0_431 br_0_431 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c431
+ bl_0_431 br_0_431 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c431
+ bl_0_431 br_0_431 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c431
+ bl_0_431 br_0_431 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c431
+ bl_0_431 br_0_431 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c431
+ bl_0_431 br_0_431 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c431
+ bl_0_431 br_0_431 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c431
+ bl_0_431 br_0_431 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c431
+ bl_0_431 br_0_431 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c431
+ bl_0_431 br_0_431 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c431
+ bl_0_431 br_0_431 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c431
+ bl_0_431 br_0_431 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c431
+ bl_0_431 br_0_431 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c431
+ bl_0_431 br_0_431 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c431
+ bl_0_431 br_0_431 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c431
+ bl_0_431 br_0_431 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c431
+ bl_0_431 br_0_431 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c432
+ bl_0_432 br_0_432 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c432
+ bl_0_432 br_0_432 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c432
+ bl_0_432 br_0_432 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c432
+ bl_0_432 br_0_432 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c432
+ bl_0_432 br_0_432 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c432
+ bl_0_432 br_0_432 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c432
+ bl_0_432 br_0_432 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c432
+ bl_0_432 br_0_432 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c432
+ bl_0_432 br_0_432 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c432
+ bl_0_432 br_0_432 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c432
+ bl_0_432 br_0_432 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c432
+ bl_0_432 br_0_432 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c432
+ bl_0_432 br_0_432 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c432
+ bl_0_432 br_0_432 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c432
+ bl_0_432 br_0_432 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c432
+ bl_0_432 br_0_432 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c432
+ bl_0_432 br_0_432 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c432
+ bl_0_432 br_0_432 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c432
+ bl_0_432 br_0_432 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c432
+ bl_0_432 br_0_432 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c432
+ bl_0_432 br_0_432 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c432
+ bl_0_432 br_0_432 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c432
+ bl_0_432 br_0_432 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c432
+ bl_0_432 br_0_432 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c432
+ bl_0_432 br_0_432 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c432
+ bl_0_432 br_0_432 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c432
+ bl_0_432 br_0_432 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c432
+ bl_0_432 br_0_432 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c432
+ bl_0_432 br_0_432 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c432
+ bl_0_432 br_0_432 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c432
+ bl_0_432 br_0_432 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c432
+ bl_0_432 br_0_432 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c432
+ bl_0_432 br_0_432 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c432
+ bl_0_432 br_0_432 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c432
+ bl_0_432 br_0_432 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c432
+ bl_0_432 br_0_432 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c432
+ bl_0_432 br_0_432 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c432
+ bl_0_432 br_0_432 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c432
+ bl_0_432 br_0_432 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c432
+ bl_0_432 br_0_432 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c432
+ bl_0_432 br_0_432 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c432
+ bl_0_432 br_0_432 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c432
+ bl_0_432 br_0_432 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c432
+ bl_0_432 br_0_432 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c432
+ bl_0_432 br_0_432 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c433
+ bl_0_433 br_0_433 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c433
+ bl_0_433 br_0_433 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c433
+ bl_0_433 br_0_433 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c433
+ bl_0_433 br_0_433 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c433
+ bl_0_433 br_0_433 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c433
+ bl_0_433 br_0_433 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c433
+ bl_0_433 br_0_433 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c433
+ bl_0_433 br_0_433 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c433
+ bl_0_433 br_0_433 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c433
+ bl_0_433 br_0_433 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c433
+ bl_0_433 br_0_433 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c433
+ bl_0_433 br_0_433 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c433
+ bl_0_433 br_0_433 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c433
+ bl_0_433 br_0_433 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c433
+ bl_0_433 br_0_433 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c433
+ bl_0_433 br_0_433 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c433
+ bl_0_433 br_0_433 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c433
+ bl_0_433 br_0_433 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c433
+ bl_0_433 br_0_433 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c433
+ bl_0_433 br_0_433 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c433
+ bl_0_433 br_0_433 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c433
+ bl_0_433 br_0_433 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c433
+ bl_0_433 br_0_433 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c433
+ bl_0_433 br_0_433 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c433
+ bl_0_433 br_0_433 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c433
+ bl_0_433 br_0_433 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c433
+ bl_0_433 br_0_433 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c433
+ bl_0_433 br_0_433 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c433
+ bl_0_433 br_0_433 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c433
+ bl_0_433 br_0_433 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c433
+ bl_0_433 br_0_433 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c433
+ bl_0_433 br_0_433 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c433
+ bl_0_433 br_0_433 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c433
+ bl_0_433 br_0_433 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c433
+ bl_0_433 br_0_433 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c433
+ bl_0_433 br_0_433 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c433
+ bl_0_433 br_0_433 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c433
+ bl_0_433 br_0_433 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c433
+ bl_0_433 br_0_433 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c433
+ bl_0_433 br_0_433 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c433
+ bl_0_433 br_0_433 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c433
+ bl_0_433 br_0_433 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c433
+ bl_0_433 br_0_433 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c433
+ bl_0_433 br_0_433 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c433
+ bl_0_433 br_0_433 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c434
+ bl_0_434 br_0_434 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c434
+ bl_0_434 br_0_434 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c434
+ bl_0_434 br_0_434 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c434
+ bl_0_434 br_0_434 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c434
+ bl_0_434 br_0_434 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c434
+ bl_0_434 br_0_434 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c434
+ bl_0_434 br_0_434 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c434
+ bl_0_434 br_0_434 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c434
+ bl_0_434 br_0_434 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c434
+ bl_0_434 br_0_434 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c434
+ bl_0_434 br_0_434 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c434
+ bl_0_434 br_0_434 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c434
+ bl_0_434 br_0_434 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c434
+ bl_0_434 br_0_434 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c434
+ bl_0_434 br_0_434 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c434
+ bl_0_434 br_0_434 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c434
+ bl_0_434 br_0_434 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c434
+ bl_0_434 br_0_434 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c434
+ bl_0_434 br_0_434 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c434
+ bl_0_434 br_0_434 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c434
+ bl_0_434 br_0_434 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c434
+ bl_0_434 br_0_434 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c434
+ bl_0_434 br_0_434 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c434
+ bl_0_434 br_0_434 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c434
+ bl_0_434 br_0_434 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c434
+ bl_0_434 br_0_434 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c434
+ bl_0_434 br_0_434 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c434
+ bl_0_434 br_0_434 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c434
+ bl_0_434 br_0_434 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c434
+ bl_0_434 br_0_434 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c434
+ bl_0_434 br_0_434 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c434
+ bl_0_434 br_0_434 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c434
+ bl_0_434 br_0_434 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c434
+ bl_0_434 br_0_434 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c434
+ bl_0_434 br_0_434 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c434
+ bl_0_434 br_0_434 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c434
+ bl_0_434 br_0_434 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c434
+ bl_0_434 br_0_434 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c434
+ bl_0_434 br_0_434 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c434
+ bl_0_434 br_0_434 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c434
+ bl_0_434 br_0_434 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c434
+ bl_0_434 br_0_434 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c434
+ bl_0_434 br_0_434 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c434
+ bl_0_434 br_0_434 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c434
+ bl_0_434 br_0_434 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c435
+ bl_0_435 br_0_435 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c435
+ bl_0_435 br_0_435 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c435
+ bl_0_435 br_0_435 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c435
+ bl_0_435 br_0_435 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c435
+ bl_0_435 br_0_435 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c435
+ bl_0_435 br_0_435 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c435
+ bl_0_435 br_0_435 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c435
+ bl_0_435 br_0_435 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c435
+ bl_0_435 br_0_435 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c435
+ bl_0_435 br_0_435 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c435
+ bl_0_435 br_0_435 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c435
+ bl_0_435 br_0_435 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c435
+ bl_0_435 br_0_435 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c435
+ bl_0_435 br_0_435 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c435
+ bl_0_435 br_0_435 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c435
+ bl_0_435 br_0_435 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c435
+ bl_0_435 br_0_435 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c435
+ bl_0_435 br_0_435 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c435
+ bl_0_435 br_0_435 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c435
+ bl_0_435 br_0_435 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c435
+ bl_0_435 br_0_435 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c435
+ bl_0_435 br_0_435 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c435
+ bl_0_435 br_0_435 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c435
+ bl_0_435 br_0_435 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c435
+ bl_0_435 br_0_435 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c435
+ bl_0_435 br_0_435 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c435
+ bl_0_435 br_0_435 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c435
+ bl_0_435 br_0_435 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c435
+ bl_0_435 br_0_435 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c435
+ bl_0_435 br_0_435 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c435
+ bl_0_435 br_0_435 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c435
+ bl_0_435 br_0_435 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c435
+ bl_0_435 br_0_435 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c435
+ bl_0_435 br_0_435 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c435
+ bl_0_435 br_0_435 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c435
+ bl_0_435 br_0_435 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c435
+ bl_0_435 br_0_435 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c435
+ bl_0_435 br_0_435 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c435
+ bl_0_435 br_0_435 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c435
+ bl_0_435 br_0_435 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c435
+ bl_0_435 br_0_435 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c435
+ bl_0_435 br_0_435 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c435
+ bl_0_435 br_0_435 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c435
+ bl_0_435 br_0_435 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c435
+ bl_0_435 br_0_435 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c436
+ bl_0_436 br_0_436 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c436
+ bl_0_436 br_0_436 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c436
+ bl_0_436 br_0_436 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c436
+ bl_0_436 br_0_436 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c436
+ bl_0_436 br_0_436 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c436
+ bl_0_436 br_0_436 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c436
+ bl_0_436 br_0_436 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c436
+ bl_0_436 br_0_436 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c436
+ bl_0_436 br_0_436 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c436
+ bl_0_436 br_0_436 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c436
+ bl_0_436 br_0_436 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c436
+ bl_0_436 br_0_436 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c436
+ bl_0_436 br_0_436 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c436
+ bl_0_436 br_0_436 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c436
+ bl_0_436 br_0_436 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c436
+ bl_0_436 br_0_436 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c436
+ bl_0_436 br_0_436 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c436
+ bl_0_436 br_0_436 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c436
+ bl_0_436 br_0_436 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c436
+ bl_0_436 br_0_436 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c436
+ bl_0_436 br_0_436 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c436
+ bl_0_436 br_0_436 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c436
+ bl_0_436 br_0_436 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c436
+ bl_0_436 br_0_436 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c436
+ bl_0_436 br_0_436 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c436
+ bl_0_436 br_0_436 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c436
+ bl_0_436 br_0_436 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c436
+ bl_0_436 br_0_436 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c436
+ bl_0_436 br_0_436 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c436
+ bl_0_436 br_0_436 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c436
+ bl_0_436 br_0_436 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c436
+ bl_0_436 br_0_436 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c436
+ bl_0_436 br_0_436 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c436
+ bl_0_436 br_0_436 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c436
+ bl_0_436 br_0_436 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c436
+ bl_0_436 br_0_436 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c436
+ bl_0_436 br_0_436 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c436
+ bl_0_436 br_0_436 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c436
+ bl_0_436 br_0_436 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c436
+ bl_0_436 br_0_436 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c436
+ bl_0_436 br_0_436 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c436
+ bl_0_436 br_0_436 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c436
+ bl_0_436 br_0_436 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c436
+ bl_0_436 br_0_436 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c436
+ bl_0_436 br_0_436 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c437
+ bl_0_437 br_0_437 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c437
+ bl_0_437 br_0_437 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c437
+ bl_0_437 br_0_437 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c437
+ bl_0_437 br_0_437 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c437
+ bl_0_437 br_0_437 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c437
+ bl_0_437 br_0_437 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c437
+ bl_0_437 br_0_437 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c437
+ bl_0_437 br_0_437 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c437
+ bl_0_437 br_0_437 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c437
+ bl_0_437 br_0_437 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c437
+ bl_0_437 br_0_437 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c437
+ bl_0_437 br_0_437 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c437
+ bl_0_437 br_0_437 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c437
+ bl_0_437 br_0_437 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c437
+ bl_0_437 br_0_437 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c437
+ bl_0_437 br_0_437 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c437
+ bl_0_437 br_0_437 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c437
+ bl_0_437 br_0_437 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c437
+ bl_0_437 br_0_437 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c437
+ bl_0_437 br_0_437 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c437
+ bl_0_437 br_0_437 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c437
+ bl_0_437 br_0_437 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c437
+ bl_0_437 br_0_437 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c437
+ bl_0_437 br_0_437 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c437
+ bl_0_437 br_0_437 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c437
+ bl_0_437 br_0_437 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c437
+ bl_0_437 br_0_437 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c437
+ bl_0_437 br_0_437 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c437
+ bl_0_437 br_0_437 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c437
+ bl_0_437 br_0_437 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c437
+ bl_0_437 br_0_437 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c437
+ bl_0_437 br_0_437 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c437
+ bl_0_437 br_0_437 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c437
+ bl_0_437 br_0_437 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c437
+ bl_0_437 br_0_437 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c437
+ bl_0_437 br_0_437 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c437
+ bl_0_437 br_0_437 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c437
+ bl_0_437 br_0_437 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c437
+ bl_0_437 br_0_437 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c437
+ bl_0_437 br_0_437 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c437
+ bl_0_437 br_0_437 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c437
+ bl_0_437 br_0_437 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c437
+ bl_0_437 br_0_437 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c437
+ bl_0_437 br_0_437 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c437
+ bl_0_437 br_0_437 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c438
+ bl_0_438 br_0_438 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c438
+ bl_0_438 br_0_438 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c438
+ bl_0_438 br_0_438 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c438
+ bl_0_438 br_0_438 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c438
+ bl_0_438 br_0_438 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c438
+ bl_0_438 br_0_438 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c438
+ bl_0_438 br_0_438 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c438
+ bl_0_438 br_0_438 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c438
+ bl_0_438 br_0_438 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c438
+ bl_0_438 br_0_438 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c438
+ bl_0_438 br_0_438 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c438
+ bl_0_438 br_0_438 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c438
+ bl_0_438 br_0_438 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c438
+ bl_0_438 br_0_438 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c438
+ bl_0_438 br_0_438 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c438
+ bl_0_438 br_0_438 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c438
+ bl_0_438 br_0_438 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c438
+ bl_0_438 br_0_438 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c438
+ bl_0_438 br_0_438 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c438
+ bl_0_438 br_0_438 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c438
+ bl_0_438 br_0_438 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c438
+ bl_0_438 br_0_438 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c438
+ bl_0_438 br_0_438 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c438
+ bl_0_438 br_0_438 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c438
+ bl_0_438 br_0_438 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c438
+ bl_0_438 br_0_438 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c438
+ bl_0_438 br_0_438 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c438
+ bl_0_438 br_0_438 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c438
+ bl_0_438 br_0_438 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c438
+ bl_0_438 br_0_438 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c438
+ bl_0_438 br_0_438 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c438
+ bl_0_438 br_0_438 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c438
+ bl_0_438 br_0_438 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c438
+ bl_0_438 br_0_438 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c438
+ bl_0_438 br_0_438 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c438
+ bl_0_438 br_0_438 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c438
+ bl_0_438 br_0_438 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c438
+ bl_0_438 br_0_438 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c438
+ bl_0_438 br_0_438 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c438
+ bl_0_438 br_0_438 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c438
+ bl_0_438 br_0_438 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c438
+ bl_0_438 br_0_438 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c438
+ bl_0_438 br_0_438 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c438
+ bl_0_438 br_0_438 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c438
+ bl_0_438 br_0_438 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c439
+ bl_0_439 br_0_439 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c439
+ bl_0_439 br_0_439 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c439
+ bl_0_439 br_0_439 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c439
+ bl_0_439 br_0_439 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c439
+ bl_0_439 br_0_439 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c439
+ bl_0_439 br_0_439 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c439
+ bl_0_439 br_0_439 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c439
+ bl_0_439 br_0_439 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c439
+ bl_0_439 br_0_439 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c439
+ bl_0_439 br_0_439 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c439
+ bl_0_439 br_0_439 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c439
+ bl_0_439 br_0_439 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c439
+ bl_0_439 br_0_439 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c439
+ bl_0_439 br_0_439 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c439
+ bl_0_439 br_0_439 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c439
+ bl_0_439 br_0_439 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c439
+ bl_0_439 br_0_439 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c439
+ bl_0_439 br_0_439 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c439
+ bl_0_439 br_0_439 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c439
+ bl_0_439 br_0_439 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c439
+ bl_0_439 br_0_439 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c439
+ bl_0_439 br_0_439 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c439
+ bl_0_439 br_0_439 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c439
+ bl_0_439 br_0_439 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c439
+ bl_0_439 br_0_439 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c439
+ bl_0_439 br_0_439 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c439
+ bl_0_439 br_0_439 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c439
+ bl_0_439 br_0_439 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c439
+ bl_0_439 br_0_439 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c439
+ bl_0_439 br_0_439 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c439
+ bl_0_439 br_0_439 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c439
+ bl_0_439 br_0_439 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c439
+ bl_0_439 br_0_439 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c439
+ bl_0_439 br_0_439 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c439
+ bl_0_439 br_0_439 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c439
+ bl_0_439 br_0_439 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c439
+ bl_0_439 br_0_439 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c439
+ bl_0_439 br_0_439 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c439
+ bl_0_439 br_0_439 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c439
+ bl_0_439 br_0_439 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c439
+ bl_0_439 br_0_439 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c439
+ bl_0_439 br_0_439 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c439
+ bl_0_439 br_0_439 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c439
+ bl_0_439 br_0_439 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c439
+ bl_0_439 br_0_439 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c440
+ bl_0_440 br_0_440 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c440
+ bl_0_440 br_0_440 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c440
+ bl_0_440 br_0_440 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c440
+ bl_0_440 br_0_440 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c440
+ bl_0_440 br_0_440 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c440
+ bl_0_440 br_0_440 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c440
+ bl_0_440 br_0_440 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c440
+ bl_0_440 br_0_440 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c440
+ bl_0_440 br_0_440 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c440
+ bl_0_440 br_0_440 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c440
+ bl_0_440 br_0_440 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c440
+ bl_0_440 br_0_440 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c440
+ bl_0_440 br_0_440 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c440
+ bl_0_440 br_0_440 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c440
+ bl_0_440 br_0_440 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c440
+ bl_0_440 br_0_440 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c440
+ bl_0_440 br_0_440 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c440
+ bl_0_440 br_0_440 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c440
+ bl_0_440 br_0_440 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c440
+ bl_0_440 br_0_440 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c440
+ bl_0_440 br_0_440 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c440
+ bl_0_440 br_0_440 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c440
+ bl_0_440 br_0_440 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c440
+ bl_0_440 br_0_440 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c440
+ bl_0_440 br_0_440 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c440
+ bl_0_440 br_0_440 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c440
+ bl_0_440 br_0_440 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c440
+ bl_0_440 br_0_440 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c440
+ bl_0_440 br_0_440 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c440
+ bl_0_440 br_0_440 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c440
+ bl_0_440 br_0_440 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c440
+ bl_0_440 br_0_440 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c440
+ bl_0_440 br_0_440 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c440
+ bl_0_440 br_0_440 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c440
+ bl_0_440 br_0_440 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c440
+ bl_0_440 br_0_440 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c440
+ bl_0_440 br_0_440 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c440
+ bl_0_440 br_0_440 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c440
+ bl_0_440 br_0_440 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c440
+ bl_0_440 br_0_440 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c440
+ bl_0_440 br_0_440 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c440
+ bl_0_440 br_0_440 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c440
+ bl_0_440 br_0_440 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c440
+ bl_0_440 br_0_440 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c440
+ bl_0_440 br_0_440 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c441
+ bl_0_441 br_0_441 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c441
+ bl_0_441 br_0_441 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c441
+ bl_0_441 br_0_441 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c441
+ bl_0_441 br_0_441 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c441
+ bl_0_441 br_0_441 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c441
+ bl_0_441 br_0_441 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c441
+ bl_0_441 br_0_441 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c441
+ bl_0_441 br_0_441 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c441
+ bl_0_441 br_0_441 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c441
+ bl_0_441 br_0_441 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c441
+ bl_0_441 br_0_441 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c441
+ bl_0_441 br_0_441 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c441
+ bl_0_441 br_0_441 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c441
+ bl_0_441 br_0_441 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c441
+ bl_0_441 br_0_441 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c441
+ bl_0_441 br_0_441 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c441
+ bl_0_441 br_0_441 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c441
+ bl_0_441 br_0_441 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c441
+ bl_0_441 br_0_441 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c441
+ bl_0_441 br_0_441 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c441
+ bl_0_441 br_0_441 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c441
+ bl_0_441 br_0_441 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c441
+ bl_0_441 br_0_441 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c441
+ bl_0_441 br_0_441 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c441
+ bl_0_441 br_0_441 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c441
+ bl_0_441 br_0_441 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c441
+ bl_0_441 br_0_441 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c441
+ bl_0_441 br_0_441 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c441
+ bl_0_441 br_0_441 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c441
+ bl_0_441 br_0_441 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c441
+ bl_0_441 br_0_441 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c441
+ bl_0_441 br_0_441 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c441
+ bl_0_441 br_0_441 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c441
+ bl_0_441 br_0_441 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c441
+ bl_0_441 br_0_441 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c441
+ bl_0_441 br_0_441 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c441
+ bl_0_441 br_0_441 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c441
+ bl_0_441 br_0_441 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c441
+ bl_0_441 br_0_441 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c441
+ bl_0_441 br_0_441 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c441
+ bl_0_441 br_0_441 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c441
+ bl_0_441 br_0_441 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c441
+ bl_0_441 br_0_441 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c441
+ bl_0_441 br_0_441 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c441
+ bl_0_441 br_0_441 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c442
+ bl_0_442 br_0_442 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c442
+ bl_0_442 br_0_442 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c442
+ bl_0_442 br_0_442 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c442
+ bl_0_442 br_0_442 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c442
+ bl_0_442 br_0_442 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c442
+ bl_0_442 br_0_442 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c442
+ bl_0_442 br_0_442 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c442
+ bl_0_442 br_0_442 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c442
+ bl_0_442 br_0_442 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c442
+ bl_0_442 br_0_442 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c442
+ bl_0_442 br_0_442 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c442
+ bl_0_442 br_0_442 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c442
+ bl_0_442 br_0_442 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c442
+ bl_0_442 br_0_442 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c442
+ bl_0_442 br_0_442 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c442
+ bl_0_442 br_0_442 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c442
+ bl_0_442 br_0_442 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c442
+ bl_0_442 br_0_442 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c442
+ bl_0_442 br_0_442 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c442
+ bl_0_442 br_0_442 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c442
+ bl_0_442 br_0_442 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c442
+ bl_0_442 br_0_442 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c442
+ bl_0_442 br_0_442 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c442
+ bl_0_442 br_0_442 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c442
+ bl_0_442 br_0_442 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c442
+ bl_0_442 br_0_442 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c442
+ bl_0_442 br_0_442 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c442
+ bl_0_442 br_0_442 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c442
+ bl_0_442 br_0_442 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c442
+ bl_0_442 br_0_442 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c442
+ bl_0_442 br_0_442 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c442
+ bl_0_442 br_0_442 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c442
+ bl_0_442 br_0_442 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c442
+ bl_0_442 br_0_442 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c442
+ bl_0_442 br_0_442 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c442
+ bl_0_442 br_0_442 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c442
+ bl_0_442 br_0_442 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c442
+ bl_0_442 br_0_442 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c442
+ bl_0_442 br_0_442 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c442
+ bl_0_442 br_0_442 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c442
+ bl_0_442 br_0_442 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c442
+ bl_0_442 br_0_442 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c442
+ bl_0_442 br_0_442 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c442
+ bl_0_442 br_0_442 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c442
+ bl_0_442 br_0_442 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c443
+ bl_0_443 br_0_443 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c443
+ bl_0_443 br_0_443 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c443
+ bl_0_443 br_0_443 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c443
+ bl_0_443 br_0_443 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c443
+ bl_0_443 br_0_443 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c443
+ bl_0_443 br_0_443 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c443
+ bl_0_443 br_0_443 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c443
+ bl_0_443 br_0_443 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c443
+ bl_0_443 br_0_443 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c443
+ bl_0_443 br_0_443 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c443
+ bl_0_443 br_0_443 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c443
+ bl_0_443 br_0_443 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c443
+ bl_0_443 br_0_443 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c443
+ bl_0_443 br_0_443 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c443
+ bl_0_443 br_0_443 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c443
+ bl_0_443 br_0_443 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c443
+ bl_0_443 br_0_443 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c443
+ bl_0_443 br_0_443 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c443
+ bl_0_443 br_0_443 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c443
+ bl_0_443 br_0_443 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c443
+ bl_0_443 br_0_443 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c443
+ bl_0_443 br_0_443 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c443
+ bl_0_443 br_0_443 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c443
+ bl_0_443 br_0_443 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c443
+ bl_0_443 br_0_443 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c443
+ bl_0_443 br_0_443 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c443
+ bl_0_443 br_0_443 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c443
+ bl_0_443 br_0_443 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c443
+ bl_0_443 br_0_443 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c443
+ bl_0_443 br_0_443 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c443
+ bl_0_443 br_0_443 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c443
+ bl_0_443 br_0_443 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c443
+ bl_0_443 br_0_443 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c443
+ bl_0_443 br_0_443 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c443
+ bl_0_443 br_0_443 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c443
+ bl_0_443 br_0_443 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c443
+ bl_0_443 br_0_443 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c443
+ bl_0_443 br_0_443 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c443
+ bl_0_443 br_0_443 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c443
+ bl_0_443 br_0_443 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c443
+ bl_0_443 br_0_443 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c443
+ bl_0_443 br_0_443 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c443
+ bl_0_443 br_0_443 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c443
+ bl_0_443 br_0_443 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c443
+ bl_0_443 br_0_443 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c444
+ bl_0_444 br_0_444 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c444
+ bl_0_444 br_0_444 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c444
+ bl_0_444 br_0_444 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c444
+ bl_0_444 br_0_444 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c444
+ bl_0_444 br_0_444 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c444
+ bl_0_444 br_0_444 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c444
+ bl_0_444 br_0_444 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c444
+ bl_0_444 br_0_444 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c444
+ bl_0_444 br_0_444 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c444
+ bl_0_444 br_0_444 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c444
+ bl_0_444 br_0_444 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c444
+ bl_0_444 br_0_444 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c444
+ bl_0_444 br_0_444 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c444
+ bl_0_444 br_0_444 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c444
+ bl_0_444 br_0_444 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c444
+ bl_0_444 br_0_444 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c444
+ bl_0_444 br_0_444 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c444
+ bl_0_444 br_0_444 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c444
+ bl_0_444 br_0_444 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c444
+ bl_0_444 br_0_444 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c444
+ bl_0_444 br_0_444 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c444
+ bl_0_444 br_0_444 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c444
+ bl_0_444 br_0_444 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c444
+ bl_0_444 br_0_444 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c444
+ bl_0_444 br_0_444 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c444
+ bl_0_444 br_0_444 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c444
+ bl_0_444 br_0_444 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c444
+ bl_0_444 br_0_444 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c444
+ bl_0_444 br_0_444 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c444
+ bl_0_444 br_0_444 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c444
+ bl_0_444 br_0_444 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c444
+ bl_0_444 br_0_444 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c444
+ bl_0_444 br_0_444 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c444
+ bl_0_444 br_0_444 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c444
+ bl_0_444 br_0_444 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c444
+ bl_0_444 br_0_444 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c444
+ bl_0_444 br_0_444 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c444
+ bl_0_444 br_0_444 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c444
+ bl_0_444 br_0_444 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c444
+ bl_0_444 br_0_444 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c444
+ bl_0_444 br_0_444 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c444
+ bl_0_444 br_0_444 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c444
+ bl_0_444 br_0_444 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c444
+ bl_0_444 br_0_444 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c444
+ bl_0_444 br_0_444 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c445
+ bl_0_445 br_0_445 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c445
+ bl_0_445 br_0_445 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c445
+ bl_0_445 br_0_445 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c445
+ bl_0_445 br_0_445 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c445
+ bl_0_445 br_0_445 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c445
+ bl_0_445 br_0_445 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c445
+ bl_0_445 br_0_445 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c445
+ bl_0_445 br_0_445 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c445
+ bl_0_445 br_0_445 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c445
+ bl_0_445 br_0_445 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c445
+ bl_0_445 br_0_445 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c445
+ bl_0_445 br_0_445 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c445
+ bl_0_445 br_0_445 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c445
+ bl_0_445 br_0_445 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c445
+ bl_0_445 br_0_445 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c445
+ bl_0_445 br_0_445 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c445
+ bl_0_445 br_0_445 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c445
+ bl_0_445 br_0_445 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c445
+ bl_0_445 br_0_445 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c445
+ bl_0_445 br_0_445 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c445
+ bl_0_445 br_0_445 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c445
+ bl_0_445 br_0_445 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c445
+ bl_0_445 br_0_445 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c445
+ bl_0_445 br_0_445 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c445
+ bl_0_445 br_0_445 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c445
+ bl_0_445 br_0_445 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c445
+ bl_0_445 br_0_445 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c445
+ bl_0_445 br_0_445 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c445
+ bl_0_445 br_0_445 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c445
+ bl_0_445 br_0_445 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c445
+ bl_0_445 br_0_445 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c445
+ bl_0_445 br_0_445 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c445
+ bl_0_445 br_0_445 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c445
+ bl_0_445 br_0_445 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c445
+ bl_0_445 br_0_445 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c445
+ bl_0_445 br_0_445 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c445
+ bl_0_445 br_0_445 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c445
+ bl_0_445 br_0_445 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c445
+ bl_0_445 br_0_445 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c445
+ bl_0_445 br_0_445 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c445
+ bl_0_445 br_0_445 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c445
+ bl_0_445 br_0_445 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c445
+ bl_0_445 br_0_445 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c445
+ bl_0_445 br_0_445 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c445
+ bl_0_445 br_0_445 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c446
+ bl_0_446 br_0_446 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c446
+ bl_0_446 br_0_446 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c446
+ bl_0_446 br_0_446 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c446
+ bl_0_446 br_0_446 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c446
+ bl_0_446 br_0_446 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c446
+ bl_0_446 br_0_446 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c446
+ bl_0_446 br_0_446 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c446
+ bl_0_446 br_0_446 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c446
+ bl_0_446 br_0_446 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c446
+ bl_0_446 br_0_446 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c446
+ bl_0_446 br_0_446 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c446
+ bl_0_446 br_0_446 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c446
+ bl_0_446 br_0_446 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c446
+ bl_0_446 br_0_446 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c446
+ bl_0_446 br_0_446 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c446
+ bl_0_446 br_0_446 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c446
+ bl_0_446 br_0_446 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c446
+ bl_0_446 br_0_446 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c446
+ bl_0_446 br_0_446 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c446
+ bl_0_446 br_0_446 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c446
+ bl_0_446 br_0_446 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c446
+ bl_0_446 br_0_446 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c446
+ bl_0_446 br_0_446 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c446
+ bl_0_446 br_0_446 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c446
+ bl_0_446 br_0_446 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c446
+ bl_0_446 br_0_446 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c446
+ bl_0_446 br_0_446 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c446
+ bl_0_446 br_0_446 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c446
+ bl_0_446 br_0_446 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c446
+ bl_0_446 br_0_446 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c446
+ bl_0_446 br_0_446 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c446
+ bl_0_446 br_0_446 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c446
+ bl_0_446 br_0_446 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c446
+ bl_0_446 br_0_446 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c446
+ bl_0_446 br_0_446 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c446
+ bl_0_446 br_0_446 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c446
+ bl_0_446 br_0_446 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c446
+ bl_0_446 br_0_446 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c446
+ bl_0_446 br_0_446 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c446
+ bl_0_446 br_0_446 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c446
+ bl_0_446 br_0_446 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c446
+ bl_0_446 br_0_446 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c446
+ bl_0_446 br_0_446 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c446
+ bl_0_446 br_0_446 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c446
+ bl_0_446 br_0_446 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c447
+ bl_0_447 br_0_447 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c447
+ bl_0_447 br_0_447 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c447
+ bl_0_447 br_0_447 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c447
+ bl_0_447 br_0_447 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c447
+ bl_0_447 br_0_447 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c447
+ bl_0_447 br_0_447 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c447
+ bl_0_447 br_0_447 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c447
+ bl_0_447 br_0_447 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c447
+ bl_0_447 br_0_447 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c447
+ bl_0_447 br_0_447 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c447
+ bl_0_447 br_0_447 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c447
+ bl_0_447 br_0_447 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c447
+ bl_0_447 br_0_447 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c447
+ bl_0_447 br_0_447 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c447
+ bl_0_447 br_0_447 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c447
+ bl_0_447 br_0_447 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c447
+ bl_0_447 br_0_447 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c447
+ bl_0_447 br_0_447 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c447
+ bl_0_447 br_0_447 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c447
+ bl_0_447 br_0_447 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c447
+ bl_0_447 br_0_447 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c447
+ bl_0_447 br_0_447 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c447
+ bl_0_447 br_0_447 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c447
+ bl_0_447 br_0_447 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c447
+ bl_0_447 br_0_447 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c447
+ bl_0_447 br_0_447 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c447
+ bl_0_447 br_0_447 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c447
+ bl_0_447 br_0_447 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c447
+ bl_0_447 br_0_447 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c447
+ bl_0_447 br_0_447 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c447
+ bl_0_447 br_0_447 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c447
+ bl_0_447 br_0_447 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c447
+ bl_0_447 br_0_447 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c447
+ bl_0_447 br_0_447 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c447
+ bl_0_447 br_0_447 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c447
+ bl_0_447 br_0_447 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c447
+ bl_0_447 br_0_447 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c447
+ bl_0_447 br_0_447 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c447
+ bl_0_447 br_0_447 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c447
+ bl_0_447 br_0_447 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c447
+ bl_0_447 br_0_447 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c447
+ bl_0_447 br_0_447 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c447
+ bl_0_447 br_0_447 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c447
+ bl_0_447 br_0_447 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c447
+ bl_0_447 br_0_447 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c448
+ bl_0_448 br_0_448 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c448
+ bl_0_448 br_0_448 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c448
+ bl_0_448 br_0_448 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c448
+ bl_0_448 br_0_448 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c448
+ bl_0_448 br_0_448 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c448
+ bl_0_448 br_0_448 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c448
+ bl_0_448 br_0_448 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c448
+ bl_0_448 br_0_448 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c448
+ bl_0_448 br_0_448 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c448
+ bl_0_448 br_0_448 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c448
+ bl_0_448 br_0_448 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c448
+ bl_0_448 br_0_448 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c448
+ bl_0_448 br_0_448 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c448
+ bl_0_448 br_0_448 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c448
+ bl_0_448 br_0_448 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c448
+ bl_0_448 br_0_448 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c448
+ bl_0_448 br_0_448 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c448
+ bl_0_448 br_0_448 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c448
+ bl_0_448 br_0_448 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c448
+ bl_0_448 br_0_448 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c448
+ bl_0_448 br_0_448 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c448
+ bl_0_448 br_0_448 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c448
+ bl_0_448 br_0_448 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c448
+ bl_0_448 br_0_448 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c448
+ bl_0_448 br_0_448 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c448
+ bl_0_448 br_0_448 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c448
+ bl_0_448 br_0_448 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c448
+ bl_0_448 br_0_448 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c448
+ bl_0_448 br_0_448 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c448
+ bl_0_448 br_0_448 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c448
+ bl_0_448 br_0_448 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c448
+ bl_0_448 br_0_448 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c448
+ bl_0_448 br_0_448 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c448
+ bl_0_448 br_0_448 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c448
+ bl_0_448 br_0_448 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c448
+ bl_0_448 br_0_448 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c448
+ bl_0_448 br_0_448 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c448
+ bl_0_448 br_0_448 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c448
+ bl_0_448 br_0_448 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c448
+ bl_0_448 br_0_448 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c448
+ bl_0_448 br_0_448 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c448
+ bl_0_448 br_0_448 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c448
+ bl_0_448 br_0_448 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c448
+ bl_0_448 br_0_448 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c448
+ bl_0_448 br_0_448 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c449
+ bl_0_449 br_0_449 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c449
+ bl_0_449 br_0_449 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c449
+ bl_0_449 br_0_449 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c449
+ bl_0_449 br_0_449 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c449
+ bl_0_449 br_0_449 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c449
+ bl_0_449 br_0_449 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c449
+ bl_0_449 br_0_449 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c449
+ bl_0_449 br_0_449 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c449
+ bl_0_449 br_0_449 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c449
+ bl_0_449 br_0_449 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c449
+ bl_0_449 br_0_449 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c449
+ bl_0_449 br_0_449 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c449
+ bl_0_449 br_0_449 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c449
+ bl_0_449 br_0_449 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c449
+ bl_0_449 br_0_449 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c449
+ bl_0_449 br_0_449 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c449
+ bl_0_449 br_0_449 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c449
+ bl_0_449 br_0_449 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c449
+ bl_0_449 br_0_449 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c449
+ bl_0_449 br_0_449 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c449
+ bl_0_449 br_0_449 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c449
+ bl_0_449 br_0_449 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c449
+ bl_0_449 br_0_449 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c449
+ bl_0_449 br_0_449 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c449
+ bl_0_449 br_0_449 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c449
+ bl_0_449 br_0_449 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c449
+ bl_0_449 br_0_449 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c449
+ bl_0_449 br_0_449 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c449
+ bl_0_449 br_0_449 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c449
+ bl_0_449 br_0_449 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c449
+ bl_0_449 br_0_449 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c449
+ bl_0_449 br_0_449 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c449
+ bl_0_449 br_0_449 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c449
+ bl_0_449 br_0_449 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c449
+ bl_0_449 br_0_449 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c449
+ bl_0_449 br_0_449 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c449
+ bl_0_449 br_0_449 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c449
+ bl_0_449 br_0_449 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c449
+ bl_0_449 br_0_449 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c449
+ bl_0_449 br_0_449 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c449
+ bl_0_449 br_0_449 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c449
+ bl_0_449 br_0_449 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c449
+ bl_0_449 br_0_449 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c449
+ bl_0_449 br_0_449 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c449
+ bl_0_449 br_0_449 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c450
+ bl_0_450 br_0_450 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c450
+ bl_0_450 br_0_450 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c450
+ bl_0_450 br_0_450 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c450
+ bl_0_450 br_0_450 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c450
+ bl_0_450 br_0_450 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c450
+ bl_0_450 br_0_450 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c450
+ bl_0_450 br_0_450 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c450
+ bl_0_450 br_0_450 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c450
+ bl_0_450 br_0_450 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c450
+ bl_0_450 br_0_450 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c450
+ bl_0_450 br_0_450 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c450
+ bl_0_450 br_0_450 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c450
+ bl_0_450 br_0_450 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c450
+ bl_0_450 br_0_450 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c450
+ bl_0_450 br_0_450 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c450
+ bl_0_450 br_0_450 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c450
+ bl_0_450 br_0_450 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c450
+ bl_0_450 br_0_450 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c450
+ bl_0_450 br_0_450 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c450
+ bl_0_450 br_0_450 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c450
+ bl_0_450 br_0_450 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c450
+ bl_0_450 br_0_450 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c450
+ bl_0_450 br_0_450 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c450
+ bl_0_450 br_0_450 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c450
+ bl_0_450 br_0_450 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c450
+ bl_0_450 br_0_450 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c450
+ bl_0_450 br_0_450 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c450
+ bl_0_450 br_0_450 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c450
+ bl_0_450 br_0_450 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c450
+ bl_0_450 br_0_450 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c450
+ bl_0_450 br_0_450 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c450
+ bl_0_450 br_0_450 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c450
+ bl_0_450 br_0_450 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c450
+ bl_0_450 br_0_450 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c450
+ bl_0_450 br_0_450 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c450
+ bl_0_450 br_0_450 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c450
+ bl_0_450 br_0_450 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c450
+ bl_0_450 br_0_450 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c450
+ bl_0_450 br_0_450 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c450
+ bl_0_450 br_0_450 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c450
+ bl_0_450 br_0_450 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c450
+ bl_0_450 br_0_450 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c450
+ bl_0_450 br_0_450 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c450
+ bl_0_450 br_0_450 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c450
+ bl_0_450 br_0_450 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c451
+ bl_0_451 br_0_451 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c451
+ bl_0_451 br_0_451 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c451
+ bl_0_451 br_0_451 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c451
+ bl_0_451 br_0_451 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c451
+ bl_0_451 br_0_451 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c451
+ bl_0_451 br_0_451 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c451
+ bl_0_451 br_0_451 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c451
+ bl_0_451 br_0_451 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c451
+ bl_0_451 br_0_451 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c451
+ bl_0_451 br_0_451 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c451
+ bl_0_451 br_0_451 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c451
+ bl_0_451 br_0_451 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c451
+ bl_0_451 br_0_451 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c451
+ bl_0_451 br_0_451 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c451
+ bl_0_451 br_0_451 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c451
+ bl_0_451 br_0_451 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c451
+ bl_0_451 br_0_451 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c451
+ bl_0_451 br_0_451 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c451
+ bl_0_451 br_0_451 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c451
+ bl_0_451 br_0_451 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c451
+ bl_0_451 br_0_451 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c451
+ bl_0_451 br_0_451 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c451
+ bl_0_451 br_0_451 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c451
+ bl_0_451 br_0_451 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c451
+ bl_0_451 br_0_451 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c451
+ bl_0_451 br_0_451 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c451
+ bl_0_451 br_0_451 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c451
+ bl_0_451 br_0_451 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c451
+ bl_0_451 br_0_451 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c451
+ bl_0_451 br_0_451 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c451
+ bl_0_451 br_0_451 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c451
+ bl_0_451 br_0_451 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c451
+ bl_0_451 br_0_451 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c451
+ bl_0_451 br_0_451 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c451
+ bl_0_451 br_0_451 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c451
+ bl_0_451 br_0_451 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c451
+ bl_0_451 br_0_451 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c451
+ bl_0_451 br_0_451 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c451
+ bl_0_451 br_0_451 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c451
+ bl_0_451 br_0_451 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c451
+ bl_0_451 br_0_451 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c451
+ bl_0_451 br_0_451 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c451
+ bl_0_451 br_0_451 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c451
+ bl_0_451 br_0_451 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c451
+ bl_0_451 br_0_451 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c452
+ bl_0_452 br_0_452 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c452
+ bl_0_452 br_0_452 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c452
+ bl_0_452 br_0_452 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c452
+ bl_0_452 br_0_452 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c452
+ bl_0_452 br_0_452 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c452
+ bl_0_452 br_0_452 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c452
+ bl_0_452 br_0_452 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c452
+ bl_0_452 br_0_452 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c452
+ bl_0_452 br_0_452 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c452
+ bl_0_452 br_0_452 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c452
+ bl_0_452 br_0_452 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c452
+ bl_0_452 br_0_452 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c452
+ bl_0_452 br_0_452 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c452
+ bl_0_452 br_0_452 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c452
+ bl_0_452 br_0_452 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c452
+ bl_0_452 br_0_452 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c452
+ bl_0_452 br_0_452 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c452
+ bl_0_452 br_0_452 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c452
+ bl_0_452 br_0_452 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c452
+ bl_0_452 br_0_452 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c452
+ bl_0_452 br_0_452 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c452
+ bl_0_452 br_0_452 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c452
+ bl_0_452 br_0_452 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c452
+ bl_0_452 br_0_452 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c452
+ bl_0_452 br_0_452 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c452
+ bl_0_452 br_0_452 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c452
+ bl_0_452 br_0_452 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c452
+ bl_0_452 br_0_452 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c452
+ bl_0_452 br_0_452 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c452
+ bl_0_452 br_0_452 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c452
+ bl_0_452 br_0_452 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c452
+ bl_0_452 br_0_452 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c452
+ bl_0_452 br_0_452 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c452
+ bl_0_452 br_0_452 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c452
+ bl_0_452 br_0_452 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c452
+ bl_0_452 br_0_452 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c452
+ bl_0_452 br_0_452 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c452
+ bl_0_452 br_0_452 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c452
+ bl_0_452 br_0_452 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c452
+ bl_0_452 br_0_452 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c452
+ bl_0_452 br_0_452 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c452
+ bl_0_452 br_0_452 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c452
+ bl_0_452 br_0_452 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c452
+ bl_0_452 br_0_452 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c452
+ bl_0_452 br_0_452 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c453
+ bl_0_453 br_0_453 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c453
+ bl_0_453 br_0_453 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c453
+ bl_0_453 br_0_453 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c453
+ bl_0_453 br_0_453 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c453
+ bl_0_453 br_0_453 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c453
+ bl_0_453 br_0_453 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c453
+ bl_0_453 br_0_453 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c453
+ bl_0_453 br_0_453 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c453
+ bl_0_453 br_0_453 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c453
+ bl_0_453 br_0_453 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c453
+ bl_0_453 br_0_453 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c453
+ bl_0_453 br_0_453 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c453
+ bl_0_453 br_0_453 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c453
+ bl_0_453 br_0_453 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c453
+ bl_0_453 br_0_453 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c453
+ bl_0_453 br_0_453 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c453
+ bl_0_453 br_0_453 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c453
+ bl_0_453 br_0_453 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c453
+ bl_0_453 br_0_453 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c453
+ bl_0_453 br_0_453 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c453
+ bl_0_453 br_0_453 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c453
+ bl_0_453 br_0_453 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c453
+ bl_0_453 br_0_453 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c453
+ bl_0_453 br_0_453 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c453
+ bl_0_453 br_0_453 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c453
+ bl_0_453 br_0_453 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c453
+ bl_0_453 br_0_453 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c453
+ bl_0_453 br_0_453 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c453
+ bl_0_453 br_0_453 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c453
+ bl_0_453 br_0_453 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c453
+ bl_0_453 br_0_453 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c453
+ bl_0_453 br_0_453 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c453
+ bl_0_453 br_0_453 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c453
+ bl_0_453 br_0_453 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c453
+ bl_0_453 br_0_453 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c453
+ bl_0_453 br_0_453 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c453
+ bl_0_453 br_0_453 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c453
+ bl_0_453 br_0_453 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c453
+ bl_0_453 br_0_453 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c453
+ bl_0_453 br_0_453 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c453
+ bl_0_453 br_0_453 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c453
+ bl_0_453 br_0_453 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c453
+ bl_0_453 br_0_453 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c453
+ bl_0_453 br_0_453 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c453
+ bl_0_453 br_0_453 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c454
+ bl_0_454 br_0_454 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c454
+ bl_0_454 br_0_454 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c454
+ bl_0_454 br_0_454 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c454
+ bl_0_454 br_0_454 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c454
+ bl_0_454 br_0_454 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c454
+ bl_0_454 br_0_454 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c454
+ bl_0_454 br_0_454 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c454
+ bl_0_454 br_0_454 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c454
+ bl_0_454 br_0_454 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c454
+ bl_0_454 br_0_454 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c454
+ bl_0_454 br_0_454 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c454
+ bl_0_454 br_0_454 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c454
+ bl_0_454 br_0_454 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c454
+ bl_0_454 br_0_454 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c454
+ bl_0_454 br_0_454 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c454
+ bl_0_454 br_0_454 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c454
+ bl_0_454 br_0_454 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c454
+ bl_0_454 br_0_454 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c454
+ bl_0_454 br_0_454 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c454
+ bl_0_454 br_0_454 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c454
+ bl_0_454 br_0_454 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c454
+ bl_0_454 br_0_454 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c454
+ bl_0_454 br_0_454 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c454
+ bl_0_454 br_0_454 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c454
+ bl_0_454 br_0_454 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c454
+ bl_0_454 br_0_454 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c454
+ bl_0_454 br_0_454 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c454
+ bl_0_454 br_0_454 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c454
+ bl_0_454 br_0_454 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c454
+ bl_0_454 br_0_454 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c454
+ bl_0_454 br_0_454 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c454
+ bl_0_454 br_0_454 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c454
+ bl_0_454 br_0_454 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c454
+ bl_0_454 br_0_454 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c454
+ bl_0_454 br_0_454 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c454
+ bl_0_454 br_0_454 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c454
+ bl_0_454 br_0_454 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c454
+ bl_0_454 br_0_454 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c454
+ bl_0_454 br_0_454 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c454
+ bl_0_454 br_0_454 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c454
+ bl_0_454 br_0_454 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c454
+ bl_0_454 br_0_454 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c454
+ bl_0_454 br_0_454 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c454
+ bl_0_454 br_0_454 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c454
+ bl_0_454 br_0_454 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c455
+ bl_0_455 br_0_455 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c455
+ bl_0_455 br_0_455 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c455
+ bl_0_455 br_0_455 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c455
+ bl_0_455 br_0_455 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c455
+ bl_0_455 br_0_455 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c455
+ bl_0_455 br_0_455 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c455
+ bl_0_455 br_0_455 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c455
+ bl_0_455 br_0_455 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c455
+ bl_0_455 br_0_455 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c455
+ bl_0_455 br_0_455 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c455
+ bl_0_455 br_0_455 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c455
+ bl_0_455 br_0_455 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c455
+ bl_0_455 br_0_455 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c455
+ bl_0_455 br_0_455 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c455
+ bl_0_455 br_0_455 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c455
+ bl_0_455 br_0_455 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c455
+ bl_0_455 br_0_455 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c455
+ bl_0_455 br_0_455 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c455
+ bl_0_455 br_0_455 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c455
+ bl_0_455 br_0_455 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c455
+ bl_0_455 br_0_455 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c455
+ bl_0_455 br_0_455 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c455
+ bl_0_455 br_0_455 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c455
+ bl_0_455 br_0_455 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c455
+ bl_0_455 br_0_455 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c455
+ bl_0_455 br_0_455 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c455
+ bl_0_455 br_0_455 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c455
+ bl_0_455 br_0_455 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c455
+ bl_0_455 br_0_455 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c455
+ bl_0_455 br_0_455 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c455
+ bl_0_455 br_0_455 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c455
+ bl_0_455 br_0_455 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c455
+ bl_0_455 br_0_455 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c455
+ bl_0_455 br_0_455 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c455
+ bl_0_455 br_0_455 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c455
+ bl_0_455 br_0_455 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c455
+ bl_0_455 br_0_455 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c455
+ bl_0_455 br_0_455 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c455
+ bl_0_455 br_0_455 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c455
+ bl_0_455 br_0_455 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c455
+ bl_0_455 br_0_455 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c455
+ bl_0_455 br_0_455 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c455
+ bl_0_455 br_0_455 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c455
+ bl_0_455 br_0_455 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c455
+ bl_0_455 br_0_455 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c456
+ bl_0_456 br_0_456 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c456
+ bl_0_456 br_0_456 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c456
+ bl_0_456 br_0_456 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c456
+ bl_0_456 br_0_456 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c456
+ bl_0_456 br_0_456 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c456
+ bl_0_456 br_0_456 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c456
+ bl_0_456 br_0_456 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c456
+ bl_0_456 br_0_456 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c456
+ bl_0_456 br_0_456 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c456
+ bl_0_456 br_0_456 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c456
+ bl_0_456 br_0_456 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c456
+ bl_0_456 br_0_456 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c456
+ bl_0_456 br_0_456 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c456
+ bl_0_456 br_0_456 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c456
+ bl_0_456 br_0_456 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c456
+ bl_0_456 br_0_456 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c456
+ bl_0_456 br_0_456 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c456
+ bl_0_456 br_0_456 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c456
+ bl_0_456 br_0_456 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c456
+ bl_0_456 br_0_456 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c456
+ bl_0_456 br_0_456 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c456
+ bl_0_456 br_0_456 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c456
+ bl_0_456 br_0_456 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c456
+ bl_0_456 br_0_456 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c456
+ bl_0_456 br_0_456 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c456
+ bl_0_456 br_0_456 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c456
+ bl_0_456 br_0_456 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c456
+ bl_0_456 br_0_456 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c456
+ bl_0_456 br_0_456 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c456
+ bl_0_456 br_0_456 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c456
+ bl_0_456 br_0_456 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c456
+ bl_0_456 br_0_456 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c456
+ bl_0_456 br_0_456 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c456
+ bl_0_456 br_0_456 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c456
+ bl_0_456 br_0_456 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c456
+ bl_0_456 br_0_456 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c456
+ bl_0_456 br_0_456 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c456
+ bl_0_456 br_0_456 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c456
+ bl_0_456 br_0_456 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c456
+ bl_0_456 br_0_456 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c456
+ bl_0_456 br_0_456 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c456
+ bl_0_456 br_0_456 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c456
+ bl_0_456 br_0_456 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c456
+ bl_0_456 br_0_456 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c456
+ bl_0_456 br_0_456 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c457
+ bl_0_457 br_0_457 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c457
+ bl_0_457 br_0_457 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c457
+ bl_0_457 br_0_457 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c457
+ bl_0_457 br_0_457 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c457
+ bl_0_457 br_0_457 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c457
+ bl_0_457 br_0_457 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c457
+ bl_0_457 br_0_457 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c457
+ bl_0_457 br_0_457 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c457
+ bl_0_457 br_0_457 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c457
+ bl_0_457 br_0_457 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c457
+ bl_0_457 br_0_457 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c457
+ bl_0_457 br_0_457 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c457
+ bl_0_457 br_0_457 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c457
+ bl_0_457 br_0_457 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c457
+ bl_0_457 br_0_457 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c457
+ bl_0_457 br_0_457 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c457
+ bl_0_457 br_0_457 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c457
+ bl_0_457 br_0_457 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c457
+ bl_0_457 br_0_457 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c457
+ bl_0_457 br_0_457 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c457
+ bl_0_457 br_0_457 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c457
+ bl_0_457 br_0_457 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c457
+ bl_0_457 br_0_457 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c457
+ bl_0_457 br_0_457 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c457
+ bl_0_457 br_0_457 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c457
+ bl_0_457 br_0_457 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c457
+ bl_0_457 br_0_457 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c457
+ bl_0_457 br_0_457 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c457
+ bl_0_457 br_0_457 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c457
+ bl_0_457 br_0_457 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c457
+ bl_0_457 br_0_457 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c457
+ bl_0_457 br_0_457 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c457
+ bl_0_457 br_0_457 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c457
+ bl_0_457 br_0_457 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c457
+ bl_0_457 br_0_457 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c457
+ bl_0_457 br_0_457 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c457
+ bl_0_457 br_0_457 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c457
+ bl_0_457 br_0_457 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c457
+ bl_0_457 br_0_457 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c457
+ bl_0_457 br_0_457 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c457
+ bl_0_457 br_0_457 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c457
+ bl_0_457 br_0_457 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c457
+ bl_0_457 br_0_457 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c457
+ bl_0_457 br_0_457 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c457
+ bl_0_457 br_0_457 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c458
+ bl_0_458 br_0_458 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c458
+ bl_0_458 br_0_458 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c458
+ bl_0_458 br_0_458 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c458
+ bl_0_458 br_0_458 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c458
+ bl_0_458 br_0_458 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c458
+ bl_0_458 br_0_458 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c458
+ bl_0_458 br_0_458 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c458
+ bl_0_458 br_0_458 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c458
+ bl_0_458 br_0_458 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c458
+ bl_0_458 br_0_458 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c458
+ bl_0_458 br_0_458 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c458
+ bl_0_458 br_0_458 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c458
+ bl_0_458 br_0_458 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c458
+ bl_0_458 br_0_458 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c458
+ bl_0_458 br_0_458 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c458
+ bl_0_458 br_0_458 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c458
+ bl_0_458 br_0_458 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c458
+ bl_0_458 br_0_458 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c458
+ bl_0_458 br_0_458 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c458
+ bl_0_458 br_0_458 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c458
+ bl_0_458 br_0_458 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c458
+ bl_0_458 br_0_458 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c458
+ bl_0_458 br_0_458 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c458
+ bl_0_458 br_0_458 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c458
+ bl_0_458 br_0_458 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c458
+ bl_0_458 br_0_458 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c458
+ bl_0_458 br_0_458 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c458
+ bl_0_458 br_0_458 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c458
+ bl_0_458 br_0_458 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c458
+ bl_0_458 br_0_458 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c458
+ bl_0_458 br_0_458 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c458
+ bl_0_458 br_0_458 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c458
+ bl_0_458 br_0_458 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c458
+ bl_0_458 br_0_458 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c458
+ bl_0_458 br_0_458 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c458
+ bl_0_458 br_0_458 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c458
+ bl_0_458 br_0_458 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c458
+ bl_0_458 br_0_458 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c458
+ bl_0_458 br_0_458 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c458
+ bl_0_458 br_0_458 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c458
+ bl_0_458 br_0_458 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c458
+ bl_0_458 br_0_458 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c458
+ bl_0_458 br_0_458 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c458
+ bl_0_458 br_0_458 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c458
+ bl_0_458 br_0_458 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c459
+ bl_0_459 br_0_459 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c459
+ bl_0_459 br_0_459 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c459
+ bl_0_459 br_0_459 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c459
+ bl_0_459 br_0_459 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c459
+ bl_0_459 br_0_459 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c459
+ bl_0_459 br_0_459 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c459
+ bl_0_459 br_0_459 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c459
+ bl_0_459 br_0_459 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c459
+ bl_0_459 br_0_459 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c459
+ bl_0_459 br_0_459 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c459
+ bl_0_459 br_0_459 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c459
+ bl_0_459 br_0_459 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c459
+ bl_0_459 br_0_459 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c459
+ bl_0_459 br_0_459 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c459
+ bl_0_459 br_0_459 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c459
+ bl_0_459 br_0_459 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c459
+ bl_0_459 br_0_459 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c459
+ bl_0_459 br_0_459 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c459
+ bl_0_459 br_0_459 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c459
+ bl_0_459 br_0_459 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c459
+ bl_0_459 br_0_459 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c459
+ bl_0_459 br_0_459 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c459
+ bl_0_459 br_0_459 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c459
+ bl_0_459 br_0_459 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c459
+ bl_0_459 br_0_459 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c459
+ bl_0_459 br_0_459 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c459
+ bl_0_459 br_0_459 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c459
+ bl_0_459 br_0_459 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c459
+ bl_0_459 br_0_459 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c459
+ bl_0_459 br_0_459 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c459
+ bl_0_459 br_0_459 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c459
+ bl_0_459 br_0_459 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c459
+ bl_0_459 br_0_459 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c459
+ bl_0_459 br_0_459 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c459
+ bl_0_459 br_0_459 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c459
+ bl_0_459 br_0_459 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c459
+ bl_0_459 br_0_459 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c459
+ bl_0_459 br_0_459 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c459
+ bl_0_459 br_0_459 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c459
+ bl_0_459 br_0_459 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c459
+ bl_0_459 br_0_459 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c459
+ bl_0_459 br_0_459 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c459
+ bl_0_459 br_0_459 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c459
+ bl_0_459 br_0_459 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c459
+ bl_0_459 br_0_459 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c460
+ bl_0_460 br_0_460 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c460
+ bl_0_460 br_0_460 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c460
+ bl_0_460 br_0_460 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c460
+ bl_0_460 br_0_460 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c460
+ bl_0_460 br_0_460 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c460
+ bl_0_460 br_0_460 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c460
+ bl_0_460 br_0_460 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c460
+ bl_0_460 br_0_460 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c460
+ bl_0_460 br_0_460 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c460
+ bl_0_460 br_0_460 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c460
+ bl_0_460 br_0_460 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c460
+ bl_0_460 br_0_460 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c460
+ bl_0_460 br_0_460 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c460
+ bl_0_460 br_0_460 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c460
+ bl_0_460 br_0_460 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c460
+ bl_0_460 br_0_460 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c460
+ bl_0_460 br_0_460 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c460
+ bl_0_460 br_0_460 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c460
+ bl_0_460 br_0_460 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c460
+ bl_0_460 br_0_460 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c460
+ bl_0_460 br_0_460 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c460
+ bl_0_460 br_0_460 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c460
+ bl_0_460 br_0_460 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c460
+ bl_0_460 br_0_460 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c460
+ bl_0_460 br_0_460 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c460
+ bl_0_460 br_0_460 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c460
+ bl_0_460 br_0_460 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c460
+ bl_0_460 br_0_460 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c460
+ bl_0_460 br_0_460 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c460
+ bl_0_460 br_0_460 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c460
+ bl_0_460 br_0_460 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c460
+ bl_0_460 br_0_460 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c460
+ bl_0_460 br_0_460 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c460
+ bl_0_460 br_0_460 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c460
+ bl_0_460 br_0_460 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c460
+ bl_0_460 br_0_460 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c460
+ bl_0_460 br_0_460 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c460
+ bl_0_460 br_0_460 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c460
+ bl_0_460 br_0_460 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c460
+ bl_0_460 br_0_460 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c460
+ bl_0_460 br_0_460 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c460
+ bl_0_460 br_0_460 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c460
+ bl_0_460 br_0_460 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c460
+ bl_0_460 br_0_460 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c460
+ bl_0_460 br_0_460 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c461
+ bl_0_461 br_0_461 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c461
+ bl_0_461 br_0_461 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c461
+ bl_0_461 br_0_461 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c461
+ bl_0_461 br_0_461 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c461
+ bl_0_461 br_0_461 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c461
+ bl_0_461 br_0_461 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c461
+ bl_0_461 br_0_461 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c461
+ bl_0_461 br_0_461 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c461
+ bl_0_461 br_0_461 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c461
+ bl_0_461 br_0_461 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c461
+ bl_0_461 br_0_461 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c461
+ bl_0_461 br_0_461 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c461
+ bl_0_461 br_0_461 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c461
+ bl_0_461 br_0_461 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c461
+ bl_0_461 br_0_461 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c461
+ bl_0_461 br_0_461 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c461
+ bl_0_461 br_0_461 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c461
+ bl_0_461 br_0_461 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c461
+ bl_0_461 br_0_461 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c461
+ bl_0_461 br_0_461 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c461
+ bl_0_461 br_0_461 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c461
+ bl_0_461 br_0_461 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c461
+ bl_0_461 br_0_461 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c461
+ bl_0_461 br_0_461 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c461
+ bl_0_461 br_0_461 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c461
+ bl_0_461 br_0_461 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c461
+ bl_0_461 br_0_461 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c461
+ bl_0_461 br_0_461 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c461
+ bl_0_461 br_0_461 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c461
+ bl_0_461 br_0_461 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c461
+ bl_0_461 br_0_461 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c461
+ bl_0_461 br_0_461 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c461
+ bl_0_461 br_0_461 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c461
+ bl_0_461 br_0_461 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c461
+ bl_0_461 br_0_461 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c461
+ bl_0_461 br_0_461 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c461
+ bl_0_461 br_0_461 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c461
+ bl_0_461 br_0_461 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c461
+ bl_0_461 br_0_461 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c461
+ bl_0_461 br_0_461 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c461
+ bl_0_461 br_0_461 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c461
+ bl_0_461 br_0_461 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c461
+ bl_0_461 br_0_461 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c461
+ bl_0_461 br_0_461 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c461
+ bl_0_461 br_0_461 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c462
+ bl_0_462 br_0_462 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c462
+ bl_0_462 br_0_462 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c462
+ bl_0_462 br_0_462 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c462
+ bl_0_462 br_0_462 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c462
+ bl_0_462 br_0_462 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c462
+ bl_0_462 br_0_462 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c462
+ bl_0_462 br_0_462 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c462
+ bl_0_462 br_0_462 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c462
+ bl_0_462 br_0_462 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c462
+ bl_0_462 br_0_462 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c462
+ bl_0_462 br_0_462 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c462
+ bl_0_462 br_0_462 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c462
+ bl_0_462 br_0_462 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c462
+ bl_0_462 br_0_462 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c462
+ bl_0_462 br_0_462 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c462
+ bl_0_462 br_0_462 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c462
+ bl_0_462 br_0_462 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c462
+ bl_0_462 br_0_462 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c462
+ bl_0_462 br_0_462 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c462
+ bl_0_462 br_0_462 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c462
+ bl_0_462 br_0_462 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c462
+ bl_0_462 br_0_462 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c462
+ bl_0_462 br_0_462 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c462
+ bl_0_462 br_0_462 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c462
+ bl_0_462 br_0_462 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c462
+ bl_0_462 br_0_462 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c462
+ bl_0_462 br_0_462 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c462
+ bl_0_462 br_0_462 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c462
+ bl_0_462 br_0_462 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c462
+ bl_0_462 br_0_462 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c462
+ bl_0_462 br_0_462 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c462
+ bl_0_462 br_0_462 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c462
+ bl_0_462 br_0_462 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c462
+ bl_0_462 br_0_462 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c462
+ bl_0_462 br_0_462 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c462
+ bl_0_462 br_0_462 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c462
+ bl_0_462 br_0_462 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c462
+ bl_0_462 br_0_462 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c462
+ bl_0_462 br_0_462 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c462
+ bl_0_462 br_0_462 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c462
+ bl_0_462 br_0_462 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c462
+ bl_0_462 br_0_462 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c462
+ bl_0_462 br_0_462 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c462
+ bl_0_462 br_0_462 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c462
+ bl_0_462 br_0_462 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c463
+ bl_0_463 br_0_463 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c463
+ bl_0_463 br_0_463 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c463
+ bl_0_463 br_0_463 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c463
+ bl_0_463 br_0_463 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c463
+ bl_0_463 br_0_463 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c463
+ bl_0_463 br_0_463 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c463
+ bl_0_463 br_0_463 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c463
+ bl_0_463 br_0_463 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c463
+ bl_0_463 br_0_463 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c463
+ bl_0_463 br_0_463 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c463
+ bl_0_463 br_0_463 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c463
+ bl_0_463 br_0_463 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c463
+ bl_0_463 br_0_463 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c463
+ bl_0_463 br_0_463 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c463
+ bl_0_463 br_0_463 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c463
+ bl_0_463 br_0_463 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c463
+ bl_0_463 br_0_463 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c463
+ bl_0_463 br_0_463 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c463
+ bl_0_463 br_0_463 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c463
+ bl_0_463 br_0_463 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c463
+ bl_0_463 br_0_463 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c463
+ bl_0_463 br_0_463 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c463
+ bl_0_463 br_0_463 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c463
+ bl_0_463 br_0_463 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c463
+ bl_0_463 br_0_463 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c463
+ bl_0_463 br_0_463 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c463
+ bl_0_463 br_0_463 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c463
+ bl_0_463 br_0_463 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c463
+ bl_0_463 br_0_463 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c463
+ bl_0_463 br_0_463 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c463
+ bl_0_463 br_0_463 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c463
+ bl_0_463 br_0_463 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c463
+ bl_0_463 br_0_463 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c463
+ bl_0_463 br_0_463 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c463
+ bl_0_463 br_0_463 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c463
+ bl_0_463 br_0_463 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c463
+ bl_0_463 br_0_463 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c463
+ bl_0_463 br_0_463 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c463
+ bl_0_463 br_0_463 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c463
+ bl_0_463 br_0_463 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c463
+ bl_0_463 br_0_463 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c463
+ bl_0_463 br_0_463 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c463
+ bl_0_463 br_0_463 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c463
+ bl_0_463 br_0_463 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c463
+ bl_0_463 br_0_463 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c464
+ bl_0_464 br_0_464 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c464
+ bl_0_464 br_0_464 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c464
+ bl_0_464 br_0_464 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c464
+ bl_0_464 br_0_464 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c464
+ bl_0_464 br_0_464 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c464
+ bl_0_464 br_0_464 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c464
+ bl_0_464 br_0_464 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c464
+ bl_0_464 br_0_464 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c464
+ bl_0_464 br_0_464 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c464
+ bl_0_464 br_0_464 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c464
+ bl_0_464 br_0_464 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c464
+ bl_0_464 br_0_464 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c464
+ bl_0_464 br_0_464 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c464
+ bl_0_464 br_0_464 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c464
+ bl_0_464 br_0_464 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c464
+ bl_0_464 br_0_464 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c464
+ bl_0_464 br_0_464 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c464
+ bl_0_464 br_0_464 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c464
+ bl_0_464 br_0_464 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c464
+ bl_0_464 br_0_464 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c464
+ bl_0_464 br_0_464 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c464
+ bl_0_464 br_0_464 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c464
+ bl_0_464 br_0_464 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c464
+ bl_0_464 br_0_464 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c464
+ bl_0_464 br_0_464 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c464
+ bl_0_464 br_0_464 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c464
+ bl_0_464 br_0_464 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c464
+ bl_0_464 br_0_464 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c464
+ bl_0_464 br_0_464 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c464
+ bl_0_464 br_0_464 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c464
+ bl_0_464 br_0_464 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c464
+ bl_0_464 br_0_464 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c464
+ bl_0_464 br_0_464 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c464
+ bl_0_464 br_0_464 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c464
+ bl_0_464 br_0_464 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c464
+ bl_0_464 br_0_464 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c464
+ bl_0_464 br_0_464 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c464
+ bl_0_464 br_0_464 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c464
+ bl_0_464 br_0_464 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c464
+ bl_0_464 br_0_464 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c464
+ bl_0_464 br_0_464 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c464
+ bl_0_464 br_0_464 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c464
+ bl_0_464 br_0_464 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c464
+ bl_0_464 br_0_464 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c464
+ bl_0_464 br_0_464 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c465
+ bl_0_465 br_0_465 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c465
+ bl_0_465 br_0_465 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c465
+ bl_0_465 br_0_465 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c465
+ bl_0_465 br_0_465 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c465
+ bl_0_465 br_0_465 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c465
+ bl_0_465 br_0_465 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c465
+ bl_0_465 br_0_465 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c465
+ bl_0_465 br_0_465 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c465
+ bl_0_465 br_0_465 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c465
+ bl_0_465 br_0_465 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c465
+ bl_0_465 br_0_465 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c465
+ bl_0_465 br_0_465 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c465
+ bl_0_465 br_0_465 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c465
+ bl_0_465 br_0_465 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c465
+ bl_0_465 br_0_465 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c465
+ bl_0_465 br_0_465 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c465
+ bl_0_465 br_0_465 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c465
+ bl_0_465 br_0_465 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c465
+ bl_0_465 br_0_465 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c465
+ bl_0_465 br_0_465 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c465
+ bl_0_465 br_0_465 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c465
+ bl_0_465 br_0_465 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c465
+ bl_0_465 br_0_465 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c465
+ bl_0_465 br_0_465 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c465
+ bl_0_465 br_0_465 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c465
+ bl_0_465 br_0_465 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c465
+ bl_0_465 br_0_465 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c465
+ bl_0_465 br_0_465 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c465
+ bl_0_465 br_0_465 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c465
+ bl_0_465 br_0_465 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c465
+ bl_0_465 br_0_465 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c465
+ bl_0_465 br_0_465 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c465
+ bl_0_465 br_0_465 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c465
+ bl_0_465 br_0_465 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c465
+ bl_0_465 br_0_465 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c465
+ bl_0_465 br_0_465 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c465
+ bl_0_465 br_0_465 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c465
+ bl_0_465 br_0_465 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c465
+ bl_0_465 br_0_465 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c465
+ bl_0_465 br_0_465 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c465
+ bl_0_465 br_0_465 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c465
+ bl_0_465 br_0_465 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c465
+ bl_0_465 br_0_465 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c465
+ bl_0_465 br_0_465 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c465
+ bl_0_465 br_0_465 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c466
+ bl_0_466 br_0_466 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c466
+ bl_0_466 br_0_466 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c466
+ bl_0_466 br_0_466 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c466
+ bl_0_466 br_0_466 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c466
+ bl_0_466 br_0_466 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c466
+ bl_0_466 br_0_466 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c466
+ bl_0_466 br_0_466 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c466
+ bl_0_466 br_0_466 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c466
+ bl_0_466 br_0_466 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c466
+ bl_0_466 br_0_466 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c466
+ bl_0_466 br_0_466 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c466
+ bl_0_466 br_0_466 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c466
+ bl_0_466 br_0_466 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c466
+ bl_0_466 br_0_466 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c466
+ bl_0_466 br_0_466 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c466
+ bl_0_466 br_0_466 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c466
+ bl_0_466 br_0_466 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c466
+ bl_0_466 br_0_466 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c466
+ bl_0_466 br_0_466 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c466
+ bl_0_466 br_0_466 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c466
+ bl_0_466 br_0_466 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c466
+ bl_0_466 br_0_466 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c466
+ bl_0_466 br_0_466 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c466
+ bl_0_466 br_0_466 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c466
+ bl_0_466 br_0_466 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c466
+ bl_0_466 br_0_466 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c466
+ bl_0_466 br_0_466 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c466
+ bl_0_466 br_0_466 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c466
+ bl_0_466 br_0_466 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c466
+ bl_0_466 br_0_466 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c466
+ bl_0_466 br_0_466 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c466
+ bl_0_466 br_0_466 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c466
+ bl_0_466 br_0_466 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c466
+ bl_0_466 br_0_466 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c466
+ bl_0_466 br_0_466 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c466
+ bl_0_466 br_0_466 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c466
+ bl_0_466 br_0_466 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c466
+ bl_0_466 br_0_466 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c466
+ bl_0_466 br_0_466 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c466
+ bl_0_466 br_0_466 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c466
+ bl_0_466 br_0_466 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c466
+ bl_0_466 br_0_466 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c466
+ bl_0_466 br_0_466 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c466
+ bl_0_466 br_0_466 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c466
+ bl_0_466 br_0_466 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c467
+ bl_0_467 br_0_467 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c467
+ bl_0_467 br_0_467 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c467
+ bl_0_467 br_0_467 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c467
+ bl_0_467 br_0_467 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c467
+ bl_0_467 br_0_467 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c467
+ bl_0_467 br_0_467 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c467
+ bl_0_467 br_0_467 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c467
+ bl_0_467 br_0_467 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c467
+ bl_0_467 br_0_467 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c467
+ bl_0_467 br_0_467 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c467
+ bl_0_467 br_0_467 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c467
+ bl_0_467 br_0_467 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c467
+ bl_0_467 br_0_467 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c467
+ bl_0_467 br_0_467 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c467
+ bl_0_467 br_0_467 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c467
+ bl_0_467 br_0_467 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c467
+ bl_0_467 br_0_467 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c467
+ bl_0_467 br_0_467 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c467
+ bl_0_467 br_0_467 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c467
+ bl_0_467 br_0_467 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c467
+ bl_0_467 br_0_467 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c467
+ bl_0_467 br_0_467 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c467
+ bl_0_467 br_0_467 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c467
+ bl_0_467 br_0_467 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c467
+ bl_0_467 br_0_467 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c467
+ bl_0_467 br_0_467 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c467
+ bl_0_467 br_0_467 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c467
+ bl_0_467 br_0_467 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c467
+ bl_0_467 br_0_467 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c467
+ bl_0_467 br_0_467 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c467
+ bl_0_467 br_0_467 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c467
+ bl_0_467 br_0_467 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c467
+ bl_0_467 br_0_467 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c467
+ bl_0_467 br_0_467 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c467
+ bl_0_467 br_0_467 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c467
+ bl_0_467 br_0_467 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c467
+ bl_0_467 br_0_467 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c467
+ bl_0_467 br_0_467 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c467
+ bl_0_467 br_0_467 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c467
+ bl_0_467 br_0_467 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c467
+ bl_0_467 br_0_467 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c467
+ bl_0_467 br_0_467 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c467
+ bl_0_467 br_0_467 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c467
+ bl_0_467 br_0_467 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c467
+ bl_0_467 br_0_467 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c468
+ bl_0_468 br_0_468 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c468
+ bl_0_468 br_0_468 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c468
+ bl_0_468 br_0_468 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c468
+ bl_0_468 br_0_468 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c468
+ bl_0_468 br_0_468 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c468
+ bl_0_468 br_0_468 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c468
+ bl_0_468 br_0_468 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c468
+ bl_0_468 br_0_468 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c468
+ bl_0_468 br_0_468 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c468
+ bl_0_468 br_0_468 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c468
+ bl_0_468 br_0_468 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c468
+ bl_0_468 br_0_468 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c468
+ bl_0_468 br_0_468 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c468
+ bl_0_468 br_0_468 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c468
+ bl_0_468 br_0_468 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c468
+ bl_0_468 br_0_468 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c468
+ bl_0_468 br_0_468 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c468
+ bl_0_468 br_0_468 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c468
+ bl_0_468 br_0_468 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c468
+ bl_0_468 br_0_468 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c468
+ bl_0_468 br_0_468 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c468
+ bl_0_468 br_0_468 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c468
+ bl_0_468 br_0_468 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c468
+ bl_0_468 br_0_468 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c468
+ bl_0_468 br_0_468 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c468
+ bl_0_468 br_0_468 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c468
+ bl_0_468 br_0_468 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c468
+ bl_0_468 br_0_468 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c468
+ bl_0_468 br_0_468 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c468
+ bl_0_468 br_0_468 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c468
+ bl_0_468 br_0_468 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c468
+ bl_0_468 br_0_468 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c468
+ bl_0_468 br_0_468 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c468
+ bl_0_468 br_0_468 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c468
+ bl_0_468 br_0_468 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c468
+ bl_0_468 br_0_468 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c468
+ bl_0_468 br_0_468 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c468
+ bl_0_468 br_0_468 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c468
+ bl_0_468 br_0_468 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c468
+ bl_0_468 br_0_468 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c468
+ bl_0_468 br_0_468 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c468
+ bl_0_468 br_0_468 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c468
+ bl_0_468 br_0_468 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c468
+ bl_0_468 br_0_468 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c468
+ bl_0_468 br_0_468 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c469
+ bl_0_469 br_0_469 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c469
+ bl_0_469 br_0_469 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c469
+ bl_0_469 br_0_469 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c469
+ bl_0_469 br_0_469 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c469
+ bl_0_469 br_0_469 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c469
+ bl_0_469 br_0_469 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c469
+ bl_0_469 br_0_469 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c469
+ bl_0_469 br_0_469 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c469
+ bl_0_469 br_0_469 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c469
+ bl_0_469 br_0_469 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c469
+ bl_0_469 br_0_469 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c469
+ bl_0_469 br_0_469 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c469
+ bl_0_469 br_0_469 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c469
+ bl_0_469 br_0_469 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c469
+ bl_0_469 br_0_469 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c469
+ bl_0_469 br_0_469 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c469
+ bl_0_469 br_0_469 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c469
+ bl_0_469 br_0_469 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c469
+ bl_0_469 br_0_469 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c469
+ bl_0_469 br_0_469 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c469
+ bl_0_469 br_0_469 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c469
+ bl_0_469 br_0_469 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c469
+ bl_0_469 br_0_469 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c469
+ bl_0_469 br_0_469 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c469
+ bl_0_469 br_0_469 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c469
+ bl_0_469 br_0_469 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c469
+ bl_0_469 br_0_469 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c469
+ bl_0_469 br_0_469 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c469
+ bl_0_469 br_0_469 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c469
+ bl_0_469 br_0_469 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c469
+ bl_0_469 br_0_469 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c469
+ bl_0_469 br_0_469 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c469
+ bl_0_469 br_0_469 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c469
+ bl_0_469 br_0_469 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c469
+ bl_0_469 br_0_469 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c469
+ bl_0_469 br_0_469 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c469
+ bl_0_469 br_0_469 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c469
+ bl_0_469 br_0_469 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c469
+ bl_0_469 br_0_469 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c469
+ bl_0_469 br_0_469 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c469
+ bl_0_469 br_0_469 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c469
+ bl_0_469 br_0_469 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c469
+ bl_0_469 br_0_469 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c469
+ bl_0_469 br_0_469 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c469
+ bl_0_469 br_0_469 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c470
+ bl_0_470 br_0_470 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c470
+ bl_0_470 br_0_470 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c470
+ bl_0_470 br_0_470 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c470
+ bl_0_470 br_0_470 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c470
+ bl_0_470 br_0_470 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c470
+ bl_0_470 br_0_470 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c470
+ bl_0_470 br_0_470 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c470
+ bl_0_470 br_0_470 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c470
+ bl_0_470 br_0_470 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c470
+ bl_0_470 br_0_470 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c470
+ bl_0_470 br_0_470 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c470
+ bl_0_470 br_0_470 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c470
+ bl_0_470 br_0_470 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c470
+ bl_0_470 br_0_470 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c470
+ bl_0_470 br_0_470 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c470
+ bl_0_470 br_0_470 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c470
+ bl_0_470 br_0_470 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c470
+ bl_0_470 br_0_470 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c470
+ bl_0_470 br_0_470 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c470
+ bl_0_470 br_0_470 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c470
+ bl_0_470 br_0_470 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c470
+ bl_0_470 br_0_470 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c470
+ bl_0_470 br_0_470 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c470
+ bl_0_470 br_0_470 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c470
+ bl_0_470 br_0_470 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c470
+ bl_0_470 br_0_470 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c470
+ bl_0_470 br_0_470 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c470
+ bl_0_470 br_0_470 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c470
+ bl_0_470 br_0_470 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c470
+ bl_0_470 br_0_470 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c470
+ bl_0_470 br_0_470 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c470
+ bl_0_470 br_0_470 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c470
+ bl_0_470 br_0_470 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c470
+ bl_0_470 br_0_470 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c470
+ bl_0_470 br_0_470 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c470
+ bl_0_470 br_0_470 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c470
+ bl_0_470 br_0_470 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c470
+ bl_0_470 br_0_470 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c470
+ bl_0_470 br_0_470 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c470
+ bl_0_470 br_0_470 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c470
+ bl_0_470 br_0_470 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c470
+ bl_0_470 br_0_470 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c470
+ bl_0_470 br_0_470 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c470
+ bl_0_470 br_0_470 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c470
+ bl_0_470 br_0_470 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c471
+ bl_0_471 br_0_471 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c471
+ bl_0_471 br_0_471 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c471
+ bl_0_471 br_0_471 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c471
+ bl_0_471 br_0_471 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c471
+ bl_0_471 br_0_471 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c471
+ bl_0_471 br_0_471 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c471
+ bl_0_471 br_0_471 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c471
+ bl_0_471 br_0_471 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c471
+ bl_0_471 br_0_471 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c471
+ bl_0_471 br_0_471 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c471
+ bl_0_471 br_0_471 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c471
+ bl_0_471 br_0_471 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c471
+ bl_0_471 br_0_471 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c471
+ bl_0_471 br_0_471 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c471
+ bl_0_471 br_0_471 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c471
+ bl_0_471 br_0_471 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c471
+ bl_0_471 br_0_471 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c471
+ bl_0_471 br_0_471 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c471
+ bl_0_471 br_0_471 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c471
+ bl_0_471 br_0_471 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c471
+ bl_0_471 br_0_471 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c471
+ bl_0_471 br_0_471 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c471
+ bl_0_471 br_0_471 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c471
+ bl_0_471 br_0_471 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c471
+ bl_0_471 br_0_471 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c471
+ bl_0_471 br_0_471 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c471
+ bl_0_471 br_0_471 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c471
+ bl_0_471 br_0_471 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c471
+ bl_0_471 br_0_471 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c471
+ bl_0_471 br_0_471 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c471
+ bl_0_471 br_0_471 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c471
+ bl_0_471 br_0_471 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c471
+ bl_0_471 br_0_471 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c471
+ bl_0_471 br_0_471 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c471
+ bl_0_471 br_0_471 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c471
+ bl_0_471 br_0_471 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c471
+ bl_0_471 br_0_471 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c471
+ bl_0_471 br_0_471 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c471
+ bl_0_471 br_0_471 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c471
+ bl_0_471 br_0_471 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c471
+ bl_0_471 br_0_471 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c471
+ bl_0_471 br_0_471 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c471
+ bl_0_471 br_0_471 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c471
+ bl_0_471 br_0_471 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c471
+ bl_0_471 br_0_471 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c472
+ bl_0_472 br_0_472 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c472
+ bl_0_472 br_0_472 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c472
+ bl_0_472 br_0_472 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c472
+ bl_0_472 br_0_472 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c472
+ bl_0_472 br_0_472 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c472
+ bl_0_472 br_0_472 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c472
+ bl_0_472 br_0_472 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c472
+ bl_0_472 br_0_472 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c472
+ bl_0_472 br_0_472 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c472
+ bl_0_472 br_0_472 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c472
+ bl_0_472 br_0_472 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c472
+ bl_0_472 br_0_472 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c472
+ bl_0_472 br_0_472 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c472
+ bl_0_472 br_0_472 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c472
+ bl_0_472 br_0_472 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c472
+ bl_0_472 br_0_472 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c472
+ bl_0_472 br_0_472 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c472
+ bl_0_472 br_0_472 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c472
+ bl_0_472 br_0_472 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c472
+ bl_0_472 br_0_472 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c472
+ bl_0_472 br_0_472 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c472
+ bl_0_472 br_0_472 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c472
+ bl_0_472 br_0_472 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c472
+ bl_0_472 br_0_472 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c472
+ bl_0_472 br_0_472 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c472
+ bl_0_472 br_0_472 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c472
+ bl_0_472 br_0_472 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c472
+ bl_0_472 br_0_472 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c472
+ bl_0_472 br_0_472 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c472
+ bl_0_472 br_0_472 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c472
+ bl_0_472 br_0_472 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c472
+ bl_0_472 br_0_472 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c472
+ bl_0_472 br_0_472 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c472
+ bl_0_472 br_0_472 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c472
+ bl_0_472 br_0_472 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c472
+ bl_0_472 br_0_472 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c472
+ bl_0_472 br_0_472 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c472
+ bl_0_472 br_0_472 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c472
+ bl_0_472 br_0_472 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c472
+ bl_0_472 br_0_472 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c472
+ bl_0_472 br_0_472 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c472
+ bl_0_472 br_0_472 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c472
+ bl_0_472 br_0_472 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c472
+ bl_0_472 br_0_472 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c472
+ bl_0_472 br_0_472 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c473
+ bl_0_473 br_0_473 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c473
+ bl_0_473 br_0_473 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c473
+ bl_0_473 br_0_473 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c473
+ bl_0_473 br_0_473 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c473
+ bl_0_473 br_0_473 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c473
+ bl_0_473 br_0_473 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c473
+ bl_0_473 br_0_473 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c473
+ bl_0_473 br_0_473 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c473
+ bl_0_473 br_0_473 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c473
+ bl_0_473 br_0_473 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c473
+ bl_0_473 br_0_473 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c473
+ bl_0_473 br_0_473 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c473
+ bl_0_473 br_0_473 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c473
+ bl_0_473 br_0_473 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c473
+ bl_0_473 br_0_473 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c473
+ bl_0_473 br_0_473 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c473
+ bl_0_473 br_0_473 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c473
+ bl_0_473 br_0_473 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c473
+ bl_0_473 br_0_473 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c473
+ bl_0_473 br_0_473 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c473
+ bl_0_473 br_0_473 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c473
+ bl_0_473 br_0_473 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c473
+ bl_0_473 br_0_473 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c473
+ bl_0_473 br_0_473 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c473
+ bl_0_473 br_0_473 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c473
+ bl_0_473 br_0_473 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c473
+ bl_0_473 br_0_473 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c473
+ bl_0_473 br_0_473 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c473
+ bl_0_473 br_0_473 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c473
+ bl_0_473 br_0_473 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c473
+ bl_0_473 br_0_473 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c473
+ bl_0_473 br_0_473 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c473
+ bl_0_473 br_0_473 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c473
+ bl_0_473 br_0_473 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c473
+ bl_0_473 br_0_473 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c473
+ bl_0_473 br_0_473 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c473
+ bl_0_473 br_0_473 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c473
+ bl_0_473 br_0_473 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c473
+ bl_0_473 br_0_473 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c473
+ bl_0_473 br_0_473 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c473
+ bl_0_473 br_0_473 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c473
+ bl_0_473 br_0_473 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c473
+ bl_0_473 br_0_473 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c473
+ bl_0_473 br_0_473 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c473
+ bl_0_473 br_0_473 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c474
+ bl_0_474 br_0_474 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c474
+ bl_0_474 br_0_474 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c474
+ bl_0_474 br_0_474 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c474
+ bl_0_474 br_0_474 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c474
+ bl_0_474 br_0_474 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c474
+ bl_0_474 br_0_474 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c474
+ bl_0_474 br_0_474 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c474
+ bl_0_474 br_0_474 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c474
+ bl_0_474 br_0_474 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c474
+ bl_0_474 br_0_474 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c474
+ bl_0_474 br_0_474 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c474
+ bl_0_474 br_0_474 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c474
+ bl_0_474 br_0_474 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c474
+ bl_0_474 br_0_474 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c474
+ bl_0_474 br_0_474 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c474
+ bl_0_474 br_0_474 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c474
+ bl_0_474 br_0_474 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c474
+ bl_0_474 br_0_474 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c474
+ bl_0_474 br_0_474 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c474
+ bl_0_474 br_0_474 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c474
+ bl_0_474 br_0_474 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c474
+ bl_0_474 br_0_474 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c474
+ bl_0_474 br_0_474 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c474
+ bl_0_474 br_0_474 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c474
+ bl_0_474 br_0_474 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c474
+ bl_0_474 br_0_474 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c474
+ bl_0_474 br_0_474 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c474
+ bl_0_474 br_0_474 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c474
+ bl_0_474 br_0_474 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c474
+ bl_0_474 br_0_474 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c474
+ bl_0_474 br_0_474 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c474
+ bl_0_474 br_0_474 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c474
+ bl_0_474 br_0_474 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c474
+ bl_0_474 br_0_474 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c474
+ bl_0_474 br_0_474 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c474
+ bl_0_474 br_0_474 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c474
+ bl_0_474 br_0_474 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c474
+ bl_0_474 br_0_474 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c474
+ bl_0_474 br_0_474 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c474
+ bl_0_474 br_0_474 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c474
+ bl_0_474 br_0_474 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c474
+ bl_0_474 br_0_474 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c474
+ bl_0_474 br_0_474 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c474
+ bl_0_474 br_0_474 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c474
+ bl_0_474 br_0_474 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c475
+ bl_0_475 br_0_475 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c475
+ bl_0_475 br_0_475 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c475
+ bl_0_475 br_0_475 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c475
+ bl_0_475 br_0_475 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c475
+ bl_0_475 br_0_475 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c475
+ bl_0_475 br_0_475 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c475
+ bl_0_475 br_0_475 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c475
+ bl_0_475 br_0_475 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c475
+ bl_0_475 br_0_475 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c475
+ bl_0_475 br_0_475 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c475
+ bl_0_475 br_0_475 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c475
+ bl_0_475 br_0_475 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c475
+ bl_0_475 br_0_475 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c475
+ bl_0_475 br_0_475 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c475
+ bl_0_475 br_0_475 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c475
+ bl_0_475 br_0_475 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c475
+ bl_0_475 br_0_475 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c475
+ bl_0_475 br_0_475 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c475
+ bl_0_475 br_0_475 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c475
+ bl_0_475 br_0_475 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c475
+ bl_0_475 br_0_475 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c475
+ bl_0_475 br_0_475 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c475
+ bl_0_475 br_0_475 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c475
+ bl_0_475 br_0_475 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c475
+ bl_0_475 br_0_475 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c475
+ bl_0_475 br_0_475 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c475
+ bl_0_475 br_0_475 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c475
+ bl_0_475 br_0_475 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c475
+ bl_0_475 br_0_475 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c475
+ bl_0_475 br_0_475 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c475
+ bl_0_475 br_0_475 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c475
+ bl_0_475 br_0_475 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c475
+ bl_0_475 br_0_475 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c475
+ bl_0_475 br_0_475 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c475
+ bl_0_475 br_0_475 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c475
+ bl_0_475 br_0_475 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c475
+ bl_0_475 br_0_475 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c475
+ bl_0_475 br_0_475 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c475
+ bl_0_475 br_0_475 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c475
+ bl_0_475 br_0_475 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c475
+ bl_0_475 br_0_475 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c475
+ bl_0_475 br_0_475 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c475
+ bl_0_475 br_0_475 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c475
+ bl_0_475 br_0_475 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c475
+ bl_0_475 br_0_475 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c476
+ bl_0_476 br_0_476 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c476
+ bl_0_476 br_0_476 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c476
+ bl_0_476 br_0_476 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c476
+ bl_0_476 br_0_476 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c476
+ bl_0_476 br_0_476 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c476
+ bl_0_476 br_0_476 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c476
+ bl_0_476 br_0_476 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c476
+ bl_0_476 br_0_476 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c476
+ bl_0_476 br_0_476 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c476
+ bl_0_476 br_0_476 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c476
+ bl_0_476 br_0_476 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c476
+ bl_0_476 br_0_476 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c476
+ bl_0_476 br_0_476 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c476
+ bl_0_476 br_0_476 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c476
+ bl_0_476 br_0_476 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c476
+ bl_0_476 br_0_476 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c476
+ bl_0_476 br_0_476 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c476
+ bl_0_476 br_0_476 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c476
+ bl_0_476 br_0_476 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c476
+ bl_0_476 br_0_476 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c476
+ bl_0_476 br_0_476 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c476
+ bl_0_476 br_0_476 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c476
+ bl_0_476 br_0_476 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c476
+ bl_0_476 br_0_476 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c476
+ bl_0_476 br_0_476 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c476
+ bl_0_476 br_0_476 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c476
+ bl_0_476 br_0_476 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c476
+ bl_0_476 br_0_476 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c476
+ bl_0_476 br_0_476 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c476
+ bl_0_476 br_0_476 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c476
+ bl_0_476 br_0_476 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c476
+ bl_0_476 br_0_476 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c476
+ bl_0_476 br_0_476 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c476
+ bl_0_476 br_0_476 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c476
+ bl_0_476 br_0_476 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c476
+ bl_0_476 br_0_476 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c476
+ bl_0_476 br_0_476 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c476
+ bl_0_476 br_0_476 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c476
+ bl_0_476 br_0_476 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c476
+ bl_0_476 br_0_476 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c476
+ bl_0_476 br_0_476 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c476
+ bl_0_476 br_0_476 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c476
+ bl_0_476 br_0_476 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c476
+ bl_0_476 br_0_476 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c476
+ bl_0_476 br_0_476 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c477
+ bl_0_477 br_0_477 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c477
+ bl_0_477 br_0_477 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c477
+ bl_0_477 br_0_477 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c477
+ bl_0_477 br_0_477 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c477
+ bl_0_477 br_0_477 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c477
+ bl_0_477 br_0_477 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c477
+ bl_0_477 br_0_477 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c477
+ bl_0_477 br_0_477 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c477
+ bl_0_477 br_0_477 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c477
+ bl_0_477 br_0_477 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c477
+ bl_0_477 br_0_477 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c477
+ bl_0_477 br_0_477 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c477
+ bl_0_477 br_0_477 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c477
+ bl_0_477 br_0_477 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c477
+ bl_0_477 br_0_477 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c477
+ bl_0_477 br_0_477 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c477
+ bl_0_477 br_0_477 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c477
+ bl_0_477 br_0_477 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c477
+ bl_0_477 br_0_477 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c477
+ bl_0_477 br_0_477 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c477
+ bl_0_477 br_0_477 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c477
+ bl_0_477 br_0_477 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c477
+ bl_0_477 br_0_477 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c477
+ bl_0_477 br_0_477 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c477
+ bl_0_477 br_0_477 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c477
+ bl_0_477 br_0_477 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c477
+ bl_0_477 br_0_477 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c477
+ bl_0_477 br_0_477 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c477
+ bl_0_477 br_0_477 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c477
+ bl_0_477 br_0_477 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c477
+ bl_0_477 br_0_477 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c477
+ bl_0_477 br_0_477 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c477
+ bl_0_477 br_0_477 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c477
+ bl_0_477 br_0_477 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c477
+ bl_0_477 br_0_477 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c477
+ bl_0_477 br_0_477 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c477
+ bl_0_477 br_0_477 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c477
+ bl_0_477 br_0_477 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c477
+ bl_0_477 br_0_477 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c477
+ bl_0_477 br_0_477 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c477
+ bl_0_477 br_0_477 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c477
+ bl_0_477 br_0_477 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c477
+ bl_0_477 br_0_477 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c477
+ bl_0_477 br_0_477 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c477
+ bl_0_477 br_0_477 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c478
+ bl_0_478 br_0_478 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c478
+ bl_0_478 br_0_478 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c478
+ bl_0_478 br_0_478 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c478
+ bl_0_478 br_0_478 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c478
+ bl_0_478 br_0_478 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c478
+ bl_0_478 br_0_478 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c478
+ bl_0_478 br_0_478 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c478
+ bl_0_478 br_0_478 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c478
+ bl_0_478 br_0_478 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c478
+ bl_0_478 br_0_478 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c478
+ bl_0_478 br_0_478 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c478
+ bl_0_478 br_0_478 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c478
+ bl_0_478 br_0_478 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c478
+ bl_0_478 br_0_478 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c478
+ bl_0_478 br_0_478 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c478
+ bl_0_478 br_0_478 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c478
+ bl_0_478 br_0_478 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c478
+ bl_0_478 br_0_478 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c478
+ bl_0_478 br_0_478 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c478
+ bl_0_478 br_0_478 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c478
+ bl_0_478 br_0_478 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c478
+ bl_0_478 br_0_478 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c478
+ bl_0_478 br_0_478 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c478
+ bl_0_478 br_0_478 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c478
+ bl_0_478 br_0_478 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c478
+ bl_0_478 br_0_478 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c478
+ bl_0_478 br_0_478 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c478
+ bl_0_478 br_0_478 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c478
+ bl_0_478 br_0_478 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c478
+ bl_0_478 br_0_478 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c478
+ bl_0_478 br_0_478 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c478
+ bl_0_478 br_0_478 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c478
+ bl_0_478 br_0_478 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c478
+ bl_0_478 br_0_478 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c478
+ bl_0_478 br_0_478 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c478
+ bl_0_478 br_0_478 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c478
+ bl_0_478 br_0_478 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c478
+ bl_0_478 br_0_478 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c478
+ bl_0_478 br_0_478 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c478
+ bl_0_478 br_0_478 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c478
+ bl_0_478 br_0_478 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c478
+ bl_0_478 br_0_478 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c478
+ bl_0_478 br_0_478 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c478
+ bl_0_478 br_0_478 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c478
+ bl_0_478 br_0_478 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c479
+ bl_0_479 br_0_479 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c479
+ bl_0_479 br_0_479 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c479
+ bl_0_479 br_0_479 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c479
+ bl_0_479 br_0_479 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c479
+ bl_0_479 br_0_479 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c479
+ bl_0_479 br_0_479 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c479
+ bl_0_479 br_0_479 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c479
+ bl_0_479 br_0_479 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c479
+ bl_0_479 br_0_479 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c479
+ bl_0_479 br_0_479 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c479
+ bl_0_479 br_0_479 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c479
+ bl_0_479 br_0_479 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c479
+ bl_0_479 br_0_479 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c479
+ bl_0_479 br_0_479 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c479
+ bl_0_479 br_0_479 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c479
+ bl_0_479 br_0_479 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c479
+ bl_0_479 br_0_479 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c479
+ bl_0_479 br_0_479 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c479
+ bl_0_479 br_0_479 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c479
+ bl_0_479 br_0_479 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c479
+ bl_0_479 br_0_479 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c479
+ bl_0_479 br_0_479 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c479
+ bl_0_479 br_0_479 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c479
+ bl_0_479 br_0_479 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c479
+ bl_0_479 br_0_479 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c479
+ bl_0_479 br_0_479 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c479
+ bl_0_479 br_0_479 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c479
+ bl_0_479 br_0_479 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c479
+ bl_0_479 br_0_479 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c479
+ bl_0_479 br_0_479 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c479
+ bl_0_479 br_0_479 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c479
+ bl_0_479 br_0_479 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c479
+ bl_0_479 br_0_479 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c479
+ bl_0_479 br_0_479 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c479
+ bl_0_479 br_0_479 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c479
+ bl_0_479 br_0_479 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c479
+ bl_0_479 br_0_479 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c479
+ bl_0_479 br_0_479 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c479
+ bl_0_479 br_0_479 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c479
+ bl_0_479 br_0_479 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c479
+ bl_0_479 br_0_479 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c479
+ bl_0_479 br_0_479 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c479
+ bl_0_479 br_0_479 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c479
+ bl_0_479 br_0_479 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c479
+ bl_0_479 br_0_479 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c480
+ bl_0_480 br_0_480 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c480
+ bl_0_480 br_0_480 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c480
+ bl_0_480 br_0_480 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c480
+ bl_0_480 br_0_480 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c480
+ bl_0_480 br_0_480 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c480
+ bl_0_480 br_0_480 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c480
+ bl_0_480 br_0_480 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c480
+ bl_0_480 br_0_480 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c480
+ bl_0_480 br_0_480 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c480
+ bl_0_480 br_0_480 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c480
+ bl_0_480 br_0_480 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c480
+ bl_0_480 br_0_480 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c480
+ bl_0_480 br_0_480 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c480
+ bl_0_480 br_0_480 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c480
+ bl_0_480 br_0_480 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c480
+ bl_0_480 br_0_480 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c480
+ bl_0_480 br_0_480 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c480
+ bl_0_480 br_0_480 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c480
+ bl_0_480 br_0_480 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c480
+ bl_0_480 br_0_480 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c480
+ bl_0_480 br_0_480 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c480
+ bl_0_480 br_0_480 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c480
+ bl_0_480 br_0_480 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c480
+ bl_0_480 br_0_480 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c480
+ bl_0_480 br_0_480 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c480
+ bl_0_480 br_0_480 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c480
+ bl_0_480 br_0_480 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c480
+ bl_0_480 br_0_480 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c480
+ bl_0_480 br_0_480 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c480
+ bl_0_480 br_0_480 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c480
+ bl_0_480 br_0_480 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c480
+ bl_0_480 br_0_480 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c480
+ bl_0_480 br_0_480 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c480
+ bl_0_480 br_0_480 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c480
+ bl_0_480 br_0_480 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c480
+ bl_0_480 br_0_480 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c480
+ bl_0_480 br_0_480 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c480
+ bl_0_480 br_0_480 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c480
+ bl_0_480 br_0_480 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c480
+ bl_0_480 br_0_480 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c480
+ bl_0_480 br_0_480 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c480
+ bl_0_480 br_0_480 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c480
+ bl_0_480 br_0_480 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c480
+ bl_0_480 br_0_480 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c480
+ bl_0_480 br_0_480 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c481
+ bl_0_481 br_0_481 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c481
+ bl_0_481 br_0_481 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c481
+ bl_0_481 br_0_481 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c481
+ bl_0_481 br_0_481 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c481
+ bl_0_481 br_0_481 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c481
+ bl_0_481 br_0_481 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c481
+ bl_0_481 br_0_481 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c481
+ bl_0_481 br_0_481 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c481
+ bl_0_481 br_0_481 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c481
+ bl_0_481 br_0_481 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c481
+ bl_0_481 br_0_481 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c481
+ bl_0_481 br_0_481 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c481
+ bl_0_481 br_0_481 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c481
+ bl_0_481 br_0_481 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c481
+ bl_0_481 br_0_481 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c481
+ bl_0_481 br_0_481 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c481
+ bl_0_481 br_0_481 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c481
+ bl_0_481 br_0_481 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c481
+ bl_0_481 br_0_481 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c481
+ bl_0_481 br_0_481 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c481
+ bl_0_481 br_0_481 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c481
+ bl_0_481 br_0_481 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c481
+ bl_0_481 br_0_481 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c481
+ bl_0_481 br_0_481 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c481
+ bl_0_481 br_0_481 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c481
+ bl_0_481 br_0_481 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c481
+ bl_0_481 br_0_481 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c481
+ bl_0_481 br_0_481 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c481
+ bl_0_481 br_0_481 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c481
+ bl_0_481 br_0_481 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c481
+ bl_0_481 br_0_481 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c481
+ bl_0_481 br_0_481 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c481
+ bl_0_481 br_0_481 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c481
+ bl_0_481 br_0_481 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c481
+ bl_0_481 br_0_481 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c481
+ bl_0_481 br_0_481 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c481
+ bl_0_481 br_0_481 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c481
+ bl_0_481 br_0_481 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c481
+ bl_0_481 br_0_481 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c481
+ bl_0_481 br_0_481 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c481
+ bl_0_481 br_0_481 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c481
+ bl_0_481 br_0_481 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c481
+ bl_0_481 br_0_481 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c481
+ bl_0_481 br_0_481 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c481
+ bl_0_481 br_0_481 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c482
+ bl_0_482 br_0_482 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c482
+ bl_0_482 br_0_482 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c482
+ bl_0_482 br_0_482 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c482
+ bl_0_482 br_0_482 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c482
+ bl_0_482 br_0_482 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c482
+ bl_0_482 br_0_482 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c482
+ bl_0_482 br_0_482 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c482
+ bl_0_482 br_0_482 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c482
+ bl_0_482 br_0_482 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c482
+ bl_0_482 br_0_482 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c482
+ bl_0_482 br_0_482 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c482
+ bl_0_482 br_0_482 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c482
+ bl_0_482 br_0_482 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c482
+ bl_0_482 br_0_482 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c482
+ bl_0_482 br_0_482 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c482
+ bl_0_482 br_0_482 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c482
+ bl_0_482 br_0_482 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c482
+ bl_0_482 br_0_482 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c482
+ bl_0_482 br_0_482 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c482
+ bl_0_482 br_0_482 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c482
+ bl_0_482 br_0_482 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c482
+ bl_0_482 br_0_482 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c482
+ bl_0_482 br_0_482 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c482
+ bl_0_482 br_0_482 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c482
+ bl_0_482 br_0_482 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c482
+ bl_0_482 br_0_482 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c482
+ bl_0_482 br_0_482 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c482
+ bl_0_482 br_0_482 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c482
+ bl_0_482 br_0_482 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c482
+ bl_0_482 br_0_482 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c482
+ bl_0_482 br_0_482 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c482
+ bl_0_482 br_0_482 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c482
+ bl_0_482 br_0_482 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c482
+ bl_0_482 br_0_482 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c482
+ bl_0_482 br_0_482 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c482
+ bl_0_482 br_0_482 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c482
+ bl_0_482 br_0_482 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c482
+ bl_0_482 br_0_482 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c482
+ bl_0_482 br_0_482 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c482
+ bl_0_482 br_0_482 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c482
+ bl_0_482 br_0_482 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c482
+ bl_0_482 br_0_482 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c482
+ bl_0_482 br_0_482 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c482
+ bl_0_482 br_0_482 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c482
+ bl_0_482 br_0_482 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c483
+ bl_0_483 br_0_483 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c483
+ bl_0_483 br_0_483 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c483
+ bl_0_483 br_0_483 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c483
+ bl_0_483 br_0_483 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c483
+ bl_0_483 br_0_483 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c483
+ bl_0_483 br_0_483 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c483
+ bl_0_483 br_0_483 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c483
+ bl_0_483 br_0_483 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c483
+ bl_0_483 br_0_483 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c483
+ bl_0_483 br_0_483 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c483
+ bl_0_483 br_0_483 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c483
+ bl_0_483 br_0_483 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c483
+ bl_0_483 br_0_483 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c483
+ bl_0_483 br_0_483 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c483
+ bl_0_483 br_0_483 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c483
+ bl_0_483 br_0_483 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c483
+ bl_0_483 br_0_483 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c483
+ bl_0_483 br_0_483 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c483
+ bl_0_483 br_0_483 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c483
+ bl_0_483 br_0_483 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c483
+ bl_0_483 br_0_483 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c483
+ bl_0_483 br_0_483 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c483
+ bl_0_483 br_0_483 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c483
+ bl_0_483 br_0_483 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c483
+ bl_0_483 br_0_483 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c483
+ bl_0_483 br_0_483 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c483
+ bl_0_483 br_0_483 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c483
+ bl_0_483 br_0_483 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c483
+ bl_0_483 br_0_483 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c483
+ bl_0_483 br_0_483 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c483
+ bl_0_483 br_0_483 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c483
+ bl_0_483 br_0_483 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c483
+ bl_0_483 br_0_483 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c483
+ bl_0_483 br_0_483 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c483
+ bl_0_483 br_0_483 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c483
+ bl_0_483 br_0_483 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c483
+ bl_0_483 br_0_483 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c483
+ bl_0_483 br_0_483 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c483
+ bl_0_483 br_0_483 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c483
+ bl_0_483 br_0_483 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c483
+ bl_0_483 br_0_483 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c483
+ bl_0_483 br_0_483 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c483
+ bl_0_483 br_0_483 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c483
+ bl_0_483 br_0_483 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c483
+ bl_0_483 br_0_483 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c484
+ bl_0_484 br_0_484 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c484
+ bl_0_484 br_0_484 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c484
+ bl_0_484 br_0_484 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c484
+ bl_0_484 br_0_484 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c484
+ bl_0_484 br_0_484 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c484
+ bl_0_484 br_0_484 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c484
+ bl_0_484 br_0_484 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c484
+ bl_0_484 br_0_484 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c484
+ bl_0_484 br_0_484 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c484
+ bl_0_484 br_0_484 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c484
+ bl_0_484 br_0_484 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c484
+ bl_0_484 br_0_484 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c484
+ bl_0_484 br_0_484 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c484
+ bl_0_484 br_0_484 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c484
+ bl_0_484 br_0_484 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c484
+ bl_0_484 br_0_484 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c484
+ bl_0_484 br_0_484 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c484
+ bl_0_484 br_0_484 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c484
+ bl_0_484 br_0_484 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c484
+ bl_0_484 br_0_484 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c484
+ bl_0_484 br_0_484 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c484
+ bl_0_484 br_0_484 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c484
+ bl_0_484 br_0_484 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c484
+ bl_0_484 br_0_484 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c484
+ bl_0_484 br_0_484 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c484
+ bl_0_484 br_0_484 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c484
+ bl_0_484 br_0_484 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c484
+ bl_0_484 br_0_484 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c484
+ bl_0_484 br_0_484 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c484
+ bl_0_484 br_0_484 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c484
+ bl_0_484 br_0_484 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c484
+ bl_0_484 br_0_484 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c484
+ bl_0_484 br_0_484 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c484
+ bl_0_484 br_0_484 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c484
+ bl_0_484 br_0_484 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c484
+ bl_0_484 br_0_484 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c484
+ bl_0_484 br_0_484 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c484
+ bl_0_484 br_0_484 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c484
+ bl_0_484 br_0_484 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c484
+ bl_0_484 br_0_484 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c484
+ bl_0_484 br_0_484 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c484
+ bl_0_484 br_0_484 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c484
+ bl_0_484 br_0_484 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c484
+ bl_0_484 br_0_484 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c484
+ bl_0_484 br_0_484 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c485
+ bl_0_485 br_0_485 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c485
+ bl_0_485 br_0_485 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c485
+ bl_0_485 br_0_485 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c485
+ bl_0_485 br_0_485 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c485
+ bl_0_485 br_0_485 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c485
+ bl_0_485 br_0_485 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c485
+ bl_0_485 br_0_485 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c485
+ bl_0_485 br_0_485 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c485
+ bl_0_485 br_0_485 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c485
+ bl_0_485 br_0_485 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c485
+ bl_0_485 br_0_485 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c485
+ bl_0_485 br_0_485 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c485
+ bl_0_485 br_0_485 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c485
+ bl_0_485 br_0_485 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c485
+ bl_0_485 br_0_485 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c485
+ bl_0_485 br_0_485 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c485
+ bl_0_485 br_0_485 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c485
+ bl_0_485 br_0_485 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c485
+ bl_0_485 br_0_485 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c485
+ bl_0_485 br_0_485 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c485
+ bl_0_485 br_0_485 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c485
+ bl_0_485 br_0_485 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c485
+ bl_0_485 br_0_485 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c485
+ bl_0_485 br_0_485 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c485
+ bl_0_485 br_0_485 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c485
+ bl_0_485 br_0_485 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c485
+ bl_0_485 br_0_485 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c485
+ bl_0_485 br_0_485 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c485
+ bl_0_485 br_0_485 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c485
+ bl_0_485 br_0_485 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c485
+ bl_0_485 br_0_485 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c485
+ bl_0_485 br_0_485 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c485
+ bl_0_485 br_0_485 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c485
+ bl_0_485 br_0_485 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c485
+ bl_0_485 br_0_485 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c485
+ bl_0_485 br_0_485 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c485
+ bl_0_485 br_0_485 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c485
+ bl_0_485 br_0_485 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c485
+ bl_0_485 br_0_485 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c485
+ bl_0_485 br_0_485 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c485
+ bl_0_485 br_0_485 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c485
+ bl_0_485 br_0_485 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c485
+ bl_0_485 br_0_485 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c485
+ bl_0_485 br_0_485 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c485
+ bl_0_485 br_0_485 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c486
+ bl_0_486 br_0_486 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c486
+ bl_0_486 br_0_486 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c486
+ bl_0_486 br_0_486 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c486
+ bl_0_486 br_0_486 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c486
+ bl_0_486 br_0_486 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c486
+ bl_0_486 br_0_486 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c486
+ bl_0_486 br_0_486 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c486
+ bl_0_486 br_0_486 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c486
+ bl_0_486 br_0_486 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c486
+ bl_0_486 br_0_486 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c486
+ bl_0_486 br_0_486 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c486
+ bl_0_486 br_0_486 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c486
+ bl_0_486 br_0_486 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c486
+ bl_0_486 br_0_486 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c486
+ bl_0_486 br_0_486 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c486
+ bl_0_486 br_0_486 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c486
+ bl_0_486 br_0_486 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c486
+ bl_0_486 br_0_486 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c486
+ bl_0_486 br_0_486 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c486
+ bl_0_486 br_0_486 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c486
+ bl_0_486 br_0_486 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c486
+ bl_0_486 br_0_486 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c486
+ bl_0_486 br_0_486 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c486
+ bl_0_486 br_0_486 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c486
+ bl_0_486 br_0_486 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c486
+ bl_0_486 br_0_486 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c486
+ bl_0_486 br_0_486 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c486
+ bl_0_486 br_0_486 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c486
+ bl_0_486 br_0_486 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c486
+ bl_0_486 br_0_486 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c486
+ bl_0_486 br_0_486 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c486
+ bl_0_486 br_0_486 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c486
+ bl_0_486 br_0_486 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c486
+ bl_0_486 br_0_486 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c486
+ bl_0_486 br_0_486 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c486
+ bl_0_486 br_0_486 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c486
+ bl_0_486 br_0_486 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c486
+ bl_0_486 br_0_486 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c486
+ bl_0_486 br_0_486 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c486
+ bl_0_486 br_0_486 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c486
+ bl_0_486 br_0_486 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c486
+ bl_0_486 br_0_486 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c486
+ bl_0_486 br_0_486 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c486
+ bl_0_486 br_0_486 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c486
+ bl_0_486 br_0_486 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c487
+ bl_0_487 br_0_487 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c487
+ bl_0_487 br_0_487 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c487
+ bl_0_487 br_0_487 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c487
+ bl_0_487 br_0_487 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c487
+ bl_0_487 br_0_487 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c487
+ bl_0_487 br_0_487 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c487
+ bl_0_487 br_0_487 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c487
+ bl_0_487 br_0_487 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c487
+ bl_0_487 br_0_487 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c487
+ bl_0_487 br_0_487 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c487
+ bl_0_487 br_0_487 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c487
+ bl_0_487 br_0_487 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c487
+ bl_0_487 br_0_487 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c487
+ bl_0_487 br_0_487 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c487
+ bl_0_487 br_0_487 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c487
+ bl_0_487 br_0_487 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c487
+ bl_0_487 br_0_487 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c487
+ bl_0_487 br_0_487 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c487
+ bl_0_487 br_0_487 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c487
+ bl_0_487 br_0_487 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c487
+ bl_0_487 br_0_487 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c487
+ bl_0_487 br_0_487 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c487
+ bl_0_487 br_0_487 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c487
+ bl_0_487 br_0_487 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c487
+ bl_0_487 br_0_487 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c487
+ bl_0_487 br_0_487 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c487
+ bl_0_487 br_0_487 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c487
+ bl_0_487 br_0_487 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c487
+ bl_0_487 br_0_487 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c487
+ bl_0_487 br_0_487 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c487
+ bl_0_487 br_0_487 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c487
+ bl_0_487 br_0_487 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c487
+ bl_0_487 br_0_487 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c487
+ bl_0_487 br_0_487 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c487
+ bl_0_487 br_0_487 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c487
+ bl_0_487 br_0_487 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c487
+ bl_0_487 br_0_487 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c487
+ bl_0_487 br_0_487 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c487
+ bl_0_487 br_0_487 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c487
+ bl_0_487 br_0_487 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c487
+ bl_0_487 br_0_487 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c487
+ bl_0_487 br_0_487 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c487
+ bl_0_487 br_0_487 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c487
+ bl_0_487 br_0_487 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c487
+ bl_0_487 br_0_487 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c488
+ bl_0_488 br_0_488 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c488
+ bl_0_488 br_0_488 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c488
+ bl_0_488 br_0_488 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c488
+ bl_0_488 br_0_488 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c488
+ bl_0_488 br_0_488 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c488
+ bl_0_488 br_0_488 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c488
+ bl_0_488 br_0_488 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c488
+ bl_0_488 br_0_488 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c488
+ bl_0_488 br_0_488 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c488
+ bl_0_488 br_0_488 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c488
+ bl_0_488 br_0_488 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c488
+ bl_0_488 br_0_488 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c488
+ bl_0_488 br_0_488 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c488
+ bl_0_488 br_0_488 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c488
+ bl_0_488 br_0_488 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c488
+ bl_0_488 br_0_488 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c488
+ bl_0_488 br_0_488 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c488
+ bl_0_488 br_0_488 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c488
+ bl_0_488 br_0_488 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c488
+ bl_0_488 br_0_488 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c488
+ bl_0_488 br_0_488 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c488
+ bl_0_488 br_0_488 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c488
+ bl_0_488 br_0_488 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c488
+ bl_0_488 br_0_488 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c488
+ bl_0_488 br_0_488 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c488
+ bl_0_488 br_0_488 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c488
+ bl_0_488 br_0_488 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c488
+ bl_0_488 br_0_488 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c488
+ bl_0_488 br_0_488 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c488
+ bl_0_488 br_0_488 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c488
+ bl_0_488 br_0_488 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c488
+ bl_0_488 br_0_488 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c488
+ bl_0_488 br_0_488 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c488
+ bl_0_488 br_0_488 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c488
+ bl_0_488 br_0_488 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c488
+ bl_0_488 br_0_488 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c488
+ bl_0_488 br_0_488 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c488
+ bl_0_488 br_0_488 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c488
+ bl_0_488 br_0_488 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c488
+ bl_0_488 br_0_488 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c488
+ bl_0_488 br_0_488 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c488
+ bl_0_488 br_0_488 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c488
+ bl_0_488 br_0_488 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c488
+ bl_0_488 br_0_488 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c488
+ bl_0_488 br_0_488 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c489
+ bl_0_489 br_0_489 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c489
+ bl_0_489 br_0_489 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c489
+ bl_0_489 br_0_489 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c489
+ bl_0_489 br_0_489 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c489
+ bl_0_489 br_0_489 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c489
+ bl_0_489 br_0_489 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c489
+ bl_0_489 br_0_489 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c489
+ bl_0_489 br_0_489 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c489
+ bl_0_489 br_0_489 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c489
+ bl_0_489 br_0_489 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c489
+ bl_0_489 br_0_489 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c489
+ bl_0_489 br_0_489 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c489
+ bl_0_489 br_0_489 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c489
+ bl_0_489 br_0_489 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c489
+ bl_0_489 br_0_489 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c489
+ bl_0_489 br_0_489 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c489
+ bl_0_489 br_0_489 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c489
+ bl_0_489 br_0_489 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c489
+ bl_0_489 br_0_489 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c489
+ bl_0_489 br_0_489 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c489
+ bl_0_489 br_0_489 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c489
+ bl_0_489 br_0_489 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c489
+ bl_0_489 br_0_489 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c489
+ bl_0_489 br_0_489 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c489
+ bl_0_489 br_0_489 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c489
+ bl_0_489 br_0_489 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c489
+ bl_0_489 br_0_489 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c489
+ bl_0_489 br_0_489 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c489
+ bl_0_489 br_0_489 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c489
+ bl_0_489 br_0_489 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c489
+ bl_0_489 br_0_489 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c489
+ bl_0_489 br_0_489 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c489
+ bl_0_489 br_0_489 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c489
+ bl_0_489 br_0_489 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c489
+ bl_0_489 br_0_489 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c489
+ bl_0_489 br_0_489 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c489
+ bl_0_489 br_0_489 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c489
+ bl_0_489 br_0_489 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c489
+ bl_0_489 br_0_489 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c489
+ bl_0_489 br_0_489 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c489
+ bl_0_489 br_0_489 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c489
+ bl_0_489 br_0_489 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c489
+ bl_0_489 br_0_489 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c489
+ bl_0_489 br_0_489 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c489
+ bl_0_489 br_0_489 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c490
+ bl_0_490 br_0_490 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c490
+ bl_0_490 br_0_490 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c490
+ bl_0_490 br_0_490 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c490
+ bl_0_490 br_0_490 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c490
+ bl_0_490 br_0_490 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c490
+ bl_0_490 br_0_490 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c490
+ bl_0_490 br_0_490 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c490
+ bl_0_490 br_0_490 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c490
+ bl_0_490 br_0_490 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c490
+ bl_0_490 br_0_490 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c490
+ bl_0_490 br_0_490 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c490
+ bl_0_490 br_0_490 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c490
+ bl_0_490 br_0_490 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c490
+ bl_0_490 br_0_490 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c490
+ bl_0_490 br_0_490 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c490
+ bl_0_490 br_0_490 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c490
+ bl_0_490 br_0_490 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c490
+ bl_0_490 br_0_490 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c490
+ bl_0_490 br_0_490 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c490
+ bl_0_490 br_0_490 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c490
+ bl_0_490 br_0_490 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c490
+ bl_0_490 br_0_490 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c490
+ bl_0_490 br_0_490 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c490
+ bl_0_490 br_0_490 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c490
+ bl_0_490 br_0_490 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c490
+ bl_0_490 br_0_490 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c490
+ bl_0_490 br_0_490 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c490
+ bl_0_490 br_0_490 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c490
+ bl_0_490 br_0_490 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c490
+ bl_0_490 br_0_490 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c490
+ bl_0_490 br_0_490 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c490
+ bl_0_490 br_0_490 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c490
+ bl_0_490 br_0_490 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c490
+ bl_0_490 br_0_490 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c490
+ bl_0_490 br_0_490 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c490
+ bl_0_490 br_0_490 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c490
+ bl_0_490 br_0_490 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c490
+ bl_0_490 br_0_490 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c490
+ bl_0_490 br_0_490 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c490
+ bl_0_490 br_0_490 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c490
+ bl_0_490 br_0_490 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c490
+ bl_0_490 br_0_490 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c490
+ bl_0_490 br_0_490 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c490
+ bl_0_490 br_0_490 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c490
+ bl_0_490 br_0_490 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c491
+ bl_0_491 br_0_491 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c491
+ bl_0_491 br_0_491 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c491
+ bl_0_491 br_0_491 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c491
+ bl_0_491 br_0_491 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c491
+ bl_0_491 br_0_491 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c491
+ bl_0_491 br_0_491 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c491
+ bl_0_491 br_0_491 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c491
+ bl_0_491 br_0_491 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c491
+ bl_0_491 br_0_491 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c491
+ bl_0_491 br_0_491 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c491
+ bl_0_491 br_0_491 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c491
+ bl_0_491 br_0_491 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c491
+ bl_0_491 br_0_491 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c491
+ bl_0_491 br_0_491 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c491
+ bl_0_491 br_0_491 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c491
+ bl_0_491 br_0_491 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c491
+ bl_0_491 br_0_491 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c491
+ bl_0_491 br_0_491 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c491
+ bl_0_491 br_0_491 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c491
+ bl_0_491 br_0_491 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c491
+ bl_0_491 br_0_491 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c491
+ bl_0_491 br_0_491 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c491
+ bl_0_491 br_0_491 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c491
+ bl_0_491 br_0_491 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c491
+ bl_0_491 br_0_491 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c491
+ bl_0_491 br_0_491 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c491
+ bl_0_491 br_0_491 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c491
+ bl_0_491 br_0_491 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c491
+ bl_0_491 br_0_491 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c491
+ bl_0_491 br_0_491 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c491
+ bl_0_491 br_0_491 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c491
+ bl_0_491 br_0_491 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c491
+ bl_0_491 br_0_491 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c491
+ bl_0_491 br_0_491 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c491
+ bl_0_491 br_0_491 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c491
+ bl_0_491 br_0_491 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c491
+ bl_0_491 br_0_491 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c491
+ bl_0_491 br_0_491 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c491
+ bl_0_491 br_0_491 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c491
+ bl_0_491 br_0_491 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c491
+ bl_0_491 br_0_491 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c491
+ bl_0_491 br_0_491 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c491
+ bl_0_491 br_0_491 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c491
+ bl_0_491 br_0_491 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c491
+ bl_0_491 br_0_491 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c492
+ bl_0_492 br_0_492 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c492
+ bl_0_492 br_0_492 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c492
+ bl_0_492 br_0_492 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c492
+ bl_0_492 br_0_492 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c492
+ bl_0_492 br_0_492 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c492
+ bl_0_492 br_0_492 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c492
+ bl_0_492 br_0_492 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c492
+ bl_0_492 br_0_492 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c492
+ bl_0_492 br_0_492 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c492
+ bl_0_492 br_0_492 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c492
+ bl_0_492 br_0_492 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c492
+ bl_0_492 br_0_492 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c492
+ bl_0_492 br_0_492 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c492
+ bl_0_492 br_0_492 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c492
+ bl_0_492 br_0_492 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c492
+ bl_0_492 br_0_492 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c492
+ bl_0_492 br_0_492 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c492
+ bl_0_492 br_0_492 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c492
+ bl_0_492 br_0_492 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c492
+ bl_0_492 br_0_492 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c492
+ bl_0_492 br_0_492 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c492
+ bl_0_492 br_0_492 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c492
+ bl_0_492 br_0_492 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c492
+ bl_0_492 br_0_492 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c492
+ bl_0_492 br_0_492 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c492
+ bl_0_492 br_0_492 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c492
+ bl_0_492 br_0_492 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c492
+ bl_0_492 br_0_492 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c492
+ bl_0_492 br_0_492 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c492
+ bl_0_492 br_0_492 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c492
+ bl_0_492 br_0_492 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c492
+ bl_0_492 br_0_492 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c492
+ bl_0_492 br_0_492 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c492
+ bl_0_492 br_0_492 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c492
+ bl_0_492 br_0_492 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c492
+ bl_0_492 br_0_492 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c492
+ bl_0_492 br_0_492 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c492
+ bl_0_492 br_0_492 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c492
+ bl_0_492 br_0_492 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c492
+ bl_0_492 br_0_492 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c492
+ bl_0_492 br_0_492 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c492
+ bl_0_492 br_0_492 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c492
+ bl_0_492 br_0_492 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c492
+ bl_0_492 br_0_492 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c492
+ bl_0_492 br_0_492 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c493
+ bl_0_493 br_0_493 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c493
+ bl_0_493 br_0_493 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c493
+ bl_0_493 br_0_493 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c493
+ bl_0_493 br_0_493 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c493
+ bl_0_493 br_0_493 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c493
+ bl_0_493 br_0_493 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c493
+ bl_0_493 br_0_493 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c493
+ bl_0_493 br_0_493 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c493
+ bl_0_493 br_0_493 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c493
+ bl_0_493 br_0_493 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c493
+ bl_0_493 br_0_493 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c493
+ bl_0_493 br_0_493 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c493
+ bl_0_493 br_0_493 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c493
+ bl_0_493 br_0_493 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c493
+ bl_0_493 br_0_493 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c493
+ bl_0_493 br_0_493 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c493
+ bl_0_493 br_0_493 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c493
+ bl_0_493 br_0_493 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c493
+ bl_0_493 br_0_493 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c493
+ bl_0_493 br_0_493 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c493
+ bl_0_493 br_0_493 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c493
+ bl_0_493 br_0_493 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c493
+ bl_0_493 br_0_493 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c493
+ bl_0_493 br_0_493 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c493
+ bl_0_493 br_0_493 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c493
+ bl_0_493 br_0_493 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c493
+ bl_0_493 br_0_493 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c493
+ bl_0_493 br_0_493 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c493
+ bl_0_493 br_0_493 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c493
+ bl_0_493 br_0_493 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c493
+ bl_0_493 br_0_493 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c493
+ bl_0_493 br_0_493 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c493
+ bl_0_493 br_0_493 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c493
+ bl_0_493 br_0_493 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c493
+ bl_0_493 br_0_493 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c493
+ bl_0_493 br_0_493 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c493
+ bl_0_493 br_0_493 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c493
+ bl_0_493 br_0_493 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c493
+ bl_0_493 br_0_493 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c493
+ bl_0_493 br_0_493 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c493
+ bl_0_493 br_0_493 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c493
+ bl_0_493 br_0_493 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c493
+ bl_0_493 br_0_493 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c493
+ bl_0_493 br_0_493 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c493
+ bl_0_493 br_0_493 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c494
+ bl_0_494 br_0_494 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c494
+ bl_0_494 br_0_494 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c494
+ bl_0_494 br_0_494 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c494
+ bl_0_494 br_0_494 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c494
+ bl_0_494 br_0_494 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c494
+ bl_0_494 br_0_494 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c494
+ bl_0_494 br_0_494 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c494
+ bl_0_494 br_0_494 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c494
+ bl_0_494 br_0_494 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c494
+ bl_0_494 br_0_494 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c494
+ bl_0_494 br_0_494 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c494
+ bl_0_494 br_0_494 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c494
+ bl_0_494 br_0_494 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c494
+ bl_0_494 br_0_494 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c494
+ bl_0_494 br_0_494 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c494
+ bl_0_494 br_0_494 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c494
+ bl_0_494 br_0_494 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c494
+ bl_0_494 br_0_494 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c494
+ bl_0_494 br_0_494 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c494
+ bl_0_494 br_0_494 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c494
+ bl_0_494 br_0_494 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c494
+ bl_0_494 br_0_494 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c494
+ bl_0_494 br_0_494 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c494
+ bl_0_494 br_0_494 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c494
+ bl_0_494 br_0_494 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c494
+ bl_0_494 br_0_494 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c494
+ bl_0_494 br_0_494 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c494
+ bl_0_494 br_0_494 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c494
+ bl_0_494 br_0_494 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c494
+ bl_0_494 br_0_494 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c494
+ bl_0_494 br_0_494 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c494
+ bl_0_494 br_0_494 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c494
+ bl_0_494 br_0_494 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c494
+ bl_0_494 br_0_494 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c494
+ bl_0_494 br_0_494 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c494
+ bl_0_494 br_0_494 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c494
+ bl_0_494 br_0_494 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c494
+ bl_0_494 br_0_494 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c494
+ bl_0_494 br_0_494 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c494
+ bl_0_494 br_0_494 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c494
+ bl_0_494 br_0_494 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c494
+ bl_0_494 br_0_494 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c494
+ bl_0_494 br_0_494 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c494
+ bl_0_494 br_0_494 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c494
+ bl_0_494 br_0_494 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c495
+ bl_0_495 br_0_495 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c495
+ bl_0_495 br_0_495 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c495
+ bl_0_495 br_0_495 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c495
+ bl_0_495 br_0_495 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c495
+ bl_0_495 br_0_495 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c495
+ bl_0_495 br_0_495 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c495
+ bl_0_495 br_0_495 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c495
+ bl_0_495 br_0_495 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c495
+ bl_0_495 br_0_495 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c495
+ bl_0_495 br_0_495 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c495
+ bl_0_495 br_0_495 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c495
+ bl_0_495 br_0_495 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c495
+ bl_0_495 br_0_495 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c495
+ bl_0_495 br_0_495 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c495
+ bl_0_495 br_0_495 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c495
+ bl_0_495 br_0_495 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c495
+ bl_0_495 br_0_495 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c495
+ bl_0_495 br_0_495 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c495
+ bl_0_495 br_0_495 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c495
+ bl_0_495 br_0_495 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c495
+ bl_0_495 br_0_495 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c495
+ bl_0_495 br_0_495 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c495
+ bl_0_495 br_0_495 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c495
+ bl_0_495 br_0_495 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c495
+ bl_0_495 br_0_495 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c495
+ bl_0_495 br_0_495 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c495
+ bl_0_495 br_0_495 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c495
+ bl_0_495 br_0_495 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c495
+ bl_0_495 br_0_495 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c495
+ bl_0_495 br_0_495 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c495
+ bl_0_495 br_0_495 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c495
+ bl_0_495 br_0_495 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c495
+ bl_0_495 br_0_495 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c495
+ bl_0_495 br_0_495 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c495
+ bl_0_495 br_0_495 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c495
+ bl_0_495 br_0_495 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c495
+ bl_0_495 br_0_495 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c495
+ bl_0_495 br_0_495 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c495
+ bl_0_495 br_0_495 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c495
+ bl_0_495 br_0_495 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c495
+ bl_0_495 br_0_495 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c495
+ bl_0_495 br_0_495 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c495
+ bl_0_495 br_0_495 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c495
+ bl_0_495 br_0_495 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c495
+ bl_0_495 br_0_495 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c496
+ bl_0_496 br_0_496 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c496
+ bl_0_496 br_0_496 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c496
+ bl_0_496 br_0_496 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c496
+ bl_0_496 br_0_496 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c496
+ bl_0_496 br_0_496 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c496
+ bl_0_496 br_0_496 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c496
+ bl_0_496 br_0_496 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c496
+ bl_0_496 br_0_496 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c496
+ bl_0_496 br_0_496 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c496
+ bl_0_496 br_0_496 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c496
+ bl_0_496 br_0_496 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c496
+ bl_0_496 br_0_496 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c496
+ bl_0_496 br_0_496 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c496
+ bl_0_496 br_0_496 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c496
+ bl_0_496 br_0_496 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c496
+ bl_0_496 br_0_496 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c496
+ bl_0_496 br_0_496 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c496
+ bl_0_496 br_0_496 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c496
+ bl_0_496 br_0_496 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c496
+ bl_0_496 br_0_496 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c496
+ bl_0_496 br_0_496 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c496
+ bl_0_496 br_0_496 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c496
+ bl_0_496 br_0_496 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c496
+ bl_0_496 br_0_496 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c496
+ bl_0_496 br_0_496 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c496
+ bl_0_496 br_0_496 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c496
+ bl_0_496 br_0_496 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c496
+ bl_0_496 br_0_496 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c496
+ bl_0_496 br_0_496 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c496
+ bl_0_496 br_0_496 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c496
+ bl_0_496 br_0_496 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c496
+ bl_0_496 br_0_496 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c496
+ bl_0_496 br_0_496 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c496
+ bl_0_496 br_0_496 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c496
+ bl_0_496 br_0_496 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c496
+ bl_0_496 br_0_496 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c496
+ bl_0_496 br_0_496 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c496
+ bl_0_496 br_0_496 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c496
+ bl_0_496 br_0_496 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c496
+ bl_0_496 br_0_496 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c496
+ bl_0_496 br_0_496 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c496
+ bl_0_496 br_0_496 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c496
+ bl_0_496 br_0_496 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c496
+ bl_0_496 br_0_496 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c496
+ bl_0_496 br_0_496 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c497
+ bl_0_497 br_0_497 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c497
+ bl_0_497 br_0_497 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c497
+ bl_0_497 br_0_497 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c497
+ bl_0_497 br_0_497 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c497
+ bl_0_497 br_0_497 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c497
+ bl_0_497 br_0_497 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c497
+ bl_0_497 br_0_497 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c497
+ bl_0_497 br_0_497 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c497
+ bl_0_497 br_0_497 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c497
+ bl_0_497 br_0_497 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c497
+ bl_0_497 br_0_497 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c497
+ bl_0_497 br_0_497 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c497
+ bl_0_497 br_0_497 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c497
+ bl_0_497 br_0_497 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c497
+ bl_0_497 br_0_497 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c497
+ bl_0_497 br_0_497 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c497
+ bl_0_497 br_0_497 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c497
+ bl_0_497 br_0_497 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c497
+ bl_0_497 br_0_497 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c497
+ bl_0_497 br_0_497 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c497
+ bl_0_497 br_0_497 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c497
+ bl_0_497 br_0_497 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c497
+ bl_0_497 br_0_497 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c497
+ bl_0_497 br_0_497 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c497
+ bl_0_497 br_0_497 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c497
+ bl_0_497 br_0_497 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c497
+ bl_0_497 br_0_497 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c497
+ bl_0_497 br_0_497 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c497
+ bl_0_497 br_0_497 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c497
+ bl_0_497 br_0_497 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c497
+ bl_0_497 br_0_497 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c497
+ bl_0_497 br_0_497 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c497
+ bl_0_497 br_0_497 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c497
+ bl_0_497 br_0_497 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c497
+ bl_0_497 br_0_497 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c497
+ bl_0_497 br_0_497 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c497
+ bl_0_497 br_0_497 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c497
+ bl_0_497 br_0_497 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c497
+ bl_0_497 br_0_497 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c497
+ bl_0_497 br_0_497 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c497
+ bl_0_497 br_0_497 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c497
+ bl_0_497 br_0_497 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c497
+ bl_0_497 br_0_497 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c497
+ bl_0_497 br_0_497 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c497
+ bl_0_497 br_0_497 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c498
+ bl_0_498 br_0_498 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c498
+ bl_0_498 br_0_498 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c498
+ bl_0_498 br_0_498 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c498
+ bl_0_498 br_0_498 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c498
+ bl_0_498 br_0_498 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c498
+ bl_0_498 br_0_498 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c498
+ bl_0_498 br_0_498 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c498
+ bl_0_498 br_0_498 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c498
+ bl_0_498 br_0_498 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c498
+ bl_0_498 br_0_498 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c498
+ bl_0_498 br_0_498 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c498
+ bl_0_498 br_0_498 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c498
+ bl_0_498 br_0_498 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c498
+ bl_0_498 br_0_498 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c498
+ bl_0_498 br_0_498 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c498
+ bl_0_498 br_0_498 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c498
+ bl_0_498 br_0_498 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c498
+ bl_0_498 br_0_498 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c498
+ bl_0_498 br_0_498 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c498
+ bl_0_498 br_0_498 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c498
+ bl_0_498 br_0_498 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c498
+ bl_0_498 br_0_498 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c498
+ bl_0_498 br_0_498 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c498
+ bl_0_498 br_0_498 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c498
+ bl_0_498 br_0_498 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c498
+ bl_0_498 br_0_498 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c498
+ bl_0_498 br_0_498 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c498
+ bl_0_498 br_0_498 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c498
+ bl_0_498 br_0_498 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c498
+ bl_0_498 br_0_498 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c498
+ bl_0_498 br_0_498 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c498
+ bl_0_498 br_0_498 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c498
+ bl_0_498 br_0_498 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c498
+ bl_0_498 br_0_498 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c498
+ bl_0_498 br_0_498 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c498
+ bl_0_498 br_0_498 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c498
+ bl_0_498 br_0_498 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c498
+ bl_0_498 br_0_498 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c498
+ bl_0_498 br_0_498 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c498
+ bl_0_498 br_0_498 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c498
+ bl_0_498 br_0_498 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c498
+ bl_0_498 br_0_498 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c498
+ bl_0_498 br_0_498 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c498
+ bl_0_498 br_0_498 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c498
+ bl_0_498 br_0_498 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c499
+ bl_0_499 br_0_499 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c499
+ bl_0_499 br_0_499 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c499
+ bl_0_499 br_0_499 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c499
+ bl_0_499 br_0_499 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c499
+ bl_0_499 br_0_499 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c499
+ bl_0_499 br_0_499 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c499
+ bl_0_499 br_0_499 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c499
+ bl_0_499 br_0_499 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c499
+ bl_0_499 br_0_499 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c499
+ bl_0_499 br_0_499 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c499
+ bl_0_499 br_0_499 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c499
+ bl_0_499 br_0_499 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c499
+ bl_0_499 br_0_499 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c499
+ bl_0_499 br_0_499 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c499
+ bl_0_499 br_0_499 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c499
+ bl_0_499 br_0_499 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c499
+ bl_0_499 br_0_499 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c499
+ bl_0_499 br_0_499 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c499
+ bl_0_499 br_0_499 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c499
+ bl_0_499 br_0_499 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c499
+ bl_0_499 br_0_499 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c499
+ bl_0_499 br_0_499 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c499
+ bl_0_499 br_0_499 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c499
+ bl_0_499 br_0_499 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c499
+ bl_0_499 br_0_499 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c499
+ bl_0_499 br_0_499 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c499
+ bl_0_499 br_0_499 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c499
+ bl_0_499 br_0_499 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c499
+ bl_0_499 br_0_499 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c499
+ bl_0_499 br_0_499 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c499
+ bl_0_499 br_0_499 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c499
+ bl_0_499 br_0_499 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c499
+ bl_0_499 br_0_499 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c499
+ bl_0_499 br_0_499 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c499
+ bl_0_499 br_0_499 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c499
+ bl_0_499 br_0_499 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c499
+ bl_0_499 br_0_499 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c499
+ bl_0_499 br_0_499 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c499
+ bl_0_499 br_0_499 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c499
+ bl_0_499 br_0_499 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c499
+ bl_0_499 br_0_499 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c499
+ bl_0_499 br_0_499 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c499
+ bl_0_499 br_0_499 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c499
+ bl_0_499 br_0_499 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c499
+ bl_0_499 br_0_499 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c500
+ bl_0_500 br_0_500 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c500
+ bl_0_500 br_0_500 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c500
+ bl_0_500 br_0_500 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c500
+ bl_0_500 br_0_500 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c500
+ bl_0_500 br_0_500 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c500
+ bl_0_500 br_0_500 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c500
+ bl_0_500 br_0_500 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c500
+ bl_0_500 br_0_500 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c500
+ bl_0_500 br_0_500 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c500
+ bl_0_500 br_0_500 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c500
+ bl_0_500 br_0_500 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c500
+ bl_0_500 br_0_500 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c500
+ bl_0_500 br_0_500 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c500
+ bl_0_500 br_0_500 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c500
+ bl_0_500 br_0_500 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c500
+ bl_0_500 br_0_500 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c500
+ bl_0_500 br_0_500 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c500
+ bl_0_500 br_0_500 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c500
+ bl_0_500 br_0_500 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c500
+ bl_0_500 br_0_500 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c500
+ bl_0_500 br_0_500 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c500
+ bl_0_500 br_0_500 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c500
+ bl_0_500 br_0_500 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c500
+ bl_0_500 br_0_500 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c500
+ bl_0_500 br_0_500 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c500
+ bl_0_500 br_0_500 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c500
+ bl_0_500 br_0_500 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c500
+ bl_0_500 br_0_500 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c500
+ bl_0_500 br_0_500 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c500
+ bl_0_500 br_0_500 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c500
+ bl_0_500 br_0_500 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c500
+ bl_0_500 br_0_500 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c500
+ bl_0_500 br_0_500 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c500
+ bl_0_500 br_0_500 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c500
+ bl_0_500 br_0_500 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c500
+ bl_0_500 br_0_500 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c500
+ bl_0_500 br_0_500 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c500
+ bl_0_500 br_0_500 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c500
+ bl_0_500 br_0_500 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c500
+ bl_0_500 br_0_500 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c500
+ bl_0_500 br_0_500 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c500
+ bl_0_500 br_0_500 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c500
+ bl_0_500 br_0_500 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c500
+ bl_0_500 br_0_500 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c500
+ bl_0_500 br_0_500 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c501
+ bl_0_501 br_0_501 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c501
+ bl_0_501 br_0_501 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c501
+ bl_0_501 br_0_501 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c501
+ bl_0_501 br_0_501 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c501
+ bl_0_501 br_0_501 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c501
+ bl_0_501 br_0_501 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c501
+ bl_0_501 br_0_501 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c501
+ bl_0_501 br_0_501 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c501
+ bl_0_501 br_0_501 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c501
+ bl_0_501 br_0_501 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c501
+ bl_0_501 br_0_501 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c501
+ bl_0_501 br_0_501 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c501
+ bl_0_501 br_0_501 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c501
+ bl_0_501 br_0_501 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c501
+ bl_0_501 br_0_501 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c501
+ bl_0_501 br_0_501 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c501
+ bl_0_501 br_0_501 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c501
+ bl_0_501 br_0_501 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c501
+ bl_0_501 br_0_501 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c501
+ bl_0_501 br_0_501 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c501
+ bl_0_501 br_0_501 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c501
+ bl_0_501 br_0_501 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c501
+ bl_0_501 br_0_501 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c501
+ bl_0_501 br_0_501 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c501
+ bl_0_501 br_0_501 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c501
+ bl_0_501 br_0_501 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c501
+ bl_0_501 br_0_501 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c501
+ bl_0_501 br_0_501 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c501
+ bl_0_501 br_0_501 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c501
+ bl_0_501 br_0_501 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c501
+ bl_0_501 br_0_501 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c501
+ bl_0_501 br_0_501 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c501
+ bl_0_501 br_0_501 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c501
+ bl_0_501 br_0_501 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c501
+ bl_0_501 br_0_501 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c501
+ bl_0_501 br_0_501 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c501
+ bl_0_501 br_0_501 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c501
+ bl_0_501 br_0_501 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c501
+ bl_0_501 br_0_501 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c501
+ bl_0_501 br_0_501 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c501
+ bl_0_501 br_0_501 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c501
+ bl_0_501 br_0_501 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c501
+ bl_0_501 br_0_501 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c501
+ bl_0_501 br_0_501 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c501
+ bl_0_501 br_0_501 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c502
+ bl_0_502 br_0_502 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c502
+ bl_0_502 br_0_502 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c502
+ bl_0_502 br_0_502 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c502
+ bl_0_502 br_0_502 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c502
+ bl_0_502 br_0_502 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c502
+ bl_0_502 br_0_502 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c502
+ bl_0_502 br_0_502 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c502
+ bl_0_502 br_0_502 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c502
+ bl_0_502 br_0_502 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c502
+ bl_0_502 br_0_502 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c502
+ bl_0_502 br_0_502 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c502
+ bl_0_502 br_0_502 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c502
+ bl_0_502 br_0_502 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c502
+ bl_0_502 br_0_502 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c502
+ bl_0_502 br_0_502 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c502
+ bl_0_502 br_0_502 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c502
+ bl_0_502 br_0_502 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c502
+ bl_0_502 br_0_502 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c502
+ bl_0_502 br_0_502 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c502
+ bl_0_502 br_0_502 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c502
+ bl_0_502 br_0_502 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c502
+ bl_0_502 br_0_502 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c502
+ bl_0_502 br_0_502 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c502
+ bl_0_502 br_0_502 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c502
+ bl_0_502 br_0_502 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c502
+ bl_0_502 br_0_502 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c502
+ bl_0_502 br_0_502 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c502
+ bl_0_502 br_0_502 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c502
+ bl_0_502 br_0_502 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c502
+ bl_0_502 br_0_502 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c502
+ bl_0_502 br_0_502 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c502
+ bl_0_502 br_0_502 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c502
+ bl_0_502 br_0_502 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c502
+ bl_0_502 br_0_502 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c502
+ bl_0_502 br_0_502 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c502
+ bl_0_502 br_0_502 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c502
+ bl_0_502 br_0_502 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c502
+ bl_0_502 br_0_502 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c502
+ bl_0_502 br_0_502 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c502
+ bl_0_502 br_0_502 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c502
+ bl_0_502 br_0_502 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c502
+ bl_0_502 br_0_502 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c502
+ bl_0_502 br_0_502 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c502
+ bl_0_502 br_0_502 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c502
+ bl_0_502 br_0_502 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c503
+ bl_0_503 br_0_503 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c503
+ bl_0_503 br_0_503 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c503
+ bl_0_503 br_0_503 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c503
+ bl_0_503 br_0_503 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c503
+ bl_0_503 br_0_503 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c503
+ bl_0_503 br_0_503 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c503
+ bl_0_503 br_0_503 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c503
+ bl_0_503 br_0_503 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c503
+ bl_0_503 br_0_503 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c503
+ bl_0_503 br_0_503 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c503
+ bl_0_503 br_0_503 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c503
+ bl_0_503 br_0_503 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c503
+ bl_0_503 br_0_503 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c503
+ bl_0_503 br_0_503 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c503
+ bl_0_503 br_0_503 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c503
+ bl_0_503 br_0_503 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c503
+ bl_0_503 br_0_503 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c503
+ bl_0_503 br_0_503 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c503
+ bl_0_503 br_0_503 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c503
+ bl_0_503 br_0_503 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c503
+ bl_0_503 br_0_503 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c503
+ bl_0_503 br_0_503 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c503
+ bl_0_503 br_0_503 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c503
+ bl_0_503 br_0_503 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c503
+ bl_0_503 br_0_503 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c503
+ bl_0_503 br_0_503 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c503
+ bl_0_503 br_0_503 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c503
+ bl_0_503 br_0_503 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c503
+ bl_0_503 br_0_503 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c503
+ bl_0_503 br_0_503 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c503
+ bl_0_503 br_0_503 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c503
+ bl_0_503 br_0_503 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c503
+ bl_0_503 br_0_503 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c503
+ bl_0_503 br_0_503 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c503
+ bl_0_503 br_0_503 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c503
+ bl_0_503 br_0_503 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c503
+ bl_0_503 br_0_503 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c503
+ bl_0_503 br_0_503 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c503
+ bl_0_503 br_0_503 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c503
+ bl_0_503 br_0_503 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c503
+ bl_0_503 br_0_503 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c503
+ bl_0_503 br_0_503 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c503
+ bl_0_503 br_0_503 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c503
+ bl_0_503 br_0_503 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c503
+ bl_0_503 br_0_503 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c504
+ bl_0_504 br_0_504 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c504
+ bl_0_504 br_0_504 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c504
+ bl_0_504 br_0_504 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c504
+ bl_0_504 br_0_504 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c504
+ bl_0_504 br_0_504 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c504
+ bl_0_504 br_0_504 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c504
+ bl_0_504 br_0_504 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c504
+ bl_0_504 br_0_504 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c504
+ bl_0_504 br_0_504 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c504
+ bl_0_504 br_0_504 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c504
+ bl_0_504 br_0_504 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c504
+ bl_0_504 br_0_504 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c504
+ bl_0_504 br_0_504 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c504
+ bl_0_504 br_0_504 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c504
+ bl_0_504 br_0_504 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c504
+ bl_0_504 br_0_504 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c504
+ bl_0_504 br_0_504 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c504
+ bl_0_504 br_0_504 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c504
+ bl_0_504 br_0_504 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c504
+ bl_0_504 br_0_504 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c504
+ bl_0_504 br_0_504 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c504
+ bl_0_504 br_0_504 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c504
+ bl_0_504 br_0_504 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c504
+ bl_0_504 br_0_504 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c504
+ bl_0_504 br_0_504 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c504
+ bl_0_504 br_0_504 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c504
+ bl_0_504 br_0_504 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c504
+ bl_0_504 br_0_504 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c504
+ bl_0_504 br_0_504 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c504
+ bl_0_504 br_0_504 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c504
+ bl_0_504 br_0_504 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c504
+ bl_0_504 br_0_504 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c504
+ bl_0_504 br_0_504 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c504
+ bl_0_504 br_0_504 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c504
+ bl_0_504 br_0_504 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c504
+ bl_0_504 br_0_504 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c504
+ bl_0_504 br_0_504 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c504
+ bl_0_504 br_0_504 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c504
+ bl_0_504 br_0_504 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c504
+ bl_0_504 br_0_504 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c504
+ bl_0_504 br_0_504 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c504
+ bl_0_504 br_0_504 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c504
+ bl_0_504 br_0_504 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c504
+ bl_0_504 br_0_504 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c504
+ bl_0_504 br_0_504 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c505
+ bl_0_505 br_0_505 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c505
+ bl_0_505 br_0_505 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c505
+ bl_0_505 br_0_505 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c505
+ bl_0_505 br_0_505 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c505
+ bl_0_505 br_0_505 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c505
+ bl_0_505 br_0_505 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c505
+ bl_0_505 br_0_505 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c505
+ bl_0_505 br_0_505 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c505
+ bl_0_505 br_0_505 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c505
+ bl_0_505 br_0_505 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c505
+ bl_0_505 br_0_505 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c505
+ bl_0_505 br_0_505 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c505
+ bl_0_505 br_0_505 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c505
+ bl_0_505 br_0_505 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c505
+ bl_0_505 br_0_505 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c505
+ bl_0_505 br_0_505 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c505
+ bl_0_505 br_0_505 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c505
+ bl_0_505 br_0_505 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c505
+ bl_0_505 br_0_505 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c505
+ bl_0_505 br_0_505 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c505
+ bl_0_505 br_0_505 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c505
+ bl_0_505 br_0_505 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c505
+ bl_0_505 br_0_505 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c505
+ bl_0_505 br_0_505 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c505
+ bl_0_505 br_0_505 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c505
+ bl_0_505 br_0_505 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c505
+ bl_0_505 br_0_505 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c505
+ bl_0_505 br_0_505 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c505
+ bl_0_505 br_0_505 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c505
+ bl_0_505 br_0_505 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c505
+ bl_0_505 br_0_505 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c505
+ bl_0_505 br_0_505 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c505
+ bl_0_505 br_0_505 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c505
+ bl_0_505 br_0_505 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c505
+ bl_0_505 br_0_505 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c505
+ bl_0_505 br_0_505 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c505
+ bl_0_505 br_0_505 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c505
+ bl_0_505 br_0_505 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c505
+ bl_0_505 br_0_505 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c505
+ bl_0_505 br_0_505 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c505
+ bl_0_505 br_0_505 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c505
+ bl_0_505 br_0_505 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c505
+ bl_0_505 br_0_505 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c505
+ bl_0_505 br_0_505 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c505
+ bl_0_505 br_0_505 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c506
+ bl_0_506 br_0_506 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c506
+ bl_0_506 br_0_506 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c506
+ bl_0_506 br_0_506 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c506
+ bl_0_506 br_0_506 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c506
+ bl_0_506 br_0_506 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c506
+ bl_0_506 br_0_506 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c506
+ bl_0_506 br_0_506 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c506
+ bl_0_506 br_0_506 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c506
+ bl_0_506 br_0_506 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c506
+ bl_0_506 br_0_506 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c506
+ bl_0_506 br_0_506 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c506
+ bl_0_506 br_0_506 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c506
+ bl_0_506 br_0_506 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c506
+ bl_0_506 br_0_506 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c506
+ bl_0_506 br_0_506 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c506
+ bl_0_506 br_0_506 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c506
+ bl_0_506 br_0_506 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c506
+ bl_0_506 br_0_506 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c506
+ bl_0_506 br_0_506 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c506
+ bl_0_506 br_0_506 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c506
+ bl_0_506 br_0_506 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c506
+ bl_0_506 br_0_506 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c506
+ bl_0_506 br_0_506 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c506
+ bl_0_506 br_0_506 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c506
+ bl_0_506 br_0_506 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c506
+ bl_0_506 br_0_506 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c506
+ bl_0_506 br_0_506 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c506
+ bl_0_506 br_0_506 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c506
+ bl_0_506 br_0_506 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c506
+ bl_0_506 br_0_506 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c506
+ bl_0_506 br_0_506 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c506
+ bl_0_506 br_0_506 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c506
+ bl_0_506 br_0_506 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c506
+ bl_0_506 br_0_506 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c506
+ bl_0_506 br_0_506 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c506
+ bl_0_506 br_0_506 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c506
+ bl_0_506 br_0_506 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c506
+ bl_0_506 br_0_506 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c506
+ bl_0_506 br_0_506 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c506
+ bl_0_506 br_0_506 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c506
+ bl_0_506 br_0_506 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c506
+ bl_0_506 br_0_506 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c506
+ bl_0_506 br_0_506 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c506
+ bl_0_506 br_0_506 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c506
+ bl_0_506 br_0_506 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c507
+ bl_0_507 br_0_507 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c507
+ bl_0_507 br_0_507 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c507
+ bl_0_507 br_0_507 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c507
+ bl_0_507 br_0_507 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c507
+ bl_0_507 br_0_507 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c507
+ bl_0_507 br_0_507 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c507
+ bl_0_507 br_0_507 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c507
+ bl_0_507 br_0_507 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c507
+ bl_0_507 br_0_507 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c507
+ bl_0_507 br_0_507 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c507
+ bl_0_507 br_0_507 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c507
+ bl_0_507 br_0_507 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c507
+ bl_0_507 br_0_507 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c507
+ bl_0_507 br_0_507 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c507
+ bl_0_507 br_0_507 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c507
+ bl_0_507 br_0_507 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c507
+ bl_0_507 br_0_507 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c507
+ bl_0_507 br_0_507 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c507
+ bl_0_507 br_0_507 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c507
+ bl_0_507 br_0_507 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c507
+ bl_0_507 br_0_507 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c507
+ bl_0_507 br_0_507 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c507
+ bl_0_507 br_0_507 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c507
+ bl_0_507 br_0_507 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c507
+ bl_0_507 br_0_507 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c507
+ bl_0_507 br_0_507 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c507
+ bl_0_507 br_0_507 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c507
+ bl_0_507 br_0_507 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c507
+ bl_0_507 br_0_507 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c507
+ bl_0_507 br_0_507 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c507
+ bl_0_507 br_0_507 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c507
+ bl_0_507 br_0_507 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c507
+ bl_0_507 br_0_507 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c507
+ bl_0_507 br_0_507 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c507
+ bl_0_507 br_0_507 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c507
+ bl_0_507 br_0_507 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c507
+ bl_0_507 br_0_507 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c507
+ bl_0_507 br_0_507 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c507
+ bl_0_507 br_0_507 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c507
+ bl_0_507 br_0_507 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c507
+ bl_0_507 br_0_507 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c507
+ bl_0_507 br_0_507 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c507
+ bl_0_507 br_0_507 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c507
+ bl_0_507 br_0_507 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c507
+ bl_0_507 br_0_507 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c508
+ bl_0_508 br_0_508 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c508
+ bl_0_508 br_0_508 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c508
+ bl_0_508 br_0_508 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c508
+ bl_0_508 br_0_508 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c508
+ bl_0_508 br_0_508 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c508
+ bl_0_508 br_0_508 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c508
+ bl_0_508 br_0_508 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c508
+ bl_0_508 br_0_508 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c508
+ bl_0_508 br_0_508 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c508
+ bl_0_508 br_0_508 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c508
+ bl_0_508 br_0_508 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c508
+ bl_0_508 br_0_508 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c508
+ bl_0_508 br_0_508 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c508
+ bl_0_508 br_0_508 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c508
+ bl_0_508 br_0_508 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c508
+ bl_0_508 br_0_508 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c508
+ bl_0_508 br_0_508 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c508
+ bl_0_508 br_0_508 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c508
+ bl_0_508 br_0_508 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c508
+ bl_0_508 br_0_508 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c508
+ bl_0_508 br_0_508 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c508
+ bl_0_508 br_0_508 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c508
+ bl_0_508 br_0_508 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c508
+ bl_0_508 br_0_508 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c508
+ bl_0_508 br_0_508 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c508
+ bl_0_508 br_0_508 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c508
+ bl_0_508 br_0_508 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c508
+ bl_0_508 br_0_508 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c508
+ bl_0_508 br_0_508 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c508
+ bl_0_508 br_0_508 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c508
+ bl_0_508 br_0_508 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c508
+ bl_0_508 br_0_508 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c508
+ bl_0_508 br_0_508 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c508
+ bl_0_508 br_0_508 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c508
+ bl_0_508 br_0_508 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c508
+ bl_0_508 br_0_508 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c508
+ bl_0_508 br_0_508 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c508
+ bl_0_508 br_0_508 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c508
+ bl_0_508 br_0_508 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c508
+ bl_0_508 br_0_508 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c508
+ bl_0_508 br_0_508 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c508
+ bl_0_508 br_0_508 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c508
+ bl_0_508 br_0_508 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c508
+ bl_0_508 br_0_508 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c508
+ bl_0_508 br_0_508 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c509
+ bl_0_509 br_0_509 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c509
+ bl_0_509 br_0_509 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c509
+ bl_0_509 br_0_509 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c509
+ bl_0_509 br_0_509 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c509
+ bl_0_509 br_0_509 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c509
+ bl_0_509 br_0_509 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c509
+ bl_0_509 br_0_509 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c509
+ bl_0_509 br_0_509 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c509
+ bl_0_509 br_0_509 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c509
+ bl_0_509 br_0_509 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c509
+ bl_0_509 br_0_509 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c509
+ bl_0_509 br_0_509 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c509
+ bl_0_509 br_0_509 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c509
+ bl_0_509 br_0_509 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c509
+ bl_0_509 br_0_509 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c509
+ bl_0_509 br_0_509 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c509
+ bl_0_509 br_0_509 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c509
+ bl_0_509 br_0_509 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c509
+ bl_0_509 br_0_509 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c509
+ bl_0_509 br_0_509 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c509
+ bl_0_509 br_0_509 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c509
+ bl_0_509 br_0_509 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c509
+ bl_0_509 br_0_509 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c509
+ bl_0_509 br_0_509 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c509
+ bl_0_509 br_0_509 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c509
+ bl_0_509 br_0_509 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c509
+ bl_0_509 br_0_509 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c509
+ bl_0_509 br_0_509 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c509
+ bl_0_509 br_0_509 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c509
+ bl_0_509 br_0_509 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c509
+ bl_0_509 br_0_509 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c509
+ bl_0_509 br_0_509 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c509
+ bl_0_509 br_0_509 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c509
+ bl_0_509 br_0_509 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c509
+ bl_0_509 br_0_509 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c509
+ bl_0_509 br_0_509 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c509
+ bl_0_509 br_0_509 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c509
+ bl_0_509 br_0_509 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c509
+ bl_0_509 br_0_509 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c509
+ bl_0_509 br_0_509 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c509
+ bl_0_509 br_0_509 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c509
+ bl_0_509 br_0_509 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c509
+ bl_0_509 br_0_509 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c509
+ bl_0_509 br_0_509 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c509
+ bl_0_509 br_0_509 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c510
+ bl_0_510 br_0_510 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c510
+ bl_0_510 br_0_510 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c510
+ bl_0_510 br_0_510 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c510
+ bl_0_510 br_0_510 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c510
+ bl_0_510 br_0_510 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c510
+ bl_0_510 br_0_510 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c510
+ bl_0_510 br_0_510 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c510
+ bl_0_510 br_0_510 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c510
+ bl_0_510 br_0_510 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c510
+ bl_0_510 br_0_510 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c510
+ bl_0_510 br_0_510 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c510
+ bl_0_510 br_0_510 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c510
+ bl_0_510 br_0_510 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c510
+ bl_0_510 br_0_510 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c510
+ bl_0_510 br_0_510 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c510
+ bl_0_510 br_0_510 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c510
+ bl_0_510 br_0_510 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c510
+ bl_0_510 br_0_510 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c510
+ bl_0_510 br_0_510 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c510
+ bl_0_510 br_0_510 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c510
+ bl_0_510 br_0_510 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c510
+ bl_0_510 br_0_510 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c510
+ bl_0_510 br_0_510 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c510
+ bl_0_510 br_0_510 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c510
+ bl_0_510 br_0_510 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c510
+ bl_0_510 br_0_510 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c510
+ bl_0_510 br_0_510 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c510
+ bl_0_510 br_0_510 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c510
+ bl_0_510 br_0_510 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c510
+ bl_0_510 br_0_510 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c510
+ bl_0_510 br_0_510 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c510
+ bl_0_510 br_0_510 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c510
+ bl_0_510 br_0_510 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c510
+ bl_0_510 br_0_510 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c510
+ bl_0_510 br_0_510 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c510
+ bl_0_510 br_0_510 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c510
+ bl_0_510 br_0_510 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c510
+ bl_0_510 br_0_510 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c510
+ bl_0_510 br_0_510 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c510
+ bl_0_510 br_0_510 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c510
+ bl_0_510 br_0_510 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c510
+ bl_0_510 br_0_510 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c510
+ bl_0_510 br_0_510 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c510
+ bl_0_510 br_0_510 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c510
+ bl_0_510 br_0_510 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r0_c511
+ bl_0_511 br_0_511 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c511
+ bl_0_511 br_0_511 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c511
+ bl_0_511 br_0_511 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c511
+ bl_0_511 br_0_511 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c511
+ bl_0_511 br_0_511 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c511
+ bl_0_511 br_0_511 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c511
+ bl_0_511 br_0_511 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c511
+ bl_0_511 br_0_511 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c511
+ bl_0_511 br_0_511 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c511
+ bl_0_511 br_0_511 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c511
+ bl_0_511 br_0_511 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c511
+ bl_0_511 br_0_511 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c511
+ bl_0_511 br_0_511 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c511
+ bl_0_511 br_0_511 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c511
+ bl_0_511 br_0_511 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c511
+ bl_0_511 br_0_511 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c511
+ bl_0_511 br_0_511 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c511
+ bl_0_511 br_0_511 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c511
+ bl_0_511 br_0_511 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c511
+ bl_0_511 br_0_511 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c511
+ bl_0_511 br_0_511 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c511
+ bl_0_511 br_0_511 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c511
+ bl_0_511 br_0_511 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c511
+ bl_0_511 br_0_511 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c511
+ bl_0_511 br_0_511 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c511
+ bl_0_511 br_0_511 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c511
+ bl_0_511 br_0_511 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c511
+ bl_0_511 br_0_511 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c511
+ bl_0_511 br_0_511 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c511
+ bl_0_511 br_0_511 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c511
+ bl_0_511 br_0_511 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c511
+ bl_0_511 br_0_511 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c511
+ bl_0_511 br_0_511 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c511
+ bl_0_511 br_0_511 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c511
+ bl_0_511 br_0_511 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c511
+ bl_0_511 br_0_511 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c511
+ bl_0_511 br_0_511 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c511
+ bl_0_511 br_0_511 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c511
+ bl_0_511 br_0_511 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c511
+ bl_0_511 br_0_511 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c511
+ bl_0_511 br_0_511 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c511
+ bl_0_511 br_0_511 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c511
+ bl_0_511 br_0_511 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c511
+ bl_0_511 br_0_511 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c511
+ bl_0_511 br_0_511 wl_0_44 vdd gnd
+ cell_1rw
.ENDS freepdk45_sram_1rw0r_45x512_bitcell_array

.SUBCKT replica_cell_1rw bl br wl vdd gnd
* Inverter 1
MM0 vdd Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 vdd Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q vdd gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q vdd vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl vdd gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_1rw


.SUBCKT freepdk45_sram_1rw0r_45x512_replica_column
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 vdd gnd
* OUTPUT: bl_0_0 
* OUTPUT: br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* POWER : vdd 
* GROUND: gnd 
Xrbc_0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ replica_cell_1rw
Xrbc_1
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ replica_cell_1rw
Xrbc_2
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ replica_cell_1rw
Xrbc_3
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ replica_cell_1rw
Xrbc_4
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ replica_cell_1rw
Xrbc_5
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ replica_cell_1rw
Xrbc_6
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ replica_cell_1rw
Xrbc_7
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ replica_cell_1rw
Xrbc_8
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ replica_cell_1rw
Xrbc_9
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ replica_cell_1rw
Xrbc_10
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ replica_cell_1rw
Xrbc_11
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ replica_cell_1rw
Xrbc_12
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ replica_cell_1rw
Xrbc_13
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ replica_cell_1rw
Xrbc_14
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ replica_cell_1rw
Xrbc_15
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ replica_cell_1rw
Xrbc_16
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ replica_cell_1rw
Xrbc_17
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ replica_cell_1rw
Xrbc_18
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ replica_cell_1rw
Xrbc_19
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ replica_cell_1rw
Xrbc_20
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ replica_cell_1rw
Xrbc_21
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ replica_cell_1rw
Xrbc_22
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ replica_cell_1rw
Xrbc_23
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ replica_cell_1rw
Xrbc_24
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ replica_cell_1rw
Xrbc_25
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ replica_cell_1rw
Xrbc_26
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ replica_cell_1rw
Xrbc_27
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ replica_cell_1rw
Xrbc_28
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ replica_cell_1rw
Xrbc_29
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ replica_cell_1rw
Xrbc_30
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ replica_cell_1rw
Xrbc_31
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ replica_cell_1rw
Xrbc_32
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ replica_cell_1rw
Xrbc_33
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ replica_cell_1rw
Xrbc_34
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ replica_cell_1rw
Xrbc_35
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ replica_cell_1rw
Xrbc_36
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ replica_cell_1rw
Xrbc_37
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ replica_cell_1rw
Xrbc_38
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ replica_cell_1rw
Xrbc_39
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ replica_cell_1rw
Xrbc_40
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ replica_cell_1rw
Xrbc_41
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ replica_cell_1rw
Xrbc_42
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ replica_cell_1rw
Xrbc_43
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ replica_cell_1rw
Xrbc_44
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ replica_cell_1rw
Xrbc_45
+ bl_0_0 br_0_0 wl_0_45 vdd gnd
+ replica_cell_1rw
.ENDS freepdk45_sram_1rw0r_45x512_replica_column

.SUBCKT dummy_cell_1rw bl br wl vdd gnd
* Inverter 1
MM0 Q_bar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Q_bar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Q_bar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Q_bar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl_noconn wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br_noconn wl Q_bar gnd NMOS_VTG W=135.00n L=50n
.ENDS dummy_cell_1rw


.SUBCKT freepdk45_sram_1rw0r_45x512_dummy_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258 br_0_258 bl_0_259
+ br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261 bl_0_262 br_0_262
+ bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265 br_0_265 bl_0_266
+ br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268 bl_0_269 br_0_269
+ bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272 br_0_272 bl_0_273
+ br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275 bl_0_276 br_0_276
+ bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279 br_0_279 bl_0_280
+ br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282 bl_0_283 br_0_283
+ bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286 br_0_286 bl_0_287
+ br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289 bl_0_290 br_0_290
+ bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293 br_0_293 bl_0_294
+ br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296 bl_0_297 br_0_297
+ bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300 br_0_300 bl_0_301
+ br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303 bl_0_304 br_0_304
+ bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307 br_0_307 bl_0_308
+ br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310 bl_0_311 br_0_311
+ bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314 br_0_314 bl_0_315
+ br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317 bl_0_318 br_0_318
+ bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321 br_0_321 bl_0_322
+ br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324 bl_0_325 br_0_325
+ bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328 br_0_328 bl_0_329
+ br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331 bl_0_332 br_0_332
+ bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335 br_0_335 bl_0_336
+ br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338 bl_0_339 br_0_339
+ bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342 br_0_342 bl_0_343
+ br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345 bl_0_346 br_0_346
+ bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349 br_0_349 bl_0_350
+ br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352 bl_0_353 br_0_353
+ bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356 br_0_356 bl_0_357
+ br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359 bl_0_360 br_0_360
+ bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363 br_0_363 bl_0_364
+ br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366 bl_0_367 br_0_367
+ bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370 br_0_370 bl_0_371
+ br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373 bl_0_374 br_0_374
+ bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377 br_0_377 bl_0_378
+ br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380 bl_0_381 br_0_381
+ bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384 br_0_384 bl_0_385
+ br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387 bl_0_388 br_0_388
+ bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391 br_0_391 bl_0_392
+ br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394 bl_0_395 br_0_395
+ bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398 br_0_398 bl_0_399
+ br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401 bl_0_402 br_0_402
+ bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405 br_0_405 bl_0_406
+ br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408 bl_0_409 br_0_409
+ bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412 br_0_412 bl_0_413
+ br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415 bl_0_416 br_0_416
+ bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419 br_0_419 bl_0_420
+ br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422 bl_0_423 br_0_423
+ bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426 br_0_426 bl_0_427
+ br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429 bl_0_430 br_0_430
+ bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433 br_0_433 bl_0_434
+ br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436 bl_0_437 br_0_437
+ bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440 br_0_440 bl_0_441
+ br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443 bl_0_444 br_0_444
+ bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447 br_0_447 bl_0_448
+ br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450 bl_0_451 br_0_451
+ bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454 br_0_454 bl_0_455
+ br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457 bl_0_458 br_0_458
+ bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461 br_0_461 bl_0_462
+ br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464 bl_0_465 br_0_465
+ bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468 br_0_468 bl_0_469
+ br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471 bl_0_472 br_0_472
+ bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475 br_0_475 bl_0_476
+ br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478 bl_0_479 br_0_479
+ bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482 br_0_482 bl_0_483
+ br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485 bl_0_486 br_0_486
+ bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489 br_0_489 bl_0_490
+ br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492 bl_0_493 br_0_493
+ bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496 br_0_496 bl_0_497
+ br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499 bl_0_500 br_0_500
+ bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503 br_0_503 bl_0_504
+ br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506 bl_0_507 br_0_507
+ bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510 br_0_510 bl_0_511
+ br_0_511 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INOUT : bl_0_257 
* INOUT : br_0_257 
* INOUT : bl_0_258 
* INOUT : br_0_258 
* INOUT : bl_0_259 
* INOUT : br_0_259 
* INOUT : bl_0_260 
* INOUT : br_0_260 
* INOUT : bl_0_261 
* INOUT : br_0_261 
* INOUT : bl_0_262 
* INOUT : br_0_262 
* INOUT : bl_0_263 
* INOUT : br_0_263 
* INOUT : bl_0_264 
* INOUT : br_0_264 
* INOUT : bl_0_265 
* INOUT : br_0_265 
* INOUT : bl_0_266 
* INOUT : br_0_266 
* INOUT : bl_0_267 
* INOUT : br_0_267 
* INOUT : bl_0_268 
* INOUT : br_0_268 
* INOUT : bl_0_269 
* INOUT : br_0_269 
* INOUT : bl_0_270 
* INOUT : br_0_270 
* INOUT : bl_0_271 
* INOUT : br_0_271 
* INOUT : bl_0_272 
* INOUT : br_0_272 
* INOUT : bl_0_273 
* INOUT : br_0_273 
* INOUT : bl_0_274 
* INOUT : br_0_274 
* INOUT : bl_0_275 
* INOUT : br_0_275 
* INOUT : bl_0_276 
* INOUT : br_0_276 
* INOUT : bl_0_277 
* INOUT : br_0_277 
* INOUT : bl_0_278 
* INOUT : br_0_278 
* INOUT : bl_0_279 
* INOUT : br_0_279 
* INOUT : bl_0_280 
* INOUT : br_0_280 
* INOUT : bl_0_281 
* INOUT : br_0_281 
* INOUT : bl_0_282 
* INOUT : br_0_282 
* INOUT : bl_0_283 
* INOUT : br_0_283 
* INOUT : bl_0_284 
* INOUT : br_0_284 
* INOUT : bl_0_285 
* INOUT : br_0_285 
* INOUT : bl_0_286 
* INOUT : br_0_286 
* INOUT : bl_0_287 
* INOUT : br_0_287 
* INOUT : bl_0_288 
* INOUT : br_0_288 
* INOUT : bl_0_289 
* INOUT : br_0_289 
* INOUT : bl_0_290 
* INOUT : br_0_290 
* INOUT : bl_0_291 
* INOUT : br_0_291 
* INOUT : bl_0_292 
* INOUT : br_0_292 
* INOUT : bl_0_293 
* INOUT : br_0_293 
* INOUT : bl_0_294 
* INOUT : br_0_294 
* INOUT : bl_0_295 
* INOUT : br_0_295 
* INOUT : bl_0_296 
* INOUT : br_0_296 
* INOUT : bl_0_297 
* INOUT : br_0_297 
* INOUT : bl_0_298 
* INOUT : br_0_298 
* INOUT : bl_0_299 
* INOUT : br_0_299 
* INOUT : bl_0_300 
* INOUT : br_0_300 
* INOUT : bl_0_301 
* INOUT : br_0_301 
* INOUT : bl_0_302 
* INOUT : br_0_302 
* INOUT : bl_0_303 
* INOUT : br_0_303 
* INOUT : bl_0_304 
* INOUT : br_0_304 
* INOUT : bl_0_305 
* INOUT : br_0_305 
* INOUT : bl_0_306 
* INOUT : br_0_306 
* INOUT : bl_0_307 
* INOUT : br_0_307 
* INOUT : bl_0_308 
* INOUT : br_0_308 
* INOUT : bl_0_309 
* INOUT : br_0_309 
* INOUT : bl_0_310 
* INOUT : br_0_310 
* INOUT : bl_0_311 
* INOUT : br_0_311 
* INOUT : bl_0_312 
* INOUT : br_0_312 
* INOUT : bl_0_313 
* INOUT : br_0_313 
* INOUT : bl_0_314 
* INOUT : br_0_314 
* INOUT : bl_0_315 
* INOUT : br_0_315 
* INOUT : bl_0_316 
* INOUT : br_0_316 
* INOUT : bl_0_317 
* INOUT : br_0_317 
* INOUT : bl_0_318 
* INOUT : br_0_318 
* INOUT : bl_0_319 
* INOUT : br_0_319 
* INOUT : bl_0_320 
* INOUT : br_0_320 
* INOUT : bl_0_321 
* INOUT : br_0_321 
* INOUT : bl_0_322 
* INOUT : br_0_322 
* INOUT : bl_0_323 
* INOUT : br_0_323 
* INOUT : bl_0_324 
* INOUT : br_0_324 
* INOUT : bl_0_325 
* INOUT : br_0_325 
* INOUT : bl_0_326 
* INOUT : br_0_326 
* INOUT : bl_0_327 
* INOUT : br_0_327 
* INOUT : bl_0_328 
* INOUT : br_0_328 
* INOUT : bl_0_329 
* INOUT : br_0_329 
* INOUT : bl_0_330 
* INOUT : br_0_330 
* INOUT : bl_0_331 
* INOUT : br_0_331 
* INOUT : bl_0_332 
* INOUT : br_0_332 
* INOUT : bl_0_333 
* INOUT : br_0_333 
* INOUT : bl_0_334 
* INOUT : br_0_334 
* INOUT : bl_0_335 
* INOUT : br_0_335 
* INOUT : bl_0_336 
* INOUT : br_0_336 
* INOUT : bl_0_337 
* INOUT : br_0_337 
* INOUT : bl_0_338 
* INOUT : br_0_338 
* INOUT : bl_0_339 
* INOUT : br_0_339 
* INOUT : bl_0_340 
* INOUT : br_0_340 
* INOUT : bl_0_341 
* INOUT : br_0_341 
* INOUT : bl_0_342 
* INOUT : br_0_342 
* INOUT : bl_0_343 
* INOUT : br_0_343 
* INOUT : bl_0_344 
* INOUT : br_0_344 
* INOUT : bl_0_345 
* INOUT : br_0_345 
* INOUT : bl_0_346 
* INOUT : br_0_346 
* INOUT : bl_0_347 
* INOUT : br_0_347 
* INOUT : bl_0_348 
* INOUT : br_0_348 
* INOUT : bl_0_349 
* INOUT : br_0_349 
* INOUT : bl_0_350 
* INOUT : br_0_350 
* INOUT : bl_0_351 
* INOUT : br_0_351 
* INOUT : bl_0_352 
* INOUT : br_0_352 
* INOUT : bl_0_353 
* INOUT : br_0_353 
* INOUT : bl_0_354 
* INOUT : br_0_354 
* INOUT : bl_0_355 
* INOUT : br_0_355 
* INOUT : bl_0_356 
* INOUT : br_0_356 
* INOUT : bl_0_357 
* INOUT : br_0_357 
* INOUT : bl_0_358 
* INOUT : br_0_358 
* INOUT : bl_0_359 
* INOUT : br_0_359 
* INOUT : bl_0_360 
* INOUT : br_0_360 
* INOUT : bl_0_361 
* INOUT : br_0_361 
* INOUT : bl_0_362 
* INOUT : br_0_362 
* INOUT : bl_0_363 
* INOUT : br_0_363 
* INOUT : bl_0_364 
* INOUT : br_0_364 
* INOUT : bl_0_365 
* INOUT : br_0_365 
* INOUT : bl_0_366 
* INOUT : br_0_366 
* INOUT : bl_0_367 
* INOUT : br_0_367 
* INOUT : bl_0_368 
* INOUT : br_0_368 
* INOUT : bl_0_369 
* INOUT : br_0_369 
* INOUT : bl_0_370 
* INOUT : br_0_370 
* INOUT : bl_0_371 
* INOUT : br_0_371 
* INOUT : bl_0_372 
* INOUT : br_0_372 
* INOUT : bl_0_373 
* INOUT : br_0_373 
* INOUT : bl_0_374 
* INOUT : br_0_374 
* INOUT : bl_0_375 
* INOUT : br_0_375 
* INOUT : bl_0_376 
* INOUT : br_0_376 
* INOUT : bl_0_377 
* INOUT : br_0_377 
* INOUT : bl_0_378 
* INOUT : br_0_378 
* INOUT : bl_0_379 
* INOUT : br_0_379 
* INOUT : bl_0_380 
* INOUT : br_0_380 
* INOUT : bl_0_381 
* INOUT : br_0_381 
* INOUT : bl_0_382 
* INOUT : br_0_382 
* INOUT : bl_0_383 
* INOUT : br_0_383 
* INOUT : bl_0_384 
* INOUT : br_0_384 
* INOUT : bl_0_385 
* INOUT : br_0_385 
* INOUT : bl_0_386 
* INOUT : br_0_386 
* INOUT : bl_0_387 
* INOUT : br_0_387 
* INOUT : bl_0_388 
* INOUT : br_0_388 
* INOUT : bl_0_389 
* INOUT : br_0_389 
* INOUT : bl_0_390 
* INOUT : br_0_390 
* INOUT : bl_0_391 
* INOUT : br_0_391 
* INOUT : bl_0_392 
* INOUT : br_0_392 
* INOUT : bl_0_393 
* INOUT : br_0_393 
* INOUT : bl_0_394 
* INOUT : br_0_394 
* INOUT : bl_0_395 
* INOUT : br_0_395 
* INOUT : bl_0_396 
* INOUT : br_0_396 
* INOUT : bl_0_397 
* INOUT : br_0_397 
* INOUT : bl_0_398 
* INOUT : br_0_398 
* INOUT : bl_0_399 
* INOUT : br_0_399 
* INOUT : bl_0_400 
* INOUT : br_0_400 
* INOUT : bl_0_401 
* INOUT : br_0_401 
* INOUT : bl_0_402 
* INOUT : br_0_402 
* INOUT : bl_0_403 
* INOUT : br_0_403 
* INOUT : bl_0_404 
* INOUT : br_0_404 
* INOUT : bl_0_405 
* INOUT : br_0_405 
* INOUT : bl_0_406 
* INOUT : br_0_406 
* INOUT : bl_0_407 
* INOUT : br_0_407 
* INOUT : bl_0_408 
* INOUT : br_0_408 
* INOUT : bl_0_409 
* INOUT : br_0_409 
* INOUT : bl_0_410 
* INOUT : br_0_410 
* INOUT : bl_0_411 
* INOUT : br_0_411 
* INOUT : bl_0_412 
* INOUT : br_0_412 
* INOUT : bl_0_413 
* INOUT : br_0_413 
* INOUT : bl_0_414 
* INOUT : br_0_414 
* INOUT : bl_0_415 
* INOUT : br_0_415 
* INOUT : bl_0_416 
* INOUT : br_0_416 
* INOUT : bl_0_417 
* INOUT : br_0_417 
* INOUT : bl_0_418 
* INOUT : br_0_418 
* INOUT : bl_0_419 
* INOUT : br_0_419 
* INOUT : bl_0_420 
* INOUT : br_0_420 
* INOUT : bl_0_421 
* INOUT : br_0_421 
* INOUT : bl_0_422 
* INOUT : br_0_422 
* INOUT : bl_0_423 
* INOUT : br_0_423 
* INOUT : bl_0_424 
* INOUT : br_0_424 
* INOUT : bl_0_425 
* INOUT : br_0_425 
* INOUT : bl_0_426 
* INOUT : br_0_426 
* INOUT : bl_0_427 
* INOUT : br_0_427 
* INOUT : bl_0_428 
* INOUT : br_0_428 
* INOUT : bl_0_429 
* INOUT : br_0_429 
* INOUT : bl_0_430 
* INOUT : br_0_430 
* INOUT : bl_0_431 
* INOUT : br_0_431 
* INOUT : bl_0_432 
* INOUT : br_0_432 
* INOUT : bl_0_433 
* INOUT : br_0_433 
* INOUT : bl_0_434 
* INOUT : br_0_434 
* INOUT : bl_0_435 
* INOUT : br_0_435 
* INOUT : bl_0_436 
* INOUT : br_0_436 
* INOUT : bl_0_437 
* INOUT : br_0_437 
* INOUT : bl_0_438 
* INOUT : br_0_438 
* INOUT : bl_0_439 
* INOUT : br_0_439 
* INOUT : bl_0_440 
* INOUT : br_0_440 
* INOUT : bl_0_441 
* INOUT : br_0_441 
* INOUT : bl_0_442 
* INOUT : br_0_442 
* INOUT : bl_0_443 
* INOUT : br_0_443 
* INOUT : bl_0_444 
* INOUT : br_0_444 
* INOUT : bl_0_445 
* INOUT : br_0_445 
* INOUT : bl_0_446 
* INOUT : br_0_446 
* INOUT : bl_0_447 
* INOUT : br_0_447 
* INOUT : bl_0_448 
* INOUT : br_0_448 
* INOUT : bl_0_449 
* INOUT : br_0_449 
* INOUT : bl_0_450 
* INOUT : br_0_450 
* INOUT : bl_0_451 
* INOUT : br_0_451 
* INOUT : bl_0_452 
* INOUT : br_0_452 
* INOUT : bl_0_453 
* INOUT : br_0_453 
* INOUT : bl_0_454 
* INOUT : br_0_454 
* INOUT : bl_0_455 
* INOUT : br_0_455 
* INOUT : bl_0_456 
* INOUT : br_0_456 
* INOUT : bl_0_457 
* INOUT : br_0_457 
* INOUT : bl_0_458 
* INOUT : br_0_458 
* INOUT : bl_0_459 
* INOUT : br_0_459 
* INOUT : bl_0_460 
* INOUT : br_0_460 
* INOUT : bl_0_461 
* INOUT : br_0_461 
* INOUT : bl_0_462 
* INOUT : br_0_462 
* INOUT : bl_0_463 
* INOUT : br_0_463 
* INOUT : bl_0_464 
* INOUT : br_0_464 
* INOUT : bl_0_465 
* INOUT : br_0_465 
* INOUT : bl_0_466 
* INOUT : br_0_466 
* INOUT : bl_0_467 
* INOUT : br_0_467 
* INOUT : bl_0_468 
* INOUT : br_0_468 
* INOUT : bl_0_469 
* INOUT : br_0_469 
* INOUT : bl_0_470 
* INOUT : br_0_470 
* INOUT : bl_0_471 
* INOUT : br_0_471 
* INOUT : bl_0_472 
* INOUT : br_0_472 
* INOUT : bl_0_473 
* INOUT : br_0_473 
* INOUT : bl_0_474 
* INOUT : br_0_474 
* INOUT : bl_0_475 
* INOUT : br_0_475 
* INOUT : bl_0_476 
* INOUT : br_0_476 
* INOUT : bl_0_477 
* INOUT : br_0_477 
* INOUT : bl_0_478 
* INOUT : br_0_478 
* INOUT : bl_0_479 
* INOUT : br_0_479 
* INOUT : bl_0_480 
* INOUT : br_0_480 
* INOUT : bl_0_481 
* INOUT : br_0_481 
* INOUT : bl_0_482 
* INOUT : br_0_482 
* INOUT : bl_0_483 
* INOUT : br_0_483 
* INOUT : bl_0_484 
* INOUT : br_0_484 
* INOUT : bl_0_485 
* INOUT : br_0_485 
* INOUT : bl_0_486 
* INOUT : br_0_486 
* INOUT : bl_0_487 
* INOUT : br_0_487 
* INOUT : bl_0_488 
* INOUT : br_0_488 
* INOUT : bl_0_489 
* INOUT : br_0_489 
* INOUT : bl_0_490 
* INOUT : br_0_490 
* INOUT : bl_0_491 
* INOUT : br_0_491 
* INOUT : bl_0_492 
* INOUT : br_0_492 
* INOUT : bl_0_493 
* INOUT : br_0_493 
* INOUT : bl_0_494 
* INOUT : br_0_494 
* INOUT : bl_0_495 
* INOUT : br_0_495 
* INOUT : bl_0_496 
* INOUT : br_0_496 
* INOUT : bl_0_497 
* INOUT : br_0_497 
* INOUT : bl_0_498 
* INOUT : br_0_498 
* INOUT : bl_0_499 
* INOUT : br_0_499 
* INOUT : bl_0_500 
* INOUT : br_0_500 
* INOUT : bl_0_501 
* INOUT : br_0_501 
* INOUT : bl_0_502 
* INOUT : br_0_502 
* INOUT : bl_0_503 
* INOUT : br_0_503 
* INOUT : bl_0_504 
* INOUT : br_0_504 
* INOUT : bl_0_505 
* INOUT : br_0_505 
* INOUT : bl_0_506 
* INOUT : br_0_506 
* INOUT : bl_0_507 
* INOUT : br_0_507 
* INOUT : bl_0_508 
* INOUT : br_0_508 
* INOUT : bl_0_509 
* INOUT : br_0_509 
* INOUT : bl_0_510 
* INOUT : br_0_510 
* INOUT : bl_0_511 
* INOUT : br_0_511 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c256
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c257
+ bl_0_257 br_0_257 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c258
+ bl_0_258 br_0_258 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c259
+ bl_0_259 br_0_259 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c260
+ bl_0_260 br_0_260 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c261
+ bl_0_261 br_0_261 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c262
+ bl_0_262 br_0_262 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c263
+ bl_0_263 br_0_263 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c264
+ bl_0_264 br_0_264 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c265
+ bl_0_265 br_0_265 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c266
+ bl_0_266 br_0_266 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c267
+ bl_0_267 br_0_267 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c268
+ bl_0_268 br_0_268 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c269
+ bl_0_269 br_0_269 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c270
+ bl_0_270 br_0_270 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c271
+ bl_0_271 br_0_271 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c272
+ bl_0_272 br_0_272 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c273
+ bl_0_273 br_0_273 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c274
+ bl_0_274 br_0_274 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c275
+ bl_0_275 br_0_275 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c276
+ bl_0_276 br_0_276 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c277
+ bl_0_277 br_0_277 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c278
+ bl_0_278 br_0_278 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c279
+ bl_0_279 br_0_279 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c280
+ bl_0_280 br_0_280 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c281
+ bl_0_281 br_0_281 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c282
+ bl_0_282 br_0_282 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c283
+ bl_0_283 br_0_283 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c284
+ bl_0_284 br_0_284 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c285
+ bl_0_285 br_0_285 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c286
+ bl_0_286 br_0_286 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c287
+ bl_0_287 br_0_287 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c288
+ bl_0_288 br_0_288 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c289
+ bl_0_289 br_0_289 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c290
+ bl_0_290 br_0_290 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c291
+ bl_0_291 br_0_291 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c292
+ bl_0_292 br_0_292 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c293
+ bl_0_293 br_0_293 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c294
+ bl_0_294 br_0_294 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c295
+ bl_0_295 br_0_295 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c296
+ bl_0_296 br_0_296 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c297
+ bl_0_297 br_0_297 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c298
+ bl_0_298 br_0_298 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c299
+ bl_0_299 br_0_299 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c300
+ bl_0_300 br_0_300 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c301
+ bl_0_301 br_0_301 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c302
+ bl_0_302 br_0_302 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c303
+ bl_0_303 br_0_303 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c304
+ bl_0_304 br_0_304 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c305
+ bl_0_305 br_0_305 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c306
+ bl_0_306 br_0_306 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c307
+ bl_0_307 br_0_307 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c308
+ bl_0_308 br_0_308 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c309
+ bl_0_309 br_0_309 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c310
+ bl_0_310 br_0_310 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c311
+ bl_0_311 br_0_311 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c312
+ bl_0_312 br_0_312 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c313
+ bl_0_313 br_0_313 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c314
+ bl_0_314 br_0_314 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c315
+ bl_0_315 br_0_315 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c316
+ bl_0_316 br_0_316 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c317
+ bl_0_317 br_0_317 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c318
+ bl_0_318 br_0_318 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c319
+ bl_0_319 br_0_319 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c320
+ bl_0_320 br_0_320 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c321
+ bl_0_321 br_0_321 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c322
+ bl_0_322 br_0_322 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c323
+ bl_0_323 br_0_323 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c324
+ bl_0_324 br_0_324 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c325
+ bl_0_325 br_0_325 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c326
+ bl_0_326 br_0_326 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c327
+ bl_0_327 br_0_327 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c328
+ bl_0_328 br_0_328 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c329
+ bl_0_329 br_0_329 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c330
+ bl_0_330 br_0_330 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c331
+ bl_0_331 br_0_331 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c332
+ bl_0_332 br_0_332 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c333
+ bl_0_333 br_0_333 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c334
+ bl_0_334 br_0_334 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c335
+ bl_0_335 br_0_335 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c336
+ bl_0_336 br_0_336 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c337
+ bl_0_337 br_0_337 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c338
+ bl_0_338 br_0_338 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c339
+ bl_0_339 br_0_339 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c340
+ bl_0_340 br_0_340 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c341
+ bl_0_341 br_0_341 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c342
+ bl_0_342 br_0_342 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c343
+ bl_0_343 br_0_343 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c344
+ bl_0_344 br_0_344 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c345
+ bl_0_345 br_0_345 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c346
+ bl_0_346 br_0_346 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c347
+ bl_0_347 br_0_347 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c348
+ bl_0_348 br_0_348 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c349
+ bl_0_349 br_0_349 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c350
+ bl_0_350 br_0_350 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c351
+ bl_0_351 br_0_351 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c352
+ bl_0_352 br_0_352 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c353
+ bl_0_353 br_0_353 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c354
+ bl_0_354 br_0_354 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c355
+ bl_0_355 br_0_355 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c356
+ bl_0_356 br_0_356 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c357
+ bl_0_357 br_0_357 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c358
+ bl_0_358 br_0_358 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c359
+ bl_0_359 br_0_359 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c360
+ bl_0_360 br_0_360 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c361
+ bl_0_361 br_0_361 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c362
+ bl_0_362 br_0_362 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c363
+ bl_0_363 br_0_363 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c364
+ bl_0_364 br_0_364 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c365
+ bl_0_365 br_0_365 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c366
+ bl_0_366 br_0_366 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c367
+ bl_0_367 br_0_367 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c368
+ bl_0_368 br_0_368 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c369
+ bl_0_369 br_0_369 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c370
+ bl_0_370 br_0_370 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c371
+ bl_0_371 br_0_371 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c372
+ bl_0_372 br_0_372 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c373
+ bl_0_373 br_0_373 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c374
+ bl_0_374 br_0_374 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c375
+ bl_0_375 br_0_375 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c376
+ bl_0_376 br_0_376 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c377
+ bl_0_377 br_0_377 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c378
+ bl_0_378 br_0_378 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c379
+ bl_0_379 br_0_379 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c380
+ bl_0_380 br_0_380 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c381
+ bl_0_381 br_0_381 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c382
+ bl_0_382 br_0_382 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c383
+ bl_0_383 br_0_383 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c384
+ bl_0_384 br_0_384 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c385
+ bl_0_385 br_0_385 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c386
+ bl_0_386 br_0_386 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c387
+ bl_0_387 br_0_387 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c388
+ bl_0_388 br_0_388 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c389
+ bl_0_389 br_0_389 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c390
+ bl_0_390 br_0_390 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c391
+ bl_0_391 br_0_391 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c392
+ bl_0_392 br_0_392 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c393
+ bl_0_393 br_0_393 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c394
+ bl_0_394 br_0_394 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c395
+ bl_0_395 br_0_395 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c396
+ bl_0_396 br_0_396 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c397
+ bl_0_397 br_0_397 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c398
+ bl_0_398 br_0_398 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c399
+ bl_0_399 br_0_399 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c400
+ bl_0_400 br_0_400 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c401
+ bl_0_401 br_0_401 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c402
+ bl_0_402 br_0_402 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c403
+ bl_0_403 br_0_403 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c404
+ bl_0_404 br_0_404 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c405
+ bl_0_405 br_0_405 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c406
+ bl_0_406 br_0_406 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c407
+ bl_0_407 br_0_407 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c408
+ bl_0_408 br_0_408 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c409
+ bl_0_409 br_0_409 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c410
+ bl_0_410 br_0_410 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c411
+ bl_0_411 br_0_411 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c412
+ bl_0_412 br_0_412 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c413
+ bl_0_413 br_0_413 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c414
+ bl_0_414 br_0_414 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c415
+ bl_0_415 br_0_415 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c416
+ bl_0_416 br_0_416 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c417
+ bl_0_417 br_0_417 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c418
+ bl_0_418 br_0_418 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c419
+ bl_0_419 br_0_419 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c420
+ bl_0_420 br_0_420 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c421
+ bl_0_421 br_0_421 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c422
+ bl_0_422 br_0_422 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c423
+ bl_0_423 br_0_423 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c424
+ bl_0_424 br_0_424 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c425
+ bl_0_425 br_0_425 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c426
+ bl_0_426 br_0_426 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c427
+ bl_0_427 br_0_427 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c428
+ bl_0_428 br_0_428 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c429
+ bl_0_429 br_0_429 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c430
+ bl_0_430 br_0_430 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c431
+ bl_0_431 br_0_431 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c432
+ bl_0_432 br_0_432 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c433
+ bl_0_433 br_0_433 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c434
+ bl_0_434 br_0_434 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c435
+ bl_0_435 br_0_435 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c436
+ bl_0_436 br_0_436 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c437
+ bl_0_437 br_0_437 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c438
+ bl_0_438 br_0_438 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c439
+ bl_0_439 br_0_439 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c440
+ bl_0_440 br_0_440 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c441
+ bl_0_441 br_0_441 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c442
+ bl_0_442 br_0_442 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c443
+ bl_0_443 br_0_443 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c444
+ bl_0_444 br_0_444 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c445
+ bl_0_445 br_0_445 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c446
+ bl_0_446 br_0_446 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c447
+ bl_0_447 br_0_447 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c448
+ bl_0_448 br_0_448 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c449
+ bl_0_449 br_0_449 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c450
+ bl_0_450 br_0_450 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c451
+ bl_0_451 br_0_451 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c452
+ bl_0_452 br_0_452 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c453
+ bl_0_453 br_0_453 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c454
+ bl_0_454 br_0_454 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c455
+ bl_0_455 br_0_455 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c456
+ bl_0_456 br_0_456 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c457
+ bl_0_457 br_0_457 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c458
+ bl_0_458 br_0_458 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c459
+ bl_0_459 br_0_459 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c460
+ bl_0_460 br_0_460 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c461
+ bl_0_461 br_0_461 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c462
+ bl_0_462 br_0_462 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c463
+ bl_0_463 br_0_463 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c464
+ bl_0_464 br_0_464 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c465
+ bl_0_465 br_0_465 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c466
+ bl_0_466 br_0_466 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c467
+ bl_0_467 br_0_467 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c468
+ bl_0_468 br_0_468 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c469
+ bl_0_469 br_0_469 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c470
+ bl_0_470 br_0_470 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c471
+ bl_0_471 br_0_471 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c472
+ bl_0_472 br_0_472 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c473
+ bl_0_473 br_0_473 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c474
+ bl_0_474 br_0_474 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c475
+ bl_0_475 br_0_475 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c476
+ bl_0_476 br_0_476 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c477
+ bl_0_477 br_0_477 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c478
+ bl_0_478 br_0_478 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c479
+ bl_0_479 br_0_479 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c480
+ bl_0_480 br_0_480 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c481
+ bl_0_481 br_0_481 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c482
+ bl_0_482 br_0_482 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c483
+ bl_0_483 br_0_483 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c484
+ bl_0_484 br_0_484 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c485
+ bl_0_485 br_0_485 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c486
+ bl_0_486 br_0_486 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c487
+ bl_0_487 br_0_487 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c488
+ bl_0_488 br_0_488 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c489
+ bl_0_489 br_0_489 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c490
+ bl_0_490 br_0_490 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c491
+ bl_0_491 br_0_491 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c492
+ bl_0_492 br_0_492 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c493
+ bl_0_493 br_0_493 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c494
+ bl_0_494 br_0_494 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c495
+ bl_0_495 br_0_495 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c496
+ bl_0_496 br_0_496 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c497
+ bl_0_497 br_0_497 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c498
+ bl_0_498 br_0_498 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c499
+ bl_0_499 br_0_499 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c500
+ bl_0_500 br_0_500 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c501
+ bl_0_501 br_0_501 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c502
+ bl_0_502 br_0_502 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c503
+ bl_0_503 br_0_503 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c504
+ bl_0_504 br_0_504 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c505
+ bl_0_505 br_0_505 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c506
+ bl_0_506 br_0_506 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c507
+ bl_0_507 br_0_507 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c508
+ bl_0_508 br_0_508 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c509
+ bl_0_509 br_0_509 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c510
+ bl_0_510 br_0_510 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c511
+ bl_0_511 br_0_511 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS freepdk45_sram_1rw0r_45x512_dummy_array

.SUBCKT freepdk45_sram_1rw0r_45x512_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258
+ br_0_258 bl_0_259 br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261
+ bl_0_262 br_0_262 bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265
+ br_0_265 bl_0_266 br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268
+ bl_0_269 br_0_269 bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272
+ br_0_272 bl_0_273 br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275
+ bl_0_276 br_0_276 bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279
+ br_0_279 bl_0_280 br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282
+ bl_0_283 br_0_283 bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286
+ br_0_286 bl_0_287 br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289
+ bl_0_290 br_0_290 bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293
+ br_0_293 bl_0_294 br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296
+ bl_0_297 br_0_297 bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300
+ br_0_300 bl_0_301 br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303
+ bl_0_304 br_0_304 bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307
+ br_0_307 bl_0_308 br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310
+ bl_0_311 br_0_311 bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314
+ br_0_314 bl_0_315 br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317
+ bl_0_318 br_0_318 bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321
+ br_0_321 bl_0_322 br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324
+ bl_0_325 br_0_325 bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328
+ br_0_328 bl_0_329 br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331
+ bl_0_332 br_0_332 bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335
+ br_0_335 bl_0_336 br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338
+ bl_0_339 br_0_339 bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342
+ br_0_342 bl_0_343 br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345
+ bl_0_346 br_0_346 bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349
+ br_0_349 bl_0_350 br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352
+ bl_0_353 br_0_353 bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356
+ br_0_356 bl_0_357 br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359
+ bl_0_360 br_0_360 bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363
+ br_0_363 bl_0_364 br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366
+ bl_0_367 br_0_367 bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370
+ br_0_370 bl_0_371 br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373
+ bl_0_374 br_0_374 bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377
+ br_0_377 bl_0_378 br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380
+ bl_0_381 br_0_381 bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384
+ br_0_384 bl_0_385 br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387
+ bl_0_388 br_0_388 bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391
+ br_0_391 bl_0_392 br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394
+ bl_0_395 br_0_395 bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398
+ br_0_398 bl_0_399 br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401
+ bl_0_402 br_0_402 bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405
+ br_0_405 bl_0_406 br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408
+ bl_0_409 br_0_409 bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412
+ br_0_412 bl_0_413 br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415
+ bl_0_416 br_0_416 bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419
+ br_0_419 bl_0_420 br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422
+ bl_0_423 br_0_423 bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426
+ br_0_426 bl_0_427 br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429
+ bl_0_430 br_0_430 bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433
+ br_0_433 bl_0_434 br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436
+ bl_0_437 br_0_437 bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440
+ br_0_440 bl_0_441 br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443
+ bl_0_444 br_0_444 bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447
+ br_0_447 bl_0_448 br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450
+ bl_0_451 br_0_451 bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454
+ br_0_454 bl_0_455 br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457
+ bl_0_458 br_0_458 bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461
+ br_0_461 bl_0_462 br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464
+ bl_0_465 br_0_465 bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468
+ br_0_468 bl_0_469 br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471
+ bl_0_472 br_0_472 bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475
+ br_0_475 bl_0_476 br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478
+ bl_0_479 br_0_479 bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482
+ br_0_482 bl_0_483 br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485
+ bl_0_486 br_0_486 bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489
+ br_0_489 bl_0_490 br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492
+ bl_0_493 br_0_493 bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496
+ br_0_496 bl_0_497 br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499
+ bl_0_500 br_0_500 bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503
+ br_0_503 bl_0_504 br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506
+ bl_0_507 br_0_507 bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510
+ br_0_510 bl_0_511 br_0_511 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3
+ wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12
+ wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20
+ wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28
+ wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36
+ wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 vdd
+ gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INOUT : bl_0_257 
* INOUT : br_0_257 
* INOUT : bl_0_258 
* INOUT : br_0_258 
* INOUT : bl_0_259 
* INOUT : br_0_259 
* INOUT : bl_0_260 
* INOUT : br_0_260 
* INOUT : bl_0_261 
* INOUT : br_0_261 
* INOUT : bl_0_262 
* INOUT : br_0_262 
* INOUT : bl_0_263 
* INOUT : br_0_263 
* INOUT : bl_0_264 
* INOUT : br_0_264 
* INOUT : bl_0_265 
* INOUT : br_0_265 
* INOUT : bl_0_266 
* INOUT : br_0_266 
* INOUT : bl_0_267 
* INOUT : br_0_267 
* INOUT : bl_0_268 
* INOUT : br_0_268 
* INOUT : bl_0_269 
* INOUT : br_0_269 
* INOUT : bl_0_270 
* INOUT : br_0_270 
* INOUT : bl_0_271 
* INOUT : br_0_271 
* INOUT : bl_0_272 
* INOUT : br_0_272 
* INOUT : bl_0_273 
* INOUT : br_0_273 
* INOUT : bl_0_274 
* INOUT : br_0_274 
* INOUT : bl_0_275 
* INOUT : br_0_275 
* INOUT : bl_0_276 
* INOUT : br_0_276 
* INOUT : bl_0_277 
* INOUT : br_0_277 
* INOUT : bl_0_278 
* INOUT : br_0_278 
* INOUT : bl_0_279 
* INOUT : br_0_279 
* INOUT : bl_0_280 
* INOUT : br_0_280 
* INOUT : bl_0_281 
* INOUT : br_0_281 
* INOUT : bl_0_282 
* INOUT : br_0_282 
* INOUT : bl_0_283 
* INOUT : br_0_283 
* INOUT : bl_0_284 
* INOUT : br_0_284 
* INOUT : bl_0_285 
* INOUT : br_0_285 
* INOUT : bl_0_286 
* INOUT : br_0_286 
* INOUT : bl_0_287 
* INOUT : br_0_287 
* INOUT : bl_0_288 
* INOUT : br_0_288 
* INOUT : bl_0_289 
* INOUT : br_0_289 
* INOUT : bl_0_290 
* INOUT : br_0_290 
* INOUT : bl_0_291 
* INOUT : br_0_291 
* INOUT : bl_0_292 
* INOUT : br_0_292 
* INOUT : bl_0_293 
* INOUT : br_0_293 
* INOUT : bl_0_294 
* INOUT : br_0_294 
* INOUT : bl_0_295 
* INOUT : br_0_295 
* INOUT : bl_0_296 
* INOUT : br_0_296 
* INOUT : bl_0_297 
* INOUT : br_0_297 
* INOUT : bl_0_298 
* INOUT : br_0_298 
* INOUT : bl_0_299 
* INOUT : br_0_299 
* INOUT : bl_0_300 
* INOUT : br_0_300 
* INOUT : bl_0_301 
* INOUT : br_0_301 
* INOUT : bl_0_302 
* INOUT : br_0_302 
* INOUT : bl_0_303 
* INOUT : br_0_303 
* INOUT : bl_0_304 
* INOUT : br_0_304 
* INOUT : bl_0_305 
* INOUT : br_0_305 
* INOUT : bl_0_306 
* INOUT : br_0_306 
* INOUT : bl_0_307 
* INOUT : br_0_307 
* INOUT : bl_0_308 
* INOUT : br_0_308 
* INOUT : bl_0_309 
* INOUT : br_0_309 
* INOUT : bl_0_310 
* INOUT : br_0_310 
* INOUT : bl_0_311 
* INOUT : br_0_311 
* INOUT : bl_0_312 
* INOUT : br_0_312 
* INOUT : bl_0_313 
* INOUT : br_0_313 
* INOUT : bl_0_314 
* INOUT : br_0_314 
* INOUT : bl_0_315 
* INOUT : br_0_315 
* INOUT : bl_0_316 
* INOUT : br_0_316 
* INOUT : bl_0_317 
* INOUT : br_0_317 
* INOUT : bl_0_318 
* INOUT : br_0_318 
* INOUT : bl_0_319 
* INOUT : br_0_319 
* INOUT : bl_0_320 
* INOUT : br_0_320 
* INOUT : bl_0_321 
* INOUT : br_0_321 
* INOUT : bl_0_322 
* INOUT : br_0_322 
* INOUT : bl_0_323 
* INOUT : br_0_323 
* INOUT : bl_0_324 
* INOUT : br_0_324 
* INOUT : bl_0_325 
* INOUT : br_0_325 
* INOUT : bl_0_326 
* INOUT : br_0_326 
* INOUT : bl_0_327 
* INOUT : br_0_327 
* INOUT : bl_0_328 
* INOUT : br_0_328 
* INOUT : bl_0_329 
* INOUT : br_0_329 
* INOUT : bl_0_330 
* INOUT : br_0_330 
* INOUT : bl_0_331 
* INOUT : br_0_331 
* INOUT : bl_0_332 
* INOUT : br_0_332 
* INOUT : bl_0_333 
* INOUT : br_0_333 
* INOUT : bl_0_334 
* INOUT : br_0_334 
* INOUT : bl_0_335 
* INOUT : br_0_335 
* INOUT : bl_0_336 
* INOUT : br_0_336 
* INOUT : bl_0_337 
* INOUT : br_0_337 
* INOUT : bl_0_338 
* INOUT : br_0_338 
* INOUT : bl_0_339 
* INOUT : br_0_339 
* INOUT : bl_0_340 
* INOUT : br_0_340 
* INOUT : bl_0_341 
* INOUT : br_0_341 
* INOUT : bl_0_342 
* INOUT : br_0_342 
* INOUT : bl_0_343 
* INOUT : br_0_343 
* INOUT : bl_0_344 
* INOUT : br_0_344 
* INOUT : bl_0_345 
* INOUT : br_0_345 
* INOUT : bl_0_346 
* INOUT : br_0_346 
* INOUT : bl_0_347 
* INOUT : br_0_347 
* INOUT : bl_0_348 
* INOUT : br_0_348 
* INOUT : bl_0_349 
* INOUT : br_0_349 
* INOUT : bl_0_350 
* INOUT : br_0_350 
* INOUT : bl_0_351 
* INOUT : br_0_351 
* INOUT : bl_0_352 
* INOUT : br_0_352 
* INOUT : bl_0_353 
* INOUT : br_0_353 
* INOUT : bl_0_354 
* INOUT : br_0_354 
* INOUT : bl_0_355 
* INOUT : br_0_355 
* INOUT : bl_0_356 
* INOUT : br_0_356 
* INOUT : bl_0_357 
* INOUT : br_0_357 
* INOUT : bl_0_358 
* INOUT : br_0_358 
* INOUT : bl_0_359 
* INOUT : br_0_359 
* INOUT : bl_0_360 
* INOUT : br_0_360 
* INOUT : bl_0_361 
* INOUT : br_0_361 
* INOUT : bl_0_362 
* INOUT : br_0_362 
* INOUT : bl_0_363 
* INOUT : br_0_363 
* INOUT : bl_0_364 
* INOUT : br_0_364 
* INOUT : bl_0_365 
* INOUT : br_0_365 
* INOUT : bl_0_366 
* INOUT : br_0_366 
* INOUT : bl_0_367 
* INOUT : br_0_367 
* INOUT : bl_0_368 
* INOUT : br_0_368 
* INOUT : bl_0_369 
* INOUT : br_0_369 
* INOUT : bl_0_370 
* INOUT : br_0_370 
* INOUT : bl_0_371 
* INOUT : br_0_371 
* INOUT : bl_0_372 
* INOUT : br_0_372 
* INOUT : bl_0_373 
* INOUT : br_0_373 
* INOUT : bl_0_374 
* INOUT : br_0_374 
* INOUT : bl_0_375 
* INOUT : br_0_375 
* INOUT : bl_0_376 
* INOUT : br_0_376 
* INOUT : bl_0_377 
* INOUT : br_0_377 
* INOUT : bl_0_378 
* INOUT : br_0_378 
* INOUT : bl_0_379 
* INOUT : br_0_379 
* INOUT : bl_0_380 
* INOUT : br_0_380 
* INOUT : bl_0_381 
* INOUT : br_0_381 
* INOUT : bl_0_382 
* INOUT : br_0_382 
* INOUT : bl_0_383 
* INOUT : br_0_383 
* INOUT : bl_0_384 
* INOUT : br_0_384 
* INOUT : bl_0_385 
* INOUT : br_0_385 
* INOUT : bl_0_386 
* INOUT : br_0_386 
* INOUT : bl_0_387 
* INOUT : br_0_387 
* INOUT : bl_0_388 
* INOUT : br_0_388 
* INOUT : bl_0_389 
* INOUT : br_0_389 
* INOUT : bl_0_390 
* INOUT : br_0_390 
* INOUT : bl_0_391 
* INOUT : br_0_391 
* INOUT : bl_0_392 
* INOUT : br_0_392 
* INOUT : bl_0_393 
* INOUT : br_0_393 
* INOUT : bl_0_394 
* INOUT : br_0_394 
* INOUT : bl_0_395 
* INOUT : br_0_395 
* INOUT : bl_0_396 
* INOUT : br_0_396 
* INOUT : bl_0_397 
* INOUT : br_0_397 
* INOUT : bl_0_398 
* INOUT : br_0_398 
* INOUT : bl_0_399 
* INOUT : br_0_399 
* INOUT : bl_0_400 
* INOUT : br_0_400 
* INOUT : bl_0_401 
* INOUT : br_0_401 
* INOUT : bl_0_402 
* INOUT : br_0_402 
* INOUT : bl_0_403 
* INOUT : br_0_403 
* INOUT : bl_0_404 
* INOUT : br_0_404 
* INOUT : bl_0_405 
* INOUT : br_0_405 
* INOUT : bl_0_406 
* INOUT : br_0_406 
* INOUT : bl_0_407 
* INOUT : br_0_407 
* INOUT : bl_0_408 
* INOUT : br_0_408 
* INOUT : bl_0_409 
* INOUT : br_0_409 
* INOUT : bl_0_410 
* INOUT : br_0_410 
* INOUT : bl_0_411 
* INOUT : br_0_411 
* INOUT : bl_0_412 
* INOUT : br_0_412 
* INOUT : bl_0_413 
* INOUT : br_0_413 
* INOUT : bl_0_414 
* INOUT : br_0_414 
* INOUT : bl_0_415 
* INOUT : br_0_415 
* INOUT : bl_0_416 
* INOUT : br_0_416 
* INOUT : bl_0_417 
* INOUT : br_0_417 
* INOUT : bl_0_418 
* INOUT : br_0_418 
* INOUT : bl_0_419 
* INOUT : br_0_419 
* INOUT : bl_0_420 
* INOUT : br_0_420 
* INOUT : bl_0_421 
* INOUT : br_0_421 
* INOUT : bl_0_422 
* INOUT : br_0_422 
* INOUT : bl_0_423 
* INOUT : br_0_423 
* INOUT : bl_0_424 
* INOUT : br_0_424 
* INOUT : bl_0_425 
* INOUT : br_0_425 
* INOUT : bl_0_426 
* INOUT : br_0_426 
* INOUT : bl_0_427 
* INOUT : br_0_427 
* INOUT : bl_0_428 
* INOUT : br_0_428 
* INOUT : bl_0_429 
* INOUT : br_0_429 
* INOUT : bl_0_430 
* INOUT : br_0_430 
* INOUT : bl_0_431 
* INOUT : br_0_431 
* INOUT : bl_0_432 
* INOUT : br_0_432 
* INOUT : bl_0_433 
* INOUT : br_0_433 
* INOUT : bl_0_434 
* INOUT : br_0_434 
* INOUT : bl_0_435 
* INOUT : br_0_435 
* INOUT : bl_0_436 
* INOUT : br_0_436 
* INOUT : bl_0_437 
* INOUT : br_0_437 
* INOUT : bl_0_438 
* INOUT : br_0_438 
* INOUT : bl_0_439 
* INOUT : br_0_439 
* INOUT : bl_0_440 
* INOUT : br_0_440 
* INOUT : bl_0_441 
* INOUT : br_0_441 
* INOUT : bl_0_442 
* INOUT : br_0_442 
* INOUT : bl_0_443 
* INOUT : br_0_443 
* INOUT : bl_0_444 
* INOUT : br_0_444 
* INOUT : bl_0_445 
* INOUT : br_0_445 
* INOUT : bl_0_446 
* INOUT : br_0_446 
* INOUT : bl_0_447 
* INOUT : br_0_447 
* INOUT : bl_0_448 
* INOUT : br_0_448 
* INOUT : bl_0_449 
* INOUT : br_0_449 
* INOUT : bl_0_450 
* INOUT : br_0_450 
* INOUT : bl_0_451 
* INOUT : br_0_451 
* INOUT : bl_0_452 
* INOUT : br_0_452 
* INOUT : bl_0_453 
* INOUT : br_0_453 
* INOUT : bl_0_454 
* INOUT : br_0_454 
* INOUT : bl_0_455 
* INOUT : br_0_455 
* INOUT : bl_0_456 
* INOUT : br_0_456 
* INOUT : bl_0_457 
* INOUT : br_0_457 
* INOUT : bl_0_458 
* INOUT : br_0_458 
* INOUT : bl_0_459 
* INOUT : br_0_459 
* INOUT : bl_0_460 
* INOUT : br_0_460 
* INOUT : bl_0_461 
* INOUT : br_0_461 
* INOUT : bl_0_462 
* INOUT : br_0_462 
* INOUT : bl_0_463 
* INOUT : br_0_463 
* INOUT : bl_0_464 
* INOUT : br_0_464 
* INOUT : bl_0_465 
* INOUT : br_0_465 
* INOUT : bl_0_466 
* INOUT : br_0_466 
* INOUT : bl_0_467 
* INOUT : br_0_467 
* INOUT : bl_0_468 
* INOUT : br_0_468 
* INOUT : bl_0_469 
* INOUT : br_0_469 
* INOUT : bl_0_470 
* INOUT : br_0_470 
* INOUT : bl_0_471 
* INOUT : br_0_471 
* INOUT : bl_0_472 
* INOUT : br_0_472 
* INOUT : bl_0_473 
* INOUT : br_0_473 
* INOUT : bl_0_474 
* INOUT : br_0_474 
* INOUT : bl_0_475 
* INOUT : br_0_475 
* INOUT : bl_0_476 
* INOUT : br_0_476 
* INOUT : bl_0_477 
* INOUT : br_0_477 
* INOUT : bl_0_478 
* INOUT : br_0_478 
* INOUT : bl_0_479 
* INOUT : br_0_479 
* INOUT : bl_0_480 
* INOUT : br_0_480 
* INOUT : bl_0_481 
* INOUT : br_0_481 
* INOUT : bl_0_482 
* INOUT : br_0_482 
* INOUT : bl_0_483 
* INOUT : br_0_483 
* INOUT : bl_0_484 
* INOUT : br_0_484 
* INOUT : bl_0_485 
* INOUT : br_0_485 
* INOUT : bl_0_486 
* INOUT : br_0_486 
* INOUT : bl_0_487 
* INOUT : br_0_487 
* INOUT : bl_0_488 
* INOUT : br_0_488 
* INOUT : bl_0_489 
* INOUT : br_0_489 
* INOUT : bl_0_490 
* INOUT : br_0_490 
* INOUT : bl_0_491 
* INOUT : br_0_491 
* INOUT : bl_0_492 
* INOUT : br_0_492 
* INOUT : bl_0_493 
* INOUT : br_0_493 
* INOUT : bl_0_494 
* INOUT : br_0_494 
* INOUT : bl_0_495 
* INOUT : br_0_495 
* INOUT : bl_0_496 
* INOUT : br_0_496 
* INOUT : bl_0_497 
* INOUT : br_0_497 
* INOUT : bl_0_498 
* INOUT : br_0_498 
* INOUT : bl_0_499 
* INOUT : br_0_499 
* INOUT : bl_0_500 
* INOUT : br_0_500 
* INOUT : bl_0_501 
* INOUT : br_0_501 
* INOUT : bl_0_502 
* INOUT : br_0_502 
* INOUT : bl_0_503 
* INOUT : br_0_503 
* INOUT : bl_0_504 
* INOUT : br_0_504 
* INOUT : bl_0_505 
* INOUT : br_0_505 
* INOUT : bl_0_506 
* INOUT : br_0_506 
* INOUT : bl_0_507 
* INOUT : br_0_507 
* INOUT : bl_0_508 
* INOUT : br_0_508 
* INOUT : bl_0_509 
* INOUT : br_0_509 
* INOUT : bl_0_510 
* INOUT : br_0_510 
* INOUT : bl_0_511 
* INOUT : br_0_511 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* POWER : vdd 
* GROUND: gnd 
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xbitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258 br_0_258 bl_0_259
+ br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261 bl_0_262 br_0_262
+ bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265 br_0_265 bl_0_266
+ br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268 bl_0_269 br_0_269
+ bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272 br_0_272 bl_0_273
+ br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275 bl_0_276 br_0_276
+ bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279 br_0_279 bl_0_280
+ br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282 bl_0_283 br_0_283
+ bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286 br_0_286 bl_0_287
+ br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289 bl_0_290 br_0_290
+ bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293 br_0_293 bl_0_294
+ br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296 bl_0_297 br_0_297
+ bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300 br_0_300 bl_0_301
+ br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303 bl_0_304 br_0_304
+ bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307 br_0_307 bl_0_308
+ br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310 bl_0_311 br_0_311
+ bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314 br_0_314 bl_0_315
+ br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317 bl_0_318 br_0_318
+ bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321 br_0_321 bl_0_322
+ br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324 bl_0_325 br_0_325
+ bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328 br_0_328 bl_0_329
+ br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331 bl_0_332 br_0_332
+ bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335 br_0_335 bl_0_336
+ br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338 bl_0_339 br_0_339
+ bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342 br_0_342 bl_0_343
+ br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345 bl_0_346 br_0_346
+ bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349 br_0_349 bl_0_350
+ br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352 bl_0_353 br_0_353
+ bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356 br_0_356 bl_0_357
+ br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359 bl_0_360 br_0_360
+ bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363 br_0_363 bl_0_364
+ br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366 bl_0_367 br_0_367
+ bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370 br_0_370 bl_0_371
+ br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373 bl_0_374 br_0_374
+ bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377 br_0_377 bl_0_378
+ br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380 bl_0_381 br_0_381
+ bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384 br_0_384 bl_0_385
+ br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387 bl_0_388 br_0_388
+ bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391 br_0_391 bl_0_392
+ br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394 bl_0_395 br_0_395
+ bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398 br_0_398 bl_0_399
+ br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401 bl_0_402 br_0_402
+ bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405 br_0_405 bl_0_406
+ br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408 bl_0_409 br_0_409
+ bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412 br_0_412 bl_0_413
+ br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415 bl_0_416 br_0_416
+ bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419 br_0_419 bl_0_420
+ br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422 bl_0_423 br_0_423
+ bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426 br_0_426 bl_0_427
+ br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429 bl_0_430 br_0_430
+ bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433 br_0_433 bl_0_434
+ br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436 bl_0_437 br_0_437
+ bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440 br_0_440 bl_0_441
+ br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443 bl_0_444 br_0_444
+ bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447 br_0_447 bl_0_448
+ br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450 bl_0_451 br_0_451
+ bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454 br_0_454 bl_0_455
+ br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457 bl_0_458 br_0_458
+ bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461 br_0_461 bl_0_462
+ br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464 bl_0_465 br_0_465
+ bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468 br_0_468 bl_0_469
+ br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471 bl_0_472 br_0_472
+ bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475 br_0_475 bl_0_476
+ br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478 bl_0_479 br_0_479
+ bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482 br_0_482 bl_0_483
+ br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485 bl_0_486 br_0_486
+ bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489 br_0_489 bl_0_490
+ br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492 bl_0_493 br_0_493
+ bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496 br_0_496 bl_0_497
+ br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499 bl_0_500 br_0_500
+ bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503 br_0_503 bl_0_504
+ br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506 bl_0_507 br_0_507
+ bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510 br_0_510 bl_0_511
+ br_0_511 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 vdd gnd
+ freepdk45_sram_1rw0r_45x512_bitcell_array
Xreplica_col_0
+ rbl_bl_0_0 rbl_br_0_0 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4
+ wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13
+ wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21
+ wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37
+ wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 vdd gnd
+ freepdk45_sram_1rw0r_45x512_replica_column
Xdummy_row_0
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258 br_0_258 bl_0_259
+ br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261 bl_0_262 br_0_262
+ bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265 br_0_265 bl_0_266
+ br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268 bl_0_269 br_0_269
+ bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272 br_0_272 bl_0_273
+ br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275 bl_0_276 br_0_276
+ bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279 br_0_279 bl_0_280
+ br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282 bl_0_283 br_0_283
+ bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286 br_0_286 bl_0_287
+ br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289 bl_0_290 br_0_290
+ bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293 br_0_293 bl_0_294
+ br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296 bl_0_297 br_0_297
+ bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300 br_0_300 bl_0_301
+ br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303 bl_0_304 br_0_304
+ bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307 br_0_307 bl_0_308
+ br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310 bl_0_311 br_0_311
+ bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314 br_0_314 bl_0_315
+ br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317 bl_0_318 br_0_318
+ bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321 br_0_321 bl_0_322
+ br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324 bl_0_325 br_0_325
+ bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328 br_0_328 bl_0_329
+ br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331 bl_0_332 br_0_332
+ bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335 br_0_335 bl_0_336
+ br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338 bl_0_339 br_0_339
+ bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342 br_0_342 bl_0_343
+ br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345 bl_0_346 br_0_346
+ bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349 br_0_349 bl_0_350
+ br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352 bl_0_353 br_0_353
+ bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356 br_0_356 bl_0_357
+ br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359 bl_0_360 br_0_360
+ bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363 br_0_363 bl_0_364
+ br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366 bl_0_367 br_0_367
+ bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370 br_0_370 bl_0_371
+ br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373 bl_0_374 br_0_374
+ bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377 br_0_377 bl_0_378
+ br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380 bl_0_381 br_0_381
+ bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384 br_0_384 bl_0_385
+ br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387 bl_0_388 br_0_388
+ bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391 br_0_391 bl_0_392
+ br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394 bl_0_395 br_0_395
+ bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398 br_0_398 bl_0_399
+ br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401 bl_0_402 br_0_402
+ bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405 br_0_405 bl_0_406
+ br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408 bl_0_409 br_0_409
+ bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412 br_0_412 bl_0_413
+ br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415 bl_0_416 br_0_416
+ bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419 br_0_419 bl_0_420
+ br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422 bl_0_423 br_0_423
+ bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426 br_0_426 bl_0_427
+ br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429 bl_0_430 br_0_430
+ bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433 br_0_433 bl_0_434
+ br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436 bl_0_437 br_0_437
+ bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440 br_0_440 bl_0_441
+ br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443 bl_0_444 br_0_444
+ bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447 br_0_447 bl_0_448
+ br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450 bl_0_451 br_0_451
+ bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454 br_0_454 bl_0_455
+ br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457 bl_0_458 br_0_458
+ bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461 br_0_461 bl_0_462
+ br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464 bl_0_465 br_0_465
+ bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468 br_0_468 bl_0_469
+ br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471 bl_0_472 br_0_472
+ bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475 br_0_475 bl_0_476
+ br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478 bl_0_479 br_0_479
+ bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482 br_0_482 bl_0_483
+ br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485 bl_0_486 br_0_486
+ bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489 br_0_489 bl_0_490
+ br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492 bl_0_493 br_0_493
+ bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496 br_0_496 bl_0_497
+ br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499 bl_0_500 br_0_500
+ bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503 br_0_503 bl_0_504
+ br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506 bl_0_507 br_0_507
+ bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510 br_0_510 bl_0_511
+ br_0_511 rbl_wl_0_0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_dummy_array
.ENDS freepdk45_sram_1rw0r_45x512_replica_bitcell_array

.SUBCKT freepdk45_sram_1rw0r_45x512_dummy_array_2
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ dummy_cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ dummy_cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ dummy_cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ dummy_cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ dummy_cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ dummy_cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ dummy_cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ dummy_cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ dummy_cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ dummy_cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ dummy_cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ dummy_cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ dummy_cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ dummy_cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ dummy_cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ dummy_cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ dummy_cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ dummy_cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ dummy_cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ dummy_cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ dummy_cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ dummy_cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ dummy_cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ dummy_cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ dummy_cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ dummy_cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ dummy_cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ dummy_cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ dummy_cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ dummy_cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ dummy_cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ dummy_cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ dummy_cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ dummy_cell_1rw
Xbit_r35_c0
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ dummy_cell_1rw
Xbit_r36_c0
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ dummy_cell_1rw
Xbit_r37_c0
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ dummy_cell_1rw
Xbit_r38_c0
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ dummy_cell_1rw
Xbit_r39_c0
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ dummy_cell_1rw
Xbit_r40_c0
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ dummy_cell_1rw
Xbit_r41_c0
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ dummy_cell_1rw
Xbit_r42_c0
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ dummy_cell_1rw
Xbit_r43_c0
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ dummy_cell_1rw
Xbit_r44_c0
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ dummy_cell_1rw
Xbit_r45_c0
+ bl_0_0 br_0_0 wl_0_45 vdd gnd
+ dummy_cell_1rw
Xbit_r46_c0
+ bl_0_0 br_0_0 wl_0_46 vdd gnd
+ dummy_cell_1rw
Xbit_r47_c0
+ bl_0_0 br_0_0 wl_0_47 vdd gnd
+ dummy_cell_1rw
.ENDS freepdk45_sram_1rw0r_45x512_dummy_array_2

.SUBCKT freepdk45_sram_1rw0r_45x512_dummy_array_1
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258 br_0_258 bl_0_259
+ br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261 bl_0_262 br_0_262
+ bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265 br_0_265 bl_0_266
+ br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268 bl_0_269 br_0_269
+ bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272 br_0_272 bl_0_273
+ br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275 bl_0_276 br_0_276
+ bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279 br_0_279 bl_0_280
+ br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282 bl_0_283 br_0_283
+ bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286 br_0_286 bl_0_287
+ br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289 bl_0_290 br_0_290
+ bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293 br_0_293 bl_0_294
+ br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296 bl_0_297 br_0_297
+ bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300 br_0_300 bl_0_301
+ br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303 bl_0_304 br_0_304
+ bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307 br_0_307 bl_0_308
+ br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310 bl_0_311 br_0_311
+ bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314 br_0_314 bl_0_315
+ br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317 bl_0_318 br_0_318
+ bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321 br_0_321 bl_0_322
+ br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324 bl_0_325 br_0_325
+ bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328 br_0_328 bl_0_329
+ br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331 bl_0_332 br_0_332
+ bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335 br_0_335 bl_0_336
+ br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338 bl_0_339 br_0_339
+ bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342 br_0_342 bl_0_343
+ br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345 bl_0_346 br_0_346
+ bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349 br_0_349 bl_0_350
+ br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352 bl_0_353 br_0_353
+ bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356 br_0_356 bl_0_357
+ br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359 bl_0_360 br_0_360
+ bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363 br_0_363 bl_0_364
+ br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366 bl_0_367 br_0_367
+ bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370 br_0_370 bl_0_371
+ br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373 bl_0_374 br_0_374
+ bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377 br_0_377 bl_0_378
+ br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380 bl_0_381 br_0_381
+ bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384 br_0_384 bl_0_385
+ br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387 bl_0_388 br_0_388
+ bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391 br_0_391 bl_0_392
+ br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394 bl_0_395 br_0_395
+ bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398 br_0_398 bl_0_399
+ br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401 bl_0_402 br_0_402
+ bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405 br_0_405 bl_0_406
+ br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408 bl_0_409 br_0_409
+ bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412 br_0_412 bl_0_413
+ br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415 bl_0_416 br_0_416
+ bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419 br_0_419 bl_0_420
+ br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422 bl_0_423 br_0_423
+ bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426 br_0_426 bl_0_427
+ br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429 bl_0_430 br_0_430
+ bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433 br_0_433 bl_0_434
+ br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436 bl_0_437 br_0_437
+ bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440 br_0_440 bl_0_441
+ br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443 bl_0_444 br_0_444
+ bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447 br_0_447 bl_0_448
+ br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450 bl_0_451 br_0_451
+ bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454 br_0_454 bl_0_455
+ br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457 bl_0_458 br_0_458
+ bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461 br_0_461 bl_0_462
+ br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464 bl_0_465 br_0_465
+ bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468 br_0_468 bl_0_469
+ br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471 bl_0_472 br_0_472
+ bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475 br_0_475 bl_0_476
+ br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478 bl_0_479 br_0_479
+ bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482 br_0_482 bl_0_483
+ br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485 bl_0_486 br_0_486
+ bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489 br_0_489 bl_0_490
+ br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492 bl_0_493 br_0_493
+ bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496 br_0_496 bl_0_497
+ br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499 bl_0_500 br_0_500
+ bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503 br_0_503 bl_0_504
+ br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506 bl_0_507 br_0_507
+ bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510 br_0_510 bl_0_511
+ br_0_511 bl_0_512 br_0_512 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INOUT : bl_0_257 
* INOUT : br_0_257 
* INOUT : bl_0_258 
* INOUT : br_0_258 
* INOUT : bl_0_259 
* INOUT : br_0_259 
* INOUT : bl_0_260 
* INOUT : br_0_260 
* INOUT : bl_0_261 
* INOUT : br_0_261 
* INOUT : bl_0_262 
* INOUT : br_0_262 
* INOUT : bl_0_263 
* INOUT : br_0_263 
* INOUT : bl_0_264 
* INOUT : br_0_264 
* INOUT : bl_0_265 
* INOUT : br_0_265 
* INOUT : bl_0_266 
* INOUT : br_0_266 
* INOUT : bl_0_267 
* INOUT : br_0_267 
* INOUT : bl_0_268 
* INOUT : br_0_268 
* INOUT : bl_0_269 
* INOUT : br_0_269 
* INOUT : bl_0_270 
* INOUT : br_0_270 
* INOUT : bl_0_271 
* INOUT : br_0_271 
* INOUT : bl_0_272 
* INOUT : br_0_272 
* INOUT : bl_0_273 
* INOUT : br_0_273 
* INOUT : bl_0_274 
* INOUT : br_0_274 
* INOUT : bl_0_275 
* INOUT : br_0_275 
* INOUT : bl_0_276 
* INOUT : br_0_276 
* INOUT : bl_0_277 
* INOUT : br_0_277 
* INOUT : bl_0_278 
* INOUT : br_0_278 
* INOUT : bl_0_279 
* INOUT : br_0_279 
* INOUT : bl_0_280 
* INOUT : br_0_280 
* INOUT : bl_0_281 
* INOUT : br_0_281 
* INOUT : bl_0_282 
* INOUT : br_0_282 
* INOUT : bl_0_283 
* INOUT : br_0_283 
* INOUT : bl_0_284 
* INOUT : br_0_284 
* INOUT : bl_0_285 
* INOUT : br_0_285 
* INOUT : bl_0_286 
* INOUT : br_0_286 
* INOUT : bl_0_287 
* INOUT : br_0_287 
* INOUT : bl_0_288 
* INOUT : br_0_288 
* INOUT : bl_0_289 
* INOUT : br_0_289 
* INOUT : bl_0_290 
* INOUT : br_0_290 
* INOUT : bl_0_291 
* INOUT : br_0_291 
* INOUT : bl_0_292 
* INOUT : br_0_292 
* INOUT : bl_0_293 
* INOUT : br_0_293 
* INOUT : bl_0_294 
* INOUT : br_0_294 
* INOUT : bl_0_295 
* INOUT : br_0_295 
* INOUT : bl_0_296 
* INOUT : br_0_296 
* INOUT : bl_0_297 
* INOUT : br_0_297 
* INOUT : bl_0_298 
* INOUT : br_0_298 
* INOUT : bl_0_299 
* INOUT : br_0_299 
* INOUT : bl_0_300 
* INOUT : br_0_300 
* INOUT : bl_0_301 
* INOUT : br_0_301 
* INOUT : bl_0_302 
* INOUT : br_0_302 
* INOUT : bl_0_303 
* INOUT : br_0_303 
* INOUT : bl_0_304 
* INOUT : br_0_304 
* INOUT : bl_0_305 
* INOUT : br_0_305 
* INOUT : bl_0_306 
* INOUT : br_0_306 
* INOUT : bl_0_307 
* INOUT : br_0_307 
* INOUT : bl_0_308 
* INOUT : br_0_308 
* INOUT : bl_0_309 
* INOUT : br_0_309 
* INOUT : bl_0_310 
* INOUT : br_0_310 
* INOUT : bl_0_311 
* INOUT : br_0_311 
* INOUT : bl_0_312 
* INOUT : br_0_312 
* INOUT : bl_0_313 
* INOUT : br_0_313 
* INOUT : bl_0_314 
* INOUT : br_0_314 
* INOUT : bl_0_315 
* INOUT : br_0_315 
* INOUT : bl_0_316 
* INOUT : br_0_316 
* INOUT : bl_0_317 
* INOUT : br_0_317 
* INOUT : bl_0_318 
* INOUT : br_0_318 
* INOUT : bl_0_319 
* INOUT : br_0_319 
* INOUT : bl_0_320 
* INOUT : br_0_320 
* INOUT : bl_0_321 
* INOUT : br_0_321 
* INOUT : bl_0_322 
* INOUT : br_0_322 
* INOUT : bl_0_323 
* INOUT : br_0_323 
* INOUT : bl_0_324 
* INOUT : br_0_324 
* INOUT : bl_0_325 
* INOUT : br_0_325 
* INOUT : bl_0_326 
* INOUT : br_0_326 
* INOUT : bl_0_327 
* INOUT : br_0_327 
* INOUT : bl_0_328 
* INOUT : br_0_328 
* INOUT : bl_0_329 
* INOUT : br_0_329 
* INOUT : bl_0_330 
* INOUT : br_0_330 
* INOUT : bl_0_331 
* INOUT : br_0_331 
* INOUT : bl_0_332 
* INOUT : br_0_332 
* INOUT : bl_0_333 
* INOUT : br_0_333 
* INOUT : bl_0_334 
* INOUT : br_0_334 
* INOUT : bl_0_335 
* INOUT : br_0_335 
* INOUT : bl_0_336 
* INOUT : br_0_336 
* INOUT : bl_0_337 
* INOUT : br_0_337 
* INOUT : bl_0_338 
* INOUT : br_0_338 
* INOUT : bl_0_339 
* INOUT : br_0_339 
* INOUT : bl_0_340 
* INOUT : br_0_340 
* INOUT : bl_0_341 
* INOUT : br_0_341 
* INOUT : bl_0_342 
* INOUT : br_0_342 
* INOUT : bl_0_343 
* INOUT : br_0_343 
* INOUT : bl_0_344 
* INOUT : br_0_344 
* INOUT : bl_0_345 
* INOUT : br_0_345 
* INOUT : bl_0_346 
* INOUT : br_0_346 
* INOUT : bl_0_347 
* INOUT : br_0_347 
* INOUT : bl_0_348 
* INOUT : br_0_348 
* INOUT : bl_0_349 
* INOUT : br_0_349 
* INOUT : bl_0_350 
* INOUT : br_0_350 
* INOUT : bl_0_351 
* INOUT : br_0_351 
* INOUT : bl_0_352 
* INOUT : br_0_352 
* INOUT : bl_0_353 
* INOUT : br_0_353 
* INOUT : bl_0_354 
* INOUT : br_0_354 
* INOUT : bl_0_355 
* INOUT : br_0_355 
* INOUT : bl_0_356 
* INOUT : br_0_356 
* INOUT : bl_0_357 
* INOUT : br_0_357 
* INOUT : bl_0_358 
* INOUT : br_0_358 
* INOUT : bl_0_359 
* INOUT : br_0_359 
* INOUT : bl_0_360 
* INOUT : br_0_360 
* INOUT : bl_0_361 
* INOUT : br_0_361 
* INOUT : bl_0_362 
* INOUT : br_0_362 
* INOUT : bl_0_363 
* INOUT : br_0_363 
* INOUT : bl_0_364 
* INOUT : br_0_364 
* INOUT : bl_0_365 
* INOUT : br_0_365 
* INOUT : bl_0_366 
* INOUT : br_0_366 
* INOUT : bl_0_367 
* INOUT : br_0_367 
* INOUT : bl_0_368 
* INOUT : br_0_368 
* INOUT : bl_0_369 
* INOUT : br_0_369 
* INOUT : bl_0_370 
* INOUT : br_0_370 
* INOUT : bl_0_371 
* INOUT : br_0_371 
* INOUT : bl_0_372 
* INOUT : br_0_372 
* INOUT : bl_0_373 
* INOUT : br_0_373 
* INOUT : bl_0_374 
* INOUT : br_0_374 
* INOUT : bl_0_375 
* INOUT : br_0_375 
* INOUT : bl_0_376 
* INOUT : br_0_376 
* INOUT : bl_0_377 
* INOUT : br_0_377 
* INOUT : bl_0_378 
* INOUT : br_0_378 
* INOUT : bl_0_379 
* INOUT : br_0_379 
* INOUT : bl_0_380 
* INOUT : br_0_380 
* INOUT : bl_0_381 
* INOUT : br_0_381 
* INOUT : bl_0_382 
* INOUT : br_0_382 
* INOUT : bl_0_383 
* INOUT : br_0_383 
* INOUT : bl_0_384 
* INOUT : br_0_384 
* INOUT : bl_0_385 
* INOUT : br_0_385 
* INOUT : bl_0_386 
* INOUT : br_0_386 
* INOUT : bl_0_387 
* INOUT : br_0_387 
* INOUT : bl_0_388 
* INOUT : br_0_388 
* INOUT : bl_0_389 
* INOUT : br_0_389 
* INOUT : bl_0_390 
* INOUT : br_0_390 
* INOUT : bl_0_391 
* INOUT : br_0_391 
* INOUT : bl_0_392 
* INOUT : br_0_392 
* INOUT : bl_0_393 
* INOUT : br_0_393 
* INOUT : bl_0_394 
* INOUT : br_0_394 
* INOUT : bl_0_395 
* INOUT : br_0_395 
* INOUT : bl_0_396 
* INOUT : br_0_396 
* INOUT : bl_0_397 
* INOUT : br_0_397 
* INOUT : bl_0_398 
* INOUT : br_0_398 
* INOUT : bl_0_399 
* INOUT : br_0_399 
* INOUT : bl_0_400 
* INOUT : br_0_400 
* INOUT : bl_0_401 
* INOUT : br_0_401 
* INOUT : bl_0_402 
* INOUT : br_0_402 
* INOUT : bl_0_403 
* INOUT : br_0_403 
* INOUT : bl_0_404 
* INOUT : br_0_404 
* INOUT : bl_0_405 
* INOUT : br_0_405 
* INOUT : bl_0_406 
* INOUT : br_0_406 
* INOUT : bl_0_407 
* INOUT : br_0_407 
* INOUT : bl_0_408 
* INOUT : br_0_408 
* INOUT : bl_0_409 
* INOUT : br_0_409 
* INOUT : bl_0_410 
* INOUT : br_0_410 
* INOUT : bl_0_411 
* INOUT : br_0_411 
* INOUT : bl_0_412 
* INOUT : br_0_412 
* INOUT : bl_0_413 
* INOUT : br_0_413 
* INOUT : bl_0_414 
* INOUT : br_0_414 
* INOUT : bl_0_415 
* INOUT : br_0_415 
* INOUT : bl_0_416 
* INOUT : br_0_416 
* INOUT : bl_0_417 
* INOUT : br_0_417 
* INOUT : bl_0_418 
* INOUT : br_0_418 
* INOUT : bl_0_419 
* INOUT : br_0_419 
* INOUT : bl_0_420 
* INOUT : br_0_420 
* INOUT : bl_0_421 
* INOUT : br_0_421 
* INOUT : bl_0_422 
* INOUT : br_0_422 
* INOUT : bl_0_423 
* INOUT : br_0_423 
* INOUT : bl_0_424 
* INOUT : br_0_424 
* INOUT : bl_0_425 
* INOUT : br_0_425 
* INOUT : bl_0_426 
* INOUT : br_0_426 
* INOUT : bl_0_427 
* INOUT : br_0_427 
* INOUT : bl_0_428 
* INOUT : br_0_428 
* INOUT : bl_0_429 
* INOUT : br_0_429 
* INOUT : bl_0_430 
* INOUT : br_0_430 
* INOUT : bl_0_431 
* INOUT : br_0_431 
* INOUT : bl_0_432 
* INOUT : br_0_432 
* INOUT : bl_0_433 
* INOUT : br_0_433 
* INOUT : bl_0_434 
* INOUT : br_0_434 
* INOUT : bl_0_435 
* INOUT : br_0_435 
* INOUT : bl_0_436 
* INOUT : br_0_436 
* INOUT : bl_0_437 
* INOUT : br_0_437 
* INOUT : bl_0_438 
* INOUT : br_0_438 
* INOUT : bl_0_439 
* INOUT : br_0_439 
* INOUT : bl_0_440 
* INOUT : br_0_440 
* INOUT : bl_0_441 
* INOUT : br_0_441 
* INOUT : bl_0_442 
* INOUT : br_0_442 
* INOUT : bl_0_443 
* INOUT : br_0_443 
* INOUT : bl_0_444 
* INOUT : br_0_444 
* INOUT : bl_0_445 
* INOUT : br_0_445 
* INOUT : bl_0_446 
* INOUT : br_0_446 
* INOUT : bl_0_447 
* INOUT : br_0_447 
* INOUT : bl_0_448 
* INOUT : br_0_448 
* INOUT : bl_0_449 
* INOUT : br_0_449 
* INOUT : bl_0_450 
* INOUT : br_0_450 
* INOUT : bl_0_451 
* INOUT : br_0_451 
* INOUT : bl_0_452 
* INOUT : br_0_452 
* INOUT : bl_0_453 
* INOUT : br_0_453 
* INOUT : bl_0_454 
* INOUT : br_0_454 
* INOUT : bl_0_455 
* INOUT : br_0_455 
* INOUT : bl_0_456 
* INOUT : br_0_456 
* INOUT : bl_0_457 
* INOUT : br_0_457 
* INOUT : bl_0_458 
* INOUT : br_0_458 
* INOUT : bl_0_459 
* INOUT : br_0_459 
* INOUT : bl_0_460 
* INOUT : br_0_460 
* INOUT : bl_0_461 
* INOUT : br_0_461 
* INOUT : bl_0_462 
* INOUT : br_0_462 
* INOUT : bl_0_463 
* INOUT : br_0_463 
* INOUT : bl_0_464 
* INOUT : br_0_464 
* INOUT : bl_0_465 
* INOUT : br_0_465 
* INOUT : bl_0_466 
* INOUT : br_0_466 
* INOUT : bl_0_467 
* INOUT : br_0_467 
* INOUT : bl_0_468 
* INOUT : br_0_468 
* INOUT : bl_0_469 
* INOUT : br_0_469 
* INOUT : bl_0_470 
* INOUT : br_0_470 
* INOUT : bl_0_471 
* INOUT : br_0_471 
* INOUT : bl_0_472 
* INOUT : br_0_472 
* INOUT : bl_0_473 
* INOUT : br_0_473 
* INOUT : bl_0_474 
* INOUT : br_0_474 
* INOUT : bl_0_475 
* INOUT : br_0_475 
* INOUT : bl_0_476 
* INOUT : br_0_476 
* INOUT : bl_0_477 
* INOUT : br_0_477 
* INOUT : bl_0_478 
* INOUT : br_0_478 
* INOUT : bl_0_479 
* INOUT : br_0_479 
* INOUT : bl_0_480 
* INOUT : br_0_480 
* INOUT : bl_0_481 
* INOUT : br_0_481 
* INOUT : bl_0_482 
* INOUT : br_0_482 
* INOUT : bl_0_483 
* INOUT : br_0_483 
* INOUT : bl_0_484 
* INOUT : br_0_484 
* INOUT : bl_0_485 
* INOUT : br_0_485 
* INOUT : bl_0_486 
* INOUT : br_0_486 
* INOUT : bl_0_487 
* INOUT : br_0_487 
* INOUT : bl_0_488 
* INOUT : br_0_488 
* INOUT : bl_0_489 
* INOUT : br_0_489 
* INOUT : bl_0_490 
* INOUT : br_0_490 
* INOUT : bl_0_491 
* INOUT : br_0_491 
* INOUT : bl_0_492 
* INOUT : br_0_492 
* INOUT : bl_0_493 
* INOUT : br_0_493 
* INOUT : bl_0_494 
* INOUT : br_0_494 
* INOUT : bl_0_495 
* INOUT : br_0_495 
* INOUT : bl_0_496 
* INOUT : br_0_496 
* INOUT : bl_0_497 
* INOUT : br_0_497 
* INOUT : bl_0_498 
* INOUT : br_0_498 
* INOUT : bl_0_499 
* INOUT : br_0_499 
* INOUT : bl_0_500 
* INOUT : br_0_500 
* INOUT : bl_0_501 
* INOUT : br_0_501 
* INOUT : bl_0_502 
* INOUT : br_0_502 
* INOUT : bl_0_503 
* INOUT : br_0_503 
* INOUT : bl_0_504 
* INOUT : br_0_504 
* INOUT : bl_0_505 
* INOUT : br_0_505 
* INOUT : bl_0_506 
* INOUT : br_0_506 
* INOUT : bl_0_507 
* INOUT : br_0_507 
* INOUT : bl_0_508 
* INOUT : br_0_508 
* INOUT : bl_0_509 
* INOUT : br_0_509 
* INOUT : bl_0_510 
* INOUT : br_0_510 
* INOUT : bl_0_511 
* INOUT : br_0_511 
* INOUT : bl_0_512 
* INOUT : br_0_512 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c256
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c257
+ bl_0_257 br_0_257 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c258
+ bl_0_258 br_0_258 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c259
+ bl_0_259 br_0_259 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c260
+ bl_0_260 br_0_260 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c261
+ bl_0_261 br_0_261 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c262
+ bl_0_262 br_0_262 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c263
+ bl_0_263 br_0_263 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c264
+ bl_0_264 br_0_264 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c265
+ bl_0_265 br_0_265 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c266
+ bl_0_266 br_0_266 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c267
+ bl_0_267 br_0_267 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c268
+ bl_0_268 br_0_268 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c269
+ bl_0_269 br_0_269 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c270
+ bl_0_270 br_0_270 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c271
+ bl_0_271 br_0_271 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c272
+ bl_0_272 br_0_272 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c273
+ bl_0_273 br_0_273 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c274
+ bl_0_274 br_0_274 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c275
+ bl_0_275 br_0_275 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c276
+ bl_0_276 br_0_276 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c277
+ bl_0_277 br_0_277 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c278
+ bl_0_278 br_0_278 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c279
+ bl_0_279 br_0_279 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c280
+ bl_0_280 br_0_280 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c281
+ bl_0_281 br_0_281 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c282
+ bl_0_282 br_0_282 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c283
+ bl_0_283 br_0_283 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c284
+ bl_0_284 br_0_284 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c285
+ bl_0_285 br_0_285 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c286
+ bl_0_286 br_0_286 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c287
+ bl_0_287 br_0_287 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c288
+ bl_0_288 br_0_288 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c289
+ bl_0_289 br_0_289 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c290
+ bl_0_290 br_0_290 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c291
+ bl_0_291 br_0_291 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c292
+ bl_0_292 br_0_292 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c293
+ bl_0_293 br_0_293 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c294
+ bl_0_294 br_0_294 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c295
+ bl_0_295 br_0_295 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c296
+ bl_0_296 br_0_296 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c297
+ bl_0_297 br_0_297 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c298
+ bl_0_298 br_0_298 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c299
+ bl_0_299 br_0_299 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c300
+ bl_0_300 br_0_300 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c301
+ bl_0_301 br_0_301 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c302
+ bl_0_302 br_0_302 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c303
+ bl_0_303 br_0_303 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c304
+ bl_0_304 br_0_304 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c305
+ bl_0_305 br_0_305 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c306
+ bl_0_306 br_0_306 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c307
+ bl_0_307 br_0_307 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c308
+ bl_0_308 br_0_308 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c309
+ bl_0_309 br_0_309 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c310
+ bl_0_310 br_0_310 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c311
+ bl_0_311 br_0_311 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c312
+ bl_0_312 br_0_312 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c313
+ bl_0_313 br_0_313 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c314
+ bl_0_314 br_0_314 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c315
+ bl_0_315 br_0_315 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c316
+ bl_0_316 br_0_316 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c317
+ bl_0_317 br_0_317 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c318
+ bl_0_318 br_0_318 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c319
+ bl_0_319 br_0_319 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c320
+ bl_0_320 br_0_320 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c321
+ bl_0_321 br_0_321 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c322
+ bl_0_322 br_0_322 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c323
+ bl_0_323 br_0_323 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c324
+ bl_0_324 br_0_324 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c325
+ bl_0_325 br_0_325 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c326
+ bl_0_326 br_0_326 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c327
+ bl_0_327 br_0_327 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c328
+ bl_0_328 br_0_328 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c329
+ bl_0_329 br_0_329 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c330
+ bl_0_330 br_0_330 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c331
+ bl_0_331 br_0_331 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c332
+ bl_0_332 br_0_332 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c333
+ bl_0_333 br_0_333 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c334
+ bl_0_334 br_0_334 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c335
+ bl_0_335 br_0_335 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c336
+ bl_0_336 br_0_336 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c337
+ bl_0_337 br_0_337 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c338
+ bl_0_338 br_0_338 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c339
+ bl_0_339 br_0_339 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c340
+ bl_0_340 br_0_340 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c341
+ bl_0_341 br_0_341 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c342
+ bl_0_342 br_0_342 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c343
+ bl_0_343 br_0_343 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c344
+ bl_0_344 br_0_344 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c345
+ bl_0_345 br_0_345 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c346
+ bl_0_346 br_0_346 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c347
+ bl_0_347 br_0_347 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c348
+ bl_0_348 br_0_348 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c349
+ bl_0_349 br_0_349 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c350
+ bl_0_350 br_0_350 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c351
+ bl_0_351 br_0_351 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c352
+ bl_0_352 br_0_352 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c353
+ bl_0_353 br_0_353 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c354
+ bl_0_354 br_0_354 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c355
+ bl_0_355 br_0_355 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c356
+ bl_0_356 br_0_356 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c357
+ bl_0_357 br_0_357 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c358
+ bl_0_358 br_0_358 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c359
+ bl_0_359 br_0_359 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c360
+ bl_0_360 br_0_360 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c361
+ bl_0_361 br_0_361 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c362
+ bl_0_362 br_0_362 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c363
+ bl_0_363 br_0_363 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c364
+ bl_0_364 br_0_364 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c365
+ bl_0_365 br_0_365 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c366
+ bl_0_366 br_0_366 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c367
+ bl_0_367 br_0_367 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c368
+ bl_0_368 br_0_368 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c369
+ bl_0_369 br_0_369 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c370
+ bl_0_370 br_0_370 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c371
+ bl_0_371 br_0_371 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c372
+ bl_0_372 br_0_372 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c373
+ bl_0_373 br_0_373 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c374
+ bl_0_374 br_0_374 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c375
+ bl_0_375 br_0_375 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c376
+ bl_0_376 br_0_376 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c377
+ bl_0_377 br_0_377 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c378
+ bl_0_378 br_0_378 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c379
+ bl_0_379 br_0_379 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c380
+ bl_0_380 br_0_380 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c381
+ bl_0_381 br_0_381 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c382
+ bl_0_382 br_0_382 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c383
+ bl_0_383 br_0_383 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c384
+ bl_0_384 br_0_384 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c385
+ bl_0_385 br_0_385 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c386
+ bl_0_386 br_0_386 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c387
+ bl_0_387 br_0_387 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c388
+ bl_0_388 br_0_388 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c389
+ bl_0_389 br_0_389 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c390
+ bl_0_390 br_0_390 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c391
+ bl_0_391 br_0_391 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c392
+ bl_0_392 br_0_392 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c393
+ bl_0_393 br_0_393 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c394
+ bl_0_394 br_0_394 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c395
+ bl_0_395 br_0_395 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c396
+ bl_0_396 br_0_396 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c397
+ bl_0_397 br_0_397 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c398
+ bl_0_398 br_0_398 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c399
+ bl_0_399 br_0_399 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c400
+ bl_0_400 br_0_400 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c401
+ bl_0_401 br_0_401 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c402
+ bl_0_402 br_0_402 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c403
+ bl_0_403 br_0_403 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c404
+ bl_0_404 br_0_404 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c405
+ bl_0_405 br_0_405 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c406
+ bl_0_406 br_0_406 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c407
+ bl_0_407 br_0_407 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c408
+ bl_0_408 br_0_408 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c409
+ bl_0_409 br_0_409 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c410
+ bl_0_410 br_0_410 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c411
+ bl_0_411 br_0_411 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c412
+ bl_0_412 br_0_412 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c413
+ bl_0_413 br_0_413 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c414
+ bl_0_414 br_0_414 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c415
+ bl_0_415 br_0_415 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c416
+ bl_0_416 br_0_416 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c417
+ bl_0_417 br_0_417 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c418
+ bl_0_418 br_0_418 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c419
+ bl_0_419 br_0_419 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c420
+ bl_0_420 br_0_420 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c421
+ bl_0_421 br_0_421 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c422
+ bl_0_422 br_0_422 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c423
+ bl_0_423 br_0_423 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c424
+ bl_0_424 br_0_424 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c425
+ bl_0_425 br_0_425 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c426
+ bl_0_426 br_0_426 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c427
+ bl_0_427 br_0_427 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c428
+ bl_0_428 br_0_428 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c429
+ bl_0_429 br_0_429 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c430
+ bl_0_430 br_0_430 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c431
+ bl_0_431 br_0_431 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c432
+ bl_0_432 br_0_432 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c433
+ bl_0_433 br_0_433 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c434
+ bl_0_434 br_0_434 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c435
+ bl_0_435 br_0_435 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c436
+ bl_0_436 br_0_436 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c437
+ bl_0_437 br_0_437 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c438
+ bl_0_438 br_0_438 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c439
+ bl_0_439 br_0_439 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c440
+ bl_0_440 br_0_440 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c441
+ bl_0_441 br_0_441 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c442
+ bl_0_442 br_0_442 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c443
+ bl_0_443 br_0_443 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c444
+ bl_0_444 br_0_444 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c445
+ bl_0_445 br_0_445 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c446
+ bl_0_446 br_0_446 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c447
+ bl_0_447 br_0_447 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c448
+ bl_0_448 br_0_448 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c449
+ bl_0_449 br_0_449 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c450
+ bl_0_450 br_0_450 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c451
+ bl_0_451 br_0_451 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c452
+ bl_0_452 br_0_452 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c453
+ bl_0_453 br_0_453 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c454
+ bl_0_454 br_0_454 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c455
+ bl_0_455 br_0_455 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c456
+ bl_0_456 br_0_456 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c457
+ bl_0_457 br_0_457 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c458
+ bl_0_458 br_0_458 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c459
+ bl_0_459 br_0_459 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c460
+ bl_0_460 br_0_460 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c461
+ bl_0_461 br_0_461 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c462
+ bl_0_462 br_0_462 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c463
+ bl_0_463 br_0_463 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c464
+ bl_0_464 br_0_464 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c465
+ bl_0_465 br_0_465 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c466
+ bl_0_466 br_0_466 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c467
+ bl_0_467 br_0_467 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c468
+ bl_0_468 br_0_468 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c469
+ bl_0_469 br_0_469 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c470
+ bl_0_470 br_0_470 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c471
+ bl_0_471 br_0_471 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c472
+ bl_0_472 br_0_472 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c473
+ bl_0_473 br_0_473 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c474
+ bl_0_474 br_0_474 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c475
+ bl_0_475 br_0_475 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c476
+ bl_0_476 br_0_476 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c477
+ bl_0_477 br_0_477 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c478
+ bl_0_478 br_0_478 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c479
+ bl_0_479 br_0_479 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c480
+ bl_0_480 br_0_480 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c481
+ bl_0_481 br_0_481 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c482
+ bl_0_482 br_0_482 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c483
+ bl_0_483 br_0_483 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c484
+ bl_0_484 br_0_484 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c485
+ bl_0_485 br_0_485 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c486
+ bl_0_486 br_0_486 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c487
+ bl_0_487 br_0_487 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c488
+ bl_0_488 br_0_488 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c489
+ bl_0_489 br_0_489 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c490
+ bl_0_490 br_0_490 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c491
+ bl_0_491 br_0_491 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c492
+ bl_0_492 br_0_492 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c493
+ bl_0_493 br_0_493 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c494
+ bl_0_494 br_0_494 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c495
+ bl_0_495 br_0_495 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c496
+ bl_0_496 br_0_496 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c497
+ bl_0_497 br_0_497 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c498
+ bl_0_498 br_0_498 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c499
+ bl_0_499 br_0_499 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c500
+ bl_0_500 br_0_500 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c501
+ bl_0_501 br_0_501 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c502
+ bl_0_502 br_0_502 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c503
+ bl_0_503 br_0_503 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c504
+ bl_0_504 br_0_504 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c505
+ bl_0_505 br_0_505 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c506
+ bl_0_506 br_0_506 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c507
+ bl_0_507 br_0_507 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c508
+ bl_0_508 br_0_508 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c509
+ bl_0_509 br_0_509 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c510
+ bl_0_510 br_0_510 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c511
+ bl_0_511 br_0_511 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c512
+ bl_0_512 br_0_512 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS freepdk45_sram_1rw0r_45x512_dummy_array_1

.SUBCKT freepdk45_sram_1rw0r_45x512_dummy_array_0
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258 br_0_258 bl_0_259
+ br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261 bl_0_262 br_0_262
+ bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265 br_0_265 bl_0_266
+ br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268 bl_0_269 br_0_269
+ bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272 br_0_272 bl_0_273
+ br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275 bl_0_276 br_0_276
+ bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279 br_0_279 bl_0_280
+ br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282 bl_0_283 br_0_283
+ bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286 br_0_286 bl_0_287
+ br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289 bl_0_290 br_0_290
+ bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293 br_0_293 bl_0_294
+ br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296 bl_0_297 br_0_297
+ bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300 br_0_300 bl_0_301
+ br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303 bl_0_304 br_0_304
+ bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307 br_0_307 bl_0_308
+ br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310 bl_0_311 br_0_311
+ bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314 br_0_314 bl_0_315
+ br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317 bl_0_318 br_0_318
+ bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321 br_0_321 bl_0_322
+ br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324 bl_0_325 br_0_325
+ bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328 br_0_328 bl_0_329
+ br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331 bl_0_332 br_0_332
+ bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335 br_0_335 bl_0_336
+ br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338 bl_0_339 br_0_339
+ bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342 br_0_342 bl_0_343
+ br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345 bl_0_346 br_0_346
+ bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349 br_0_349 bl_0_350
+ br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352 bl_0_353 br_0_353
+ bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356 br_0_356 bl_0_357
+ br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359 bl_0_360 br_0_360
+ bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363 br_0_363 bl_0_364
+ br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366 bl_0_367 br_0_367
+ bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370 br_0_370 bl_0_371
+ br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373 bl_0_374 br_0_374
+ bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377 br_0_377 bl_0_378
+ br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380 bl_0_381 br_0_381
+ bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384 br_0_384 bl_0_385
+ br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387 bl_0_388 br_0_388
+ bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391 br_0_391 bl_0_392
+ br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394 bl_0_395 br_0_395
+ bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398 br_0_398 bl_0_399
+ br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401 bl_0_402 br_0_402
+ bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405 br_0_405 bl_0_406
+ br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408 bl_0_409 br_0_409
+ bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412 br_0_412 bl_0_413
+ br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415 bl_0_416 br_0_416
+ bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419 br_0_419 bl_0_420
+ br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422 bl_0_423 br_0_423
+ bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426 br_0_426 bl_0_427
+ br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429 bl_0_430 br_0_430
+ bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433 br_0_433 bl_0_434
+ br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436 bl_0_437 br_0_437
+ bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440 br_0_440 bl_0_441
+ br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443 bl_0_444 br_0_444
+ bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447 br_0_447 bl_0_448
+ br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450 bl_0_451 br_0_451
+ bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454 br_0_454 bl_0_455
+ br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457 bl_0_458 br_0_458
+ bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461 br_0_461 bl_0_462
+ br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464 bl_0_465 br_0_465
+ bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468 br_0_468 bl_0_469
+ br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471 bl_0_472 br_0_472
+ bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475 br_0_475 bl_0_476
+ br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478 bl_0_479 br_0_479
+ bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482 br_0_482 bl_0_483
+ br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485 bl_0_486 br_0_486
+ bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489 br_0_489 bl_0_490
+ br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492 bl_0_493 br_0_493
+ bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496 br_0_496 bl_0_497
+ br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499 bl_0_500 br_0_500
+ bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503 br_0_503 bl_0_504
+ br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506 bl_0_507 br_0_507
+ bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510 br_0_510 bl_0_511
+ br_0_511 bl_0_512 br_0_512 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INOUT : bl_0_257 
* INOUT : br_0_257 
* INOUT : bl_0_258 
* INOUT : br_0_258 
* INOUT : bl_0_259 
* INOUT : br_0_259 
* INOUT : bl_0_260 
* INOUT : br_0_260 
* INOUT : bl_0_261 
* INOUT : br_0_261 
* INOUT : bl_0_262 
* INOUT : br_0_262 
* INOUT : bl_0_263 
* INOUT : br_0_263 
* INOUT : bl_0_264 
* INOUT : br_0_264 
* INOUT : bl_0_265 
* INOUT : br_0_265 
* INOUT : bl_0_266 
* INOUT : br_0_266 
* INOUT : bl_0_267 
* INOUT : br_0_267 
* INOUT : bl_0_268 
* INOUT : br_0_268 
* INOUT : bl_0_269 
* INOUT : br_0_269 
* INOUT : bl_0_270 
* INOUT : br_0_270 
* INOUT : bl_0_271 
* INOUT : br_0_271 
* INOUT : bl_0_272 
* INOUT : br_0_272 
* INOUT : bl_0_273 
* INOUT : br_0_273 
* INOUT : bl_0_274 
* INOUT : br_0_274 
* INOUT : bl_0_275 
* INOUT : br_0_275 
* INOUT : bl_0_276 
* INOUT : br_0_276 
* INOUT : bl_0_277 
* INOUT : br_0_277 
* INOUT : bl_0_278 
* INOUT : br_0_278 
* INOUT : bl_0_279 
* INOUT : br_0_279 
* INOUT : bl_0_280 
* INOUT : br_0_280 
* INOUT : bl_0_281 
* INOUT : br_0_281 
* INOUT : bl_0_282 
* INOUT : br_0_282 
* INOUT : bl_0_283 
* INOUT : br_0_283 
* INOUT : bl_0_284 
* INOUT : br_0_284 
* INOUT : bl_0_285 
* INOUT : br_0_285 
* INOUT : bl_0_286 
* INOUT : br_0_286 
* INOUT : bl_0_287 
* INOUT : br_0_287 
* INOUT : bl_0_288 
* INOUT : br_0_288 
* INOUT : bl_0_289 
* INOUT : br_0_289 
* INOUT : bl_0_290 
* INOUT : br_0_290 
* INOUT : bl_0_291 
* INOUT : br_0_291 
* INOUT : bl_0_292 
* INOUT : br_0_292 
* INOUT : bl_0_293 
* INOUT : br_0_293 
* INOUT : bl_0_294 
* INOUT : br_0_294 
* INOUT : bl_0_295 
* INOUT : br_0_295 
* INOUT : bl_0_296 
* INOUT : br_0_296 
* INOUT : bl_0_297 
* INOUT : br_0_297 
* INOUT : bl_0_298 
* INOUT : br_0_298 
* INOUT : bl_0_299 
* INOUT : br_0_299 
* INOUT : bl_0_300 
* INOUT : br_0_300 
* INOUT : bl_0_301 
* INOUT : br_0_301 
* INOUT : bl_0_302 
* INOUT : br_0_302 
* INOUT : bl_0_303 
* INOUT : br_0_303 
* INOUT : bl_0_304 
* INOUT : br_0_304 
* INOUT : bl_0_305 
* INOUT : br_0_305 
* INOUT : bl_0_306 
* INOUT : br_0_306 
* INOUT : bl_0_307 
* INOUT : br_0_307 
* INOUT : bl_0_308 
* INOUT : br_0_308 
* INOUT : bl_0_309 
* INOUT : br_0_309 
* INOUT : bl_0_310 
* INOUT : br_0_310 
* INOUT : bl_0_311 
* INOUT : br_0_311 
* INOUT : bl_0_312 
* INOUT : br_0_312 
* INOUT : bl_0_313 
* INOUT : br_0_313 
* INOUT : bl_0_314 
* INOUT : br_0_314 
* INOUT : bl_0_315 
* INOUT : br_0_315 
* INOUT : bl_0_316 
* INOUT : br_0_316 
* INOUT : bl_0_317 
* INOUT : br_0_317 
* INOUT : bl_0_318 
* INOUT : br_0_318 
* INOUT : bl_0_319 
* INOUT : br_0_319 
* INOUT : bl_0_320 
* INOUT : br_0_320 
* INOUT : bl_0_321 
* INOUT : br_0_321 
* INOUT : bl_0_322 
* INOUT : br_0_322 
* INOUT : bl_0_323 
* INOUT : br_0_323 
* INOUT : bl_0_324 
* INOUT : br_0_324 
* INOUT : bl_0_325 
* INOUT : br_0_325 
* INOUT : bl_0_326 
* INOUT : br_0_326 
* INOUT : bl_0_327 
* INOUT : br_0_327 
* INOUT : bl_0_328 
* INOUT : br_0_328 
* INOUT : bl_0_329 
* INOUT : br_0_329 
* INOUT : bl_0_330 
* INOUT : br_0_330 
* INOUT : bl_0_331 
* INOUT : br_0_331 
* INOUT : bl_0_332 
* INOUT : br_0_332 
* INOUT : bl_0_333 
* INOUT : br_0_333 
* INOUT : bl_0_334 
* INOUT : br_0_334 
* INOUT : bl_0_335 
* INOUT : br_0_335 
* INOUT : bl_0_336 
* INOUT : br_0_336 
* INOUT : bl_0_337 
* INOUT : br_0_337 
* INOUT : bl_0_338 
* INOUT : br_0_338 
* INOUT : bl_0_339 
* INOUT : br_0_339 
* INOUT : bl_0_340 
* INOUT : br_0_340 
* INOUT : bl_0_341 
* INOUT : br_0_341 
* INOUT : bl_0_342 
* INOUT : br_0_342 
* INOUT : bl_0_343 
* INOUT : br_0_343 
* INOUT : bl_0_344 
* INOUT : br_0_344 
* INOUT : bl_0_345 
* INOUT : br_0_345 
* INOUT : bl_0_346 
* INOUT : br_0_346 
* INOUT : bl_0_347 
* INOUT : br_0_347 
* INOUT : bl_0_348 
* INOUT : br_0_348 
* INOUT : bl_0_349 
* INOUT : br_0_349 
* INOUT : bl_0_350 
* INOUT : br_0_350 
* INOUT : bl_0_351 
* INOUT : br_0_351 
* INOUT : bl_0_352 
* INOUT : br_0_352 
* INOUT : bl_0_353 
* INOUT : br_0_353 
* INOUT : bl_0_354 
* INOUT : br_0_354 
* INOUT : bl_0_355 
* INOUT : br_0_355 
* INOUT : bl_0_356 
* INOUT : br_0_356 
* INOUT : bl_0_357 
* INOUT : br_0_357 
* INOUT : bl_0_358 
* INOUT : br_0_358 
* INOUT : bl_0_359 
* INOUT : br_0_359 
* INOUT : bl_0_360 
* INOUT : br_0_360 
* INOUT : bl_0_361 
* INOUT : br_0_361 
* INOUT : bl_0_362 
* INOUT : br_0_362 
* INOUT : bl_0_363 
* INOUT : br_0_363 
* INOUT : bl_0_364 
* INOUT : br_0_364 
* INOUT : bl_0_365 
* INOUT : br_0_365 
* INOUT : bl_0_366 
* INOUT : br_0_366 
* INOUT : bl_0_367 
* INOUT : br_0_367 
* INOUT : bl_0_368 
* INOUT : br_0_368 
* INOUT : bl_0_369 
* INOUT : br_0_369 
* INOUT : bl_0_370 
* INOUT : br_0_370 
* INOUT : bl_0_371 
* INOUT : br_0_371 
* INOUT : bl_0_372 
* INOUT : br_0_372 
* INOUT : bl_0_373 
* INOUT : br_0_373 
* INOUT : bl_0_374 
* INOUT : br_0_374 
* INOUT : bl_0_375 
* INOUT : br_0_375 
* INOUT : bl_0_376 
* INOUT : br_0_376 
* INOUT : bl_0_377 
* INOUT : br_0_377 
* INOUT : bl_0_378 
* INOUT : br_0_378 
* INOUT : bl_0_379 
* INOUT : br_0_379 
* INOUT : bl_0_380 
* INOUT : br_0_380 
* INOUT : bl_0_381 
* INOUT : br_0_381 
* INOUT : bl_0_382 
* INOUT : br_0_382 
* INOUT : bl_0_383 
* INOUT : br_0_383 
* INOUT : bl_0_384 
* INOUT : br_0_384 
* INOUT : bl_0_385 
* INOUT : br_0_385 
* INOUT : bl_0_386 
* INOUT : br_0_386 
* INOUT : bl_0_387 
* INOUT : br_0_387 
* INOUT : bl_0_388 
* INOUT : br_0_388 
* INOUT : bl_0_389 
* INOUT : br_0_389 
* INOUT : bl_0_390 
* INOUT : br_0_390 
* INOUT : bl_0_391 
* INOUT : br_0_391 
* INOUT : bl_0_392 
* INOUT : br_0_392 
* INOUT : bl_0_393 
* INOUT : br_0_393 
* INOUT : bl_0_394 
* INOUT : br_0_394 
* INOUT : bl_0_395 
* INOUT : br_0_395 
* INOUT : bl_0_396 
* INOUT : br_0_396 
* INOUT : bl_0_397 
* INOUT : br_0_397 
* INOUT : bl_0_398 
* INOUT : br_0_398 
* INOUT : bl_0_399 
* INOUT : br_0_399 
* INOUT : bl_0_400 
* INOUT : br_0_400 
* INOUT : bl_0_401 
* INOUT : br_0_401 
* INOUT : bl_0_402 
* INOUT : br_0_402 
* INOUT : bl_0_403 
* INOUT : br_0_403 
* INOUT : bl_0_404 
* INOUT : br_0_404 
* INOUT : bl_0_405 
* INOUT : br_0_405 
* INOUT : bl_0_406 
* INOUT : br_0_406 
* INOUT : bl_0_407 
* INOUT : br_0_407 
* INOUT : bl_0_408 
* INOUT : br_0_408 
* INOUT : bl_0_409 
* INOUT : br_0_409 
* INOUT : bl_0_410 
* INOUT : br_0_410 
* INOUT : bl_0_411 
* INOUT : br_0_411 
* INOUT : bl_0_412 
* INOUT : br_0_412 
* INOUT : bl_0_413 
* INOUT : br_0_413 
* INOUT : bl_0_414 
* INOUT : br_0_414 
* INOUT : bl_0_415 
* INOUT : br_0_415 
* INOUT : bl_0_416 
* INOUT : br_0_416 
* INOUT : bl_0_417 
* INOUT : br_0_417 
* INOUT : bl_0_418 
* INOUT : br_0_418 
* INOUT : bl_0_419 
* INOUT : br_0_419 
* INOUT : bl_0_420 
* INOUT : br_0_420 
* INOUT : bl_0_421 
* INOUT : br_0_421 
* INOUT : bl_0_422 
* INOUT : br_0_422 
* INOUT : bl_0_423 
* INOUT : br_0_423 
* INOUT : bl_0_424 
* INOUT : br_0_424 
* INOUT : bl_0_425 
* INOUT : br_0_425 
* INOUT : bl_0_426 
* INOUT : br_0_426 
* INOUT : bl_0_427 
* INOUT : br_0_427 
* INOUT : bl_0_428 
* INOUT : br_0_428 
* INOUT : bl_0_429 
* INOUT : br_0_429 
* INOUT : bl_0_430 
* INOUT : br_0_430 
* INOUT : bl_0_431 
* INOUT : br_0_431 
* INOUT : bl_0_432 
* INOUT : br_0_432 
* INOUT : bl_0_433 
* INOUT : br_0_433 
* INOUT : bl_0_434 
* INOUT : br_0_434 
* INOUT : bl_0_435 
* INOUT : br_0_435 
* INOUT : bl_0_436 
* INOUT : br_0_436 
* INOUT : bl_0_437 
* INOUT : br_0_437 
* INOUT : bl_0_438 
* INOUT : br_0_438 
* INOUT : bl_0_439 
* INOUT : br_0_439 
* INOUT : bl_0_440 
* INOUT : br_0_440 
* INOUT : bl_0_441 
* INOUT : br_0_441 
* INOUT : bl_0_442 
* INOUT : br_0_442 
* INOUT : bl_0_443 
* INOUT : br_0_443 
* INOUT : bl_0_444 
* INOUT : br_0_444 
* INOUT : bl_0_445 
* INOUT : br_0_445 
* INOUT : bl_0_446 
* INOUT : br_0_446 
* INOUT : bl_0_447 
* INOUT : br_0_447 
* INOUT : bl_0_448 
* INOUT : br_0_448 
* INOUT : bl_0_449 
* INOUT : br_0_449 
* INOUT : bl_0_450 
* INOUT : br_0_450 
* INOUT : bl_0_451 
* INOUT : br_0_451 
* INOUT : bl_0_452 
* INOUT : br_0_452 
* INOUT : bl_0_453 
* INOUT : br_0_453 
* INOUT : bl_0_454 
* INOUT : br_0_454 
* INOUT : bl_0_455 
* INOUT : br_0_455 
* INOUT : bl_0_456 
* INOUT : br_0_456 
* INOUT : bl_0_457 
* INOUT : br_0_457 
* INOUT : bl_0_458 
* INOUT : br_0_458 
* INOUT : bl_0_459 
* INOUT : br_0_459 
* INOUT : bl_0_460 
* INOUT : br_0_460 
* INOUT : bl_0_461 
* INOUT : br_0_461 
* INOUT : bl_0_462 
* INOUT : br_0_462 
* INOUT : bl_0_463 
* INOUT : br_0_463 
* INOUT : bl_0_464 
* INOUT : br_0_464 
* INOUT : bl_0_465 
* INOUT : br_0_465 
* INOUT : bl_0_466 
* INOUT : br_0_466 
* INOUT : bl_0_467 
* INOUT : br_0_467 
* INOUT : bl_0_468 
* INOUT : br_0_468 
* INOUT : bl_0_469 
* INOUT : br_0_469 
* INOUT : bl_0_470 
* INOUT : br_0_470 
* INOUT : bl_0_471 
* INOUT : br_0_471 
* INOUT : bl_0_472 
* INOUT : br_0_472 
* INOUT : bl_0_473 
* INOUT : br_0_473 
* INOUT : bl_0_474 
* INOUT : br_0_474 
* INOUT : bl_0_475 
* INOUT : br_0_475 
* INOUT : bl_0_476 
* INOUT : br_0_476 
* INOUT : bl_0_477 
* INOUT : br_0_477 
* INOUT : bl_0_478 
* INOUT : br_0_478 
* INOUT : bl_0_479 
* INOUT : br_0_479 
* INOUT : bl_0_480 
* INOUT : br_0_480 
* INOUT : bl_0_481 
* INOUT : br_0_481 
* INOUT : bl_0_482 
* INOUT : br_0_482 
* INOUT : bl_0_483 
* INOUT : br_0_483 
* INOUT : bl_0_484 
* INOUT : br_0_484 
* INOUT : bl_0_485 
* INOUT : br_0_485 
* INOUT : bl_0_486 
* INOUT : br_0_486 
* INOUT : bl_0_487 
* INOUT : br_0_487 
* INOUT : bl_0_488 
* INOUT : br_0_488 
* INOUT : bl_0_489 
* INOUT : br_0_489 
* INOUT : bl_0_490 
* INOUT : br_0_490 
* INOUT : bl_0_491 
* INOUT : br_0_491 
* INOUT : bl_0_492 
* INOUT : br_0_492 
* INOUT : bl_0_493 
* INOUT : br_0_493 
* INOUT : bl_0_494 
* INOUT : br_0_494 
* INOUT : bl_0_495 
* INOUT : br_0_495 
* INOUT : bl_0_496 
* INOUT : br_0_496 
* INOUT : bl_0_497 
* INOUT : br_0_497 
* INOUT : bl_0_498 
* INOUT : br_0_498 
* INOUT : bl_0_499 
* INOUT : br_0_499 
* INOUT : bl_0_500 
* INOUT : br_0_500 
* INOUT : bl_0_501 
* INOUT : br_0_501 
* INOUT : bl_0_502 
* INOUT : br_0_502 
* INOUT : bl_0_503 
* INOUT : br_0_503 
* INOUT : bl_0_504 
* INOUT : br_0_504 
* INOUT : bl_0_505 
* INOUT : br_0_505 
* INOUT : bl_0_506 
* INOUT : br_0_506 
* INOUT : bl_0_507 
* INOUT : br_0_507 
* INOUT : bl_0_508 
* INOUT : br_0_508 
* INOUT : bl_0_509 
* INOUT : br_0_509 
* INOUT : bl_0_510 
* INOUT : br_0_510 
* INOUT : bl_0_511 
* INOUT : br_0_511 
* INOUT : bl_0_512 
* INOUT : br_0_512 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c256
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c257
+ bl_0_257 br_0_257 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c258
+ bl_0_258 br_0_258 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c259
+ bl_0_259 br_0_259 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c260
+ bl_0_260 br_0_260 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c261
+ bl_0_261 br_0_261 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c262
+ bl_0_262 br_0_262 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c263
+ bl_0_263 br_0_263 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c264
+ bl_0_264 br_0_264 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c265
+ bl_0_265 br_0_265 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c266
+ bl_0_266 br_0_266 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c267
+ bl_0_267 br_0_267 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c268
+ bl_0_268 br_0_268 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c269
+ bl_0_269 br_0_269 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c270
+ bl_0_270 br_0_270 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c271
+ bl_0_271 br_0_271 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c272
+ bl_0_272 br_0_272 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c273
+ bl_0_273 br_0_273 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c274
+ bl_0_274 br_0_274 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c275
+ bl_0_275 br_0_275 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c276
+ bl_0_276 br_0_276 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c277
+ bl_0_277 br_0_277 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c278
+ bl_0_278 br_0_278 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c279
+ bl_0_279 br_0_279 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c280
+ bl_0_280 br_0_280 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c281
+ bl_0_281 br_0_281 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c282
+ bl_0_282 br_0_282 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c283
+ bl_0_283 br_0_283 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c284
+ bl_0_284 br_0_284 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c285
+ bl_0_285 br_0_285 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c286
+ bl_0_286 br_0_286 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c287
+ bl_0_287 br_0_287 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c288
+ bl_0_288 br_0_288 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c289
+ bl_0_289 br_0_289 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c290
+ bl_0_290 br_0_290 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c291
+ bl_0_291 br_0_291 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c292
+ bl_0_292 br_0_292 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c293
+ bl_0_293 br_0_293 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c294
+ bl_0_294 br_0_294 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c295
+ bl_0_295 br_0_295 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c296
+ bl_0_296 br_0_296 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c297
+ bl_0_297 br_0_297 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c298
+ bl_0_298 br_0_298 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c299
+ bl_0_299 br_0_299 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c300
+ bl_0_300 br_0_300 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c301
+ bl_0_301 br_0_301 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c302
+ bl_0_302 br_0_302 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c303
+ bl_0_303 br_0_303 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c304
+ bl_0_304 br_0_304 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c305
+ bl_0_305 br_0_305 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c306
+ bl_0_306 br_0_306 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c307
+ bl_0_307 br_0_307 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c308
+ bl_0_308 br_0_308 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c309
+ bl_0_309 br_0_309 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c310
+ bl_0_310 br_0_310 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c311
+ bl_0_311 br_0_311 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c312
+ bl_0_312 br_0_312 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c313
+ bl_0_313 br_0_313 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c314
+ bl_0_314 br_0_314 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c315
+ bl_0_315 br_0_315 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c316
+ bl_0_316 br_0_316 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c317
+ bl_0_317 br_0_317 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c318
+ bl_0_318 br_0_318 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c319
+ bl_0_319 br_0_319 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c320
+ bl_0_320 br_0_320 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c321
+ bl_0_321 br_0_321 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c322
+ bl_0_322 br_0_322 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c323
+ bl_0_323 br_0_323 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c324
+ bl_0_324 br_0_324 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c325
+ bl_0_325 br_0_325 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c326
+ bl_0_326 br_0_326 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c327
+ bl_0_327 br_0_327 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c328
+ bl_0_328 br_0_328 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c329
+ bl_0_329 br_0_329 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c330
+ bl_0_330 br_0_330 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c331
+ bl_0_331 br_0_331 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c332
+ bl_0_332 br_0_332 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c333
+ bl_0_333 br_0_333 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c334
+ bl_0_334 br_0_334 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c335
+ bl_0_335 br_0_335 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c336
+ bl_0_336 br_0_336 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c337
+ bl_0_337 br_0_337 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c338
+ bl_0_338 br_0_338 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c339
+ bl_0_339 br_0_339 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c340
+ bl_0_340 br_0_340 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c341
+ bl_0_341 br_0_341 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c342
+ bl_0_342 br_0_342 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c343
+ bl_0_343 br_0_343 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c344
+ bl_0_344 br_0_344 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c345
+ bl_0_345 br_0_345 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c346
+ bl_0_346 br_0_346 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c347
+ bl_0_347 br_0_347 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c348
+ bl_0_348 br_0_348 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c349
+ bl_0_349 br_0_349 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c350
+ bl_0_350 br_0_350 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c351
+ bl_0_351 br_0_351 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c352
+ bl_0_352 br_0_352 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c353
+ bl_0_353 br_0_353 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c354
+ bl_0_354 br_0_354 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c355
+ bl_0_355 br_0_355 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c356
+ bl_0_356 br_0_356 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c357
+ bl_0_357 br_0_357 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c358
+ bl_0_358 br_0_358 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c359
+ bl_0_359 br_0_359 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c360
+ bl_0_360 br_0_360 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c361
+ bl_0_361 br_0_361 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c362
+ bl_0_362 br_0_362 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c363
+ bl_0_363 br_0_363 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c364
+ bl_0_364 br_0_364 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c365
+ bl_0_365 br_0_365 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c366
+ bl_0_366 br_0_366 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c367
+ bl_0_367 br_0_367 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c368
+ bl_0_368 br_0_368 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c369
+ bl_0_369 br_0_369 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c370
+ bl_0_370 br_0_370 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c371
+ bl_0_371 br_0_371 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c372
+ bl_0_372 br_0_372 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c373
+ bl_0_373 br_0_373 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c374
+ bl_0_374 br_0_374 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c375
+ bl_0_375 br_0_375 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c376
+ bl_0_376 br_0_376 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c377
+ bl_0_377 br_0_377 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c378
+ bl_0_378 br_0_378 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c379
+ bl_0_379 br_0_379 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c380
+ bl_0_380 br_0_380 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c381
+ bl_0_381 br_0_381 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c382
+ bl_0_382 br_0_382 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c383
+ bl_0_383 br_0_383 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c384
+ bl_0_384 br_0_384 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c385
+ bl_0_385 br_0_385 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c386
+ bl_0_386 br_0_386 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c387
+ bl_0_387 br_0_387 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c388
+ bl_0_388 br_0_388 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c389
+ bl_0_389 br_0_389 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c390
+ bl_0_390 br_0_390 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c391
+ bl_0_391 br_0_391 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c392
+ bl_0_392 br_0_392 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c393
+ bl_0_393 br_0_393 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c394
+ bl_0_394 br_0_394 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c395
+ bl_0_395 br_0_395 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c396
+ bl_0_396 br_0_396 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c397
+ bl_0_397 br_0_397 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c398
+ bl_0_398 br_0_398 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c399
+ bl_0_399 br_0_399 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c400
+ bl_0_400 br_0_400 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c401
+ bl_0_401 br_0_401 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c402
+ bl_0_402 br_0_402 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c403
+ bl_0_403 br_0_403 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c404
+ bl_0_404 br_0_404 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c405
+ bl_0_405 br_0_405 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c406
+ bl_0_406 br_0_406 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c407
+ bl_0_407 br_0_407 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c408
+ bl_0_408 br_0_408 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c409
+ bl_0_409 br_0_409 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c410
+ bl_0_410 br_0_410 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c411
+ bl_0_411 br_0_411 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c412
+ bl_0_412 br_0_412 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c413
+ bl_0_413 br_0_413 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c414
+ bl_0_414 br_0_414 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c415
+ bl_0_415 br_0_415 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c416
+ bl_0_416 br_0_416 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c417
+ bl_0_417 br_0_417 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c418
+ bl_0_418 br_0_418 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c419
+ bl_0_419 br_0_419 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c420
+ bl_0_420 br_0_420 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c421
+ bl_0_421 br_0_421 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c422
+ bl_0_422 br_0_422 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c423
+ bl_0_423 br_0_423 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c424
+ bl_0_424 br_0_424 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c425
+ bl_0_425 br_0_425 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c426
+ bl_0_426 br_0_426 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c427
+ bl_0_427 br_0_427 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c428
+ bl_0_428 br_0_428 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c429
+ bl_0_429 br_0_429 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c430
+ bl_0_430 br_0_430 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c431
+ bl_0_431 br_0_431 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c432
+ bl_0_432 br_0_432 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c433
+ bl_0_433 br_0_433 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c434
+ bl_0_434 br_0_434 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c435
+ bl_0_435 br_0_435 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c436
+ bl_0_436 br_0_436 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c437
+ bl_0_437 br_0_437 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c438
+ bl_0_438 br_0_438 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c439
+ bl_0_439 br_0_439 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c440
+ bl_0_440 br_0_440 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c441
+ bl_0_441 br_0_441 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c442
+ bl_0_442 br_0_442 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c443
+ bl_0_443 br_0_443 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c444
+ bl_0_444 br_0_444 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c445
+ bl_0_445 br_0_445 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c446
+ bl_0_446 br_0_446 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c447
+ bl_0_447 br_0_447 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c448
+ bl_0_448 br_0_448 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c449
+ bl_0_449 br_0_449 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c450
+ bl_0_450 br_0_450 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c451
+ bl_0_451 br_0_451 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c452
+ bl_0_452 br_0_452 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c453
+ bl_0_453 br_0_453 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c454
+ bl_0_454 br_0_454 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c455
+ bl_0_455 br_0_455 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c456
+ bl_0_456 br_0_456 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c457
+ bl_0_457 br_0_457 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c458
+ bl_0_458 br_0_458 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c459
+ bl_0_459 br_0_459 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c460
+ bl_0_460 br_0_460 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c461
+ bl_0_461 br_0_461 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c462
+ bl_0_462 br_0_462 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c463
+ bl_0_463 br_0_463 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c464
+ bl_0_464 br_0_464 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c465
+ bl_0_465 br_0_465 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c466
+ bl_0_466 br_0_466 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c467
+ bl_0_467 br_0_467 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c468
+ bl_0_468 br_0_468 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c469
+ bl_0_469 br_0_469 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c470
+ bl_0_470 br_0_470 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c471
+ bl_0_471 br_0_471 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c472
+ bl_0_472 br_0_472 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c473
+ bl_0_473 br_0_473 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c474
+ bl_0_474 br_0_474 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c475
+ bl_0_475 br_0_475 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c476
+ bl_0_476 br_0_476 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c477
+ bl_0_477 br_0_477 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c478
+ bl_0_478 br_0_478 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c479
+ bl_0_479 br_0_479 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c480
+ bl_0_480 br_0_480 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c481
+ bl_0_481 br_0_481 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c482
+ bl_0_482 br_0_482 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c483
+ bl_0_483 br_0_483 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c484
+ bl_0_484 br_0_484 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c485
+ bl_0_485 br_0_485 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c486
+ bl_0_486 br_0_486 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c487
+ bl_0_487 br_0_487 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c488
+ bl_0_488 br_0_488 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c489
+ bl_0_489 br_0_489 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c490
+ bl_0_490 br_0_490 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c491
+ bl_0_491 br_0_491 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c492
+ bl_0_492 br_0_492 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c493
+ bl_0_493 br_0_493 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c494
+ bl_0_494 br_0_494 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c495
+ bl_0_495 br_0_495 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c496
+ bl_0_496 br_0_496 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c497
+ bl_0_497 br_0_497 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c498
+ bl_0_498 br_0_498 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c499
+ bl_0_499 br_0_499 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c500
+ bl_0_500 br_0_500 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c501
+ bl_0_501 br_0_501 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c502
+ bl_0_502 br_0_502 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c503
+ bl_0_503 br_0_503 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c504
+ bl_0_504 br_0_504 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c505
+ bl_0_505 br_0_505 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c506
+ bl_0_506 br_0_506 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c507
+ bl_0_507 br_0_507 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c508
+ bl_0_508 br_0_508 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c509
+ bl_0_509 br_0_509 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c510
+ bl_0_510 br_0_510 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c511
+ bl_0_511 br_0_511 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c512
+ bl_0_512 br_0_512 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS freepdk45_sram_1rw0r_45x512_dummy_array_0

.SUBCKT freepdk45_sram_1rw0r_45x512_dummy_array_3
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ dummy_cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ dummy_cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ dummy_cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ dummy_cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ dummy_cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ dummy_cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ dummy_cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ dummy_cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ dummy_cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ dummy_cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ dummy_cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ dummy_cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ dummy_cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ dummy_cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ dummy_cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ dummy_cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ dummy_cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ dummy_cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ dummy_cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ dummy_cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ dummy_cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ dummy_cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ dummy_cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ dummy_cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ dummy_cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ dummy_cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ dummy_cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ dummy_cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ dummy_cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ dummy_cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ dummy_cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ dummy_cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ dummy_cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ dummy_cell_1rw
Xbit_r35_c0
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ dummy_cell_1rw
Xbit_r36_c0
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ dummy_cell_1rw
Xbit_r37_c0
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ dummy_cell_1rw
Xbit_r38_c0
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ dummy_cell_1rw
Xbit_r39_c0
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ dummy_cell_1rw
Xbit_r40_c0
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ dummy_cell_1rw
Xbit_r41_c0
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ dummy_cell_1rw
Xbit_r42_c0
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ dummy_cell_1rw
Xbit_r43_c0
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ dummy_cell_1rw
Xbit_r44_c0
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ dummy_cell_1rw
Xbit_r45_c0
+ bl_0_0 br_0_0 wl_0_45 vdd gnd
+ dummy_cell_1rw
Xbit_r46_c0
+ bl_0_0 br_0_0 wl_0_46 vdd gnd
+ dummy_cell_1rw
Xbit_r47_c0
+ bl_0_0 br_0_0 wl_0_47 vdd gnd
+ dummy_cell_1rw
.ENDS freepdk45_sram_1rw0r_45x512_dummy_array_3

.SUBCKT freepdk45_sram_1rw0r_45x512_capped_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258
+ br_0_258 bl_0_259 br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261
+ bl_0_262 br_0_262 bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265
+ br_0_265 bl_0_266 br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268
+ bl_0_269 br_0_269 bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272
+ br_0_272 bl_0_273 br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275
+ bl_0_276 br_0_276 bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279
+ br_0_279 bl_0_280 br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282
+ bl_0_283 br_0_283 bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286
+ br_0_286 bl_0_287 br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289
+ bl_0_290 br_0_290 bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293
+ br_0_293 bl_0_294 br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296
+ bl_0_297 br_0_297 bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300
+ br_0_300 bl_0_301 br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303
+ bl_0_304 br_0_304 bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307
+ br_0_307 bl_0_308 br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310
+ bl_0_311 br_0_311 bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314
+ br_0_314 bl_0_315 br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317
+ bl_0_318 br_0_318 bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321
+ br_0_321 bl_0_322 br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324
+ bl_0_325 br_0_325 bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328
+ br_0_328 bl_0_329 br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331
+ bl_0_332 br_0_332 bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335
+ br_0_335 bl_0_336 br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338
+ bl_0_339 br_0_339 bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342
+ br_0_342 bl_0_343 br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345
+ bl_0_346 br_0_346 bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349
+ br_0_349 bl_0_350 br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352
+ bl_0_353 br_0_353 bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356
+ br_0_356 bl_0_357 br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359
+ bl_0_360 br_0_360 bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363
+ br_0_363 bl_0_364 br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366
+ bl_0_367 br_0_367 bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370
+ br_0_370 bl_0_371 br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373
+ bl_0_374 br_0_374 bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377
+ br_0_377 bl_0_378 br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380
+ bl_0_381 br_0_381 bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384
+ br_0_384 bl_0_385 br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387
+ bl_0_388 br_0_388 bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391
+ br_0_391 bl_0_392 br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394
+ bl_0_395 br_0_395 bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398
+ br_0_398 bl_0_399 br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401
+ bl_0_402 br_0_402 bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405
+ br_0_405 bl_0_406 br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408
+ bl_0_409 br_0_409 bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412
+ br_0_412 bl_0_413 br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415
+ bl_0_416 br_0_416 bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419
+ br_0_419 bl_0_420 br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422
+ bl_0_423 br_0_423 bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426
+ br_0_426 bl_0_427 br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429
+ bl_0_430 br_0_430 bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433
+ br_0_433 bl_0_434 br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436
+ bl_0_437 br_0_437 bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440
+ br_0_440 bl_0_441 br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443
+ bl_0_444 br_0_444 bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447
+ br_0_447 bl_0_448 br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450
+ bl_0_451 br_0_451 bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454
+ br_0_454 bl_0_455 br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457
+ bl_0_458 br_0_458 bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461
+ br_0_461 bl_0_462 br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464
+ bl_0_465 br_0_465 bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468
+ br_0_468 bl_0_469 br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471
+ bl_0_472 br_0_472 bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475
+ br_0_475 bl_0_476 br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478
+ bl_0_479 br_0_479 bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482
+ br_0_482 bl_0_483 br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485
+ bl_0_486 br_0_486 bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489
+ br_0_489 bl_0_490 br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492
+ bl_0_493 br_0_493 bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496
+ br_0_496 bl_0_497 br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499
+ bl_0_500 br_0_500 bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503
+ br_0_503 bl_0_504 br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506
+ bl_0_507 br_0_507 bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510
+ br_0_510 bl_0_511 br_0_511 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3
+ wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12
+ wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20
+ wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28
+ wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36
+ wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 vdd
+ gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INOUT : bl_0_257 
* INOUT : br_0_257 
* INOUT : bl_0_258 
* INOUT : br_0_258 
* INOUT : bl_0_259 
* INOUT : br_0_259 
* INOUT : bl_0_260 
* INOUT : br_0_260 
* INOUT : bl_0_261 
* INOUT : br_0_261 
* INOUT : bl_0_262 
* INOUT : br_0_262 
* INOUT : bl_0_263 
* INOUT : br_0_263 
* INOUT : bl_0_264 
* INOUT : br_0_264 
* INOUT : bl_0_265 
* INOUT : br_0_265 
* INOUT : bl_0_266 
* INOUT : br_0_266 
* INOUT : bl_0_267 
* INOUT : br_0_267 
* INOUT : bl_0_268 
* INOUT : br_0_268 
* INOUT : bl_0_269 
* INOUT : br_0_269 
* INOUT : bl_0_270 
* INOUT : br_0_270 
* INOUT : bl_0_271 
* INOUT : br_0_271 
* INOUT : bl_0_272 
* INOUT : br_0_272 
* INOUT : bl_0_273 
* INOUT : br_0_273 
* INOUT : bl_0_274 
* INOUT : br_0_274 
* INOUT : bl_0_275 
* INOUT : br_0_275 
* INOUT : bl_0_276 
* INOUT : br_0_276 
* INOUT : bl_0_277 
* INOUT : br_0_277 
* INOUT : bl_0_278 
* INOUT : br_0_278 
* INOUT : bl_0_279 
* INOUT : br_0_279 
* INOUT : bl_0_280 
* INOUT : br_0_280 
* INOUT : bl_0_281 
* INOUT : br_0_281 
* INOUT : bl_0_282 
* INOUT : br_0_282 
* INOUT : bl_0_283 
* INOUT : br_0_283 
* INOUT : bl_0_284 
* INOUT : br_0_284 
* INOUT : bl_0_285 
* INOUT : br_0_285 
* INOUT : bl_0_286 
* INOUT : br_0_286 
* INOUT : bl_0_287 
* INOUT : br_0_287 
* INOUT : bl_0_288 
* INOUT : br_0_288 
* INOUT : bl_0_289 
* INOUT : br_0_289 
* INOUT : bl_0_290 
* INOUT : br_0_290 
* INOUT : bl_0_291 
* INOUT : br_0_291 
* INOUT : bl_0_292 
* INOUT : br_0_292 
* INOUT : bl_0_293 
* INOUT : br_0_293 
* INOUT : bl_0_294 
* INOUT : br_0_294 
* INOUT : bl_0_295 
* INOUT : br_0_295 
* INOUT : bl_0_296 
* INOUT : br_0_296 
* INOUT : bl_0_297 
* INOUT : br_0_297 
* INOUT : bl_0_298 
* INOUT : br_0_298 
* INOUT : bl_0_299 
* INOUT : br_0_299 
* INOUT : bl_0_300 
* INOUT : br_0_300 
* INOUT : bl_0_301 
* INOUT : br_0_301 
* INOUT : bl_0_302 
* INOUT : br_0_302 
* INOUT : bl_0_303 
* INOUT : br_0_303 
* INOUT : bl_0_304 
* INOUT : br_0_304 
* INOUT : bl_0_305 
* INOUT : br_0_305 
* INOUT : bl_0_306 
* INOUT : br_0_306 
* INOUT : bl_0_307 
* INOUT : br_0_307 
* INOUT : bl_0_308 
* INOUT : br_0_308 
* INOUT : bl_0_309 
* INOUT : br_0_309 
* INOUT : bl_0_310 
* INOUT : br_0_310 
* INOUT : bl_0_311 
* INOUT : br_0_311 
* INOUT : bl_0_312 
* INOUT : br_0_312 
* INOUT : bl_0_313 
* INOUT : br_0_313 
* INOUT : bl_0_314 
* INOUT : br_0_314 
* INOUT : bl_0_315 
* INOUT : br_0_315 
* INOUT : bl_0_316 
* INOUT : br_0_316 
* INOUT : bl_0_317 
* INOUT : br_0_317 
* INOUT : bl_0_318 
* INOUT : br_0_318 
* INOUT : bl_0_319 
* INOUT : br_0_319 
* INOUT : bl_0_320 
* INOUT : br_0_320 
* INOUT : bl_0_321 
* INOUT : br_0_321 
* INOUT : bl_0_322 
* INOUT : br_0_322 
* INOUT : bl_0_323 
* INOUT : br_0_323 
* INOUT : bl_0_324 
* INOUT : br_0_324 
* INOUT : bl_0_325 
* INOUT : br_0_325 
* INOUT : bl_0_326 
* INOUT : br_0_326 
* INOUT : bl_0_327 
* INOUT : br_0_327 
* INOUT : bl_0_328 
* INOUT : br_0_328 
* INOUT : bl_0_329 
* INOUT : br_0_329 
* INOUT : bl_0_330 
* INOUT : br_0_330 
* INOUT : bl_0_331 
* INOUT : br_0_331 
* INOUT : bl_0_332 
* INOUT : br_0_332 
* INOUT : bl_0_333 
* INOUT : br_0_333 
* INOUT : bl_0_334 
* INOUT : br_0_334 
* INOUT : bl_0_335 
* INOUT : br_0_335 
* INOUT : bl_0_336 
* INOUT : br_0_336 
* INOUT : bl_0_337 
* INOUT : br_0_337 
* INOUT : bl_0_338 
* INOUT : br_0_338 
* INOUT : bl_0_339 
* INOUT : br_0_339 
* INOUT : bl_0_340 
* INOUT : br_0_340 
* INOUT : bl_0_341 
* INOUT : br_0_341 
* INOUT : bl_0_342 
* INOUT : br_0_342 
* INOUT : bl_0_343 
* INOUT : br_0_343 
* INOUT : bl_0_344 
* INOUT : br_0_344 
* INOUT : bl_0_345 
* INOUT : br_0_345 
* INOUT : bl_0_346 
* INOUT : br_0_346 
* INOUT : bl_0_347 
* INOUT : br_0_347 
* INOUT : bl_0_348 
* INOUT : br_0_348 
* INOUT : bl_0_349 
* INOUT : br_0_349 
* INOUT : bl_0_350 
* INOUT : br_0_350 
* INOUT : bl_0_351 
* INOUT : br_0_351 
* INOUT : bl_0_352 
* INOUT : br_0_352 
* INOUT : bl_0_353 
* INOUT : br_0_353 
* INOUT : bl_0_354 
* INOUT : br_0_354 
* INOUT : bl_0_355 
* INOUT : br_0_355 
* INOUT : bl_0_356 
* INOUT : br_0_356 
* INOUT : bl_0_357 
* INOUT : br_0_357 
* INOUT : bl_0_358 
* INOUT : br_0_358 
* INOUT : bl_0_359 
* INOUT : br_0_359 
* INOUT : bl_0_360 
* INOUT : br_0_360 
* INOUT : bl_0_361 
* INOUT : br_0_361 
* INOUT : bl_0_362 
* INOUT : br_0_362 
* INOUT : bl_0_363 
* INOUT : br_0_363 
* INOUT : bl_0_364 
* INOUT : br_0_364 
* INOUT : bl_0_365 
* INOUT : br_0_365 
* INOUT : bl_0_366 
* INOUT : br_0_366 
* INOUT : bl_0_367 
* INOUT : br_0_367 
* INOUT : bl_0_368 
* INOUT : br_0_368 
* INOUT : bl_0_369 
* INOUT : br_0_369 
* INOUT : bl_0_370 
* INOUT : br_0_370 
* INOUT : bl_0_371 
* INOUT : br_0_371 
* INOUT : bl_0_372 
* INOUT : br_0_372 
* INOUT : bl_0_373 
* INOUT : br_0_373 
* INOUT : bl_0_374 
* INOUT : br_0_374 
* INOUT : bl_0_375 
* INOUT : br_0_375 
* INOUT : bl_0_376 
* INOUT : br_0_376 
* INOUT : bl_0_377 
* INOUT : br_0_377 
* INOUT : bl_0_378 
* INOUT : br_0_378 
* INOUT : bl_0_379 
* INOUT : br_0_379 
* INOUT : bl_0_380 
* INOUT : br_0_380 
* INOUT : bl_0_381 
* INOUT : br_0_381 
* INOUT : bl_0_382 
* INOUT : br_0_382 
* INOUT : bl_0_383 
* INOUT : br_0_383 
* INOUT : bl_0_384 
* INOUT : br_0_384 
* INOUT : bl_0_385 
* INOUT : br_0_385 
* INOUT : bl_0_386 
* INOUT : br_0_386 
* INOUT : bl_0_387 
* INOUT : br_0_387 
* INOUT : bl_0_388 
* INOUT : br_0_388 
* INOUT : bl_0_389 
* INOUT : br_0_389 
* INOUT : bl_0_390 
* INOUT : br_0_390 
* INOUT : bl_0_391 
* INOUT : br_0_391 
* INOUT : bl_0_392 
* INOUT : br_0_392 
* INOUT : bl_0_393 
* INOUT : br_0_393 
* INOUT : bl_0_394 
* INOUT : br_0_394 
* INOUT : bl_0_395 
* INOUT : br_0_395 
* INOUT : bl_0_396 
* INOUT : br_0_396 
* INOUT : bl_0_397 
* INOUT : br_0_397 
* INOUT : bl_0_398 
* INOUT : br_0_398 
* INOUT : bl_0_399 
* INOUT : br_0_399 
* INOUT : bl_0_400 
* INOUT : br_0_400 
* INOUT : bl_0_401 
* INOUT : br_0_401 
* INOUT : bl_0_402 
* INOUT : br_0_402 
* INOUT : bl_0_403 
* INOUT : br_0_403 
* INOUT : bl_0_404 
* INOUT : br_0_404 
* INOUT : bl_0_405 
* INOUT : br_0_405 
* INOUT : bl_0_406 
* INOUT : br_0_406 
* INOUT : bl_0_407 
* INOUT : br_0_407 
* INOUT : bl_0_408 
* INOUT : br_0_408 
* INOUT : bl_0_409 
* INOUT : br_0_409 
* INOUT : bl_0_410 
* INOUT : br_0_410 
* INOUT : bl_0_411 
* INOUT : br_0_411 
* INOUT : bl_0_412 
* INOUT : br_0_412 
* INOUT : bl_0_413 
* INOUT : br_0_413 
* INOUT : bl_0_414 
* INOUT : br_0_414 
* INOUT : bl_0_415 
* INOUT : br_0_415 
* INOUT : bl_0_416 
* INOUT : br_0_416 
* INOUT : bl_0_417 
* INOUT : br_0_417 
* INOUT : bl_0_418 
* INOUT : br_0_418 
* INOUT : bl_0_419 
* INOUT : br_0_419 
* INOUT : bl_0_420 
* INOUT : br_0_420 
* INOUT : bl_0_421 
* INOUT : br_0_421 
* INOUT : bl_0_422 
* INOUT : br_0_422 
* INOUT : bl_0_423 
* INOUT : br_0_423 
* INOUT : bl_0_424 
* INOUT : br_0_424 
* INOUT : bl_0_425 
* INOUT : br_0_425 
* INOUT : bl_0_426 
* INOUT : br_0_426 
* INOUT : bl_0_427 
* INOUT : br_0_427 
* INOUT : bl_0_428 
* INOUT : br_0_428 
* INOUT : bl_0_429 
* INOUT : br_0_429 
* INOUT : bl_0_430 
* INOUT : br_0_430 
* INOUT : bl_0_431 
* INOUT : br_0_431 
* INOUT : bl_0_432 
* INOUT : br_0_432 
* INOUT : bl_0_433 
* INOUT : br_0_433 
* INOUT : bl_0_434 
* INOUT : br_0_434 
* INOUT : bl_0_435 
* INOUT : br_0_435 
* INOUT : bl_0_436 
* INOUT : br_0_436 
* INOUT : bl_0_437 
* INOUT : br_0_437 
* INOUT : bl_0_438 
* INOUT : br_0_438 
* INOUT : bl_0_439 
* INOUT : br_0_439 
* INOUT : bl_0_440 
* INOUT : br_0_440 
* INOUT : bl_0_441 
* INOUT : br_0_441 
* INOUT : bl_0_442 
* INOUT : br_0_442 
* INOUT : bl_0_443 
* INOUT : br_0_443 
* INOUT : bl_0_444 
* INOUT : br_0_444 
* INOUT : bl_0_445 
* INOUT : br_0_445 
* INOUT : bl_0_446 
* INOUT : br_0_446 
* INOUT : bl_0_447 
* INOUT : br_0_447 
* INOUT : bl_0_448 
* INOUT : br_0_448 
* INOUT : bl_0_449 
* INOUT : br_0_449 
* INOUT : bl_0_450 
* INOUT : br_0_450 
* INOUT : bl_0_451 
* INOUT : br_0_451 
* INOUT : bl_0_452 
* INOUT : br_0_452 
* INOUT : bl_0_453 
* INOUT : br_0_453 
* INOUT : bl_0_454 
* INOUT : br_0_454 
* INOUT : bl_0_455 
* INOUT : br_0_455 
* INOUT : bl_0_456 
* INOUT : br_0_456 
* INOUT : bl_0_457 
* INOUT : br_0_457 
* INOUT : bl_0_458 
* INOUT : br_0_458 
* INOUT : bl_0_459 
* INOUT : br_0_459 
* INOUT : bl_0_460 
* INOUT : br_0_460 
* INOUT : bl_0_461 
* INOUT : br_0_461 
* INOUT : bl_0_462 
* INOUT : br_0_462 
* INOUT : bl_0_463 
* INOUT : br_0_463 
* INOUT : bl_0_464 
* INOUT : br_0_464 
* INOUT : bl_0_465 
* INOUT : br_0_465 
* INOUT : bl_0_466 
* INOUT : br_0_466 
* INOUT : bl_0_467 
* INOUT : br_0_467 
* INOUT : bl_0_468 
* INOUT : br_0_468 
* INOUT : bl_0_469 
* INOUT : br_0_469 
* INOUT : bl_0_470 
* INOUT : br_0_470 
* INOUT : bl_0_471 
* INOUT : br_0_471 
* INOUT : bl_0_472 
* INOUT : br_0_472 
* INOUT : bl_0_473 
* INOUT : br_0_473 
* INOUT : bl_0_474 
* INOUT : br_0_474 
* INOUT : bl_0_475 
* INOUT : br_0_475 
* INOUT : bl_0_476 
* INOUT : br_0_476 
* INOUT : bl_0_477 
* INOUT : br_0_477 
* INOUT : bl_0_478 
* INOUT : br_0_478 
* INOUT : bl_0_479 
* INOUT : br_0_479 
* INOUT : bl_0_480 
* INOUT : br_0_480 
* INOUT : bl_0_481 
* INOUT : br_0_481 
* INOUT : bl_0_482 
* INOUT : br_0_482 
* INOUT : bl_0_483 
* INOUT : br_0_483 
* INOUT : bl_0_484 
* INOUT : br_0_484 
* INOUT : bl_0_485 
* INOUT : br_0_485 
* INOUT : bl_0_486 
* INOUT : br_0_486 
* INOUT : bl_0_487 
* INOUT : br_0_487 
* INOUT : bl_0_488 
* INOUT : br_0_488 
* INOUT : bl_0_489 
* INOUT : br_0_489 
* INOUT : bl_0_490 
* INOUT : br_0_490 
* INOUT : bl_0_491 
* INOUT : br_0_491 
* INOUT : bl_0_492 
* INOUT : br_0_492 
* INOUT : bl_0_493 
* INOUT : br_0_493 
* INOUT : bl_0_494 
* INOUT : br_0_494 
* INOUT : bl_0_495 
* INOUT : br_0_495 
* INOUT : bl_0_496 
* INOUT : br_0_496 
* INOUT : bl_0_497 
* INOUT : br_0_497 
* INOUT : bl_0_498 
* INOUT : br_0_498 
* INOUT : bl_0_499 
* INOUT : br_0_499 
* INOUT : bl_0_500 
* INOUT : br_0_500 
* INOUT : bl_0_501 
* INOUT : br_0_501 
* INOUT : bl_0_502 
* INOUT : br_0_502 
* INOUT : bl_0_503 
* INOUT : br_0_503 
* INOUT : bl_0_504 
* INOUT : br_0_504 
* INOUT : bl_0_505 
* INOUT : br_0_505 
* INOUT : bl_0_506 
* INOUT : br_0_506 
* INOUT : bl_0_507 
* INOUT : br_0_507 
* INOUT : bl_0_508 
* INOUT : br_0_508 
* INOUT : bl_0_509 
* INOUT : br_0_509 
* INOUT : bl_0_510 
* INOUT : br_0_510 
* INOUT : bl_0_511 
* INOUT : br_0_511 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* POWER : vdd 
* GROUND: gnd 
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xreplica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258
+ br_0_258 bl_0_259 br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261
+ bl_0_262 br_0_262 bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265
+ br_0_265 bl_0_266 br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268
+ bl_0_269 br_0_269 bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272
+ br_0_272 bl_0_273 br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275
+ bl_0_276 br_0_276 bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279
+ br_0_279 bl_0_280 br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282
+ bl_0_283 br_0_283 bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286
+ br_0_286 bl_0_287 br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289
+ bl_0_290 br_0_290 bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293
+ br_0_293 bl_0_294 br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296
+ bl_0_297 br_0_297 bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300
+ br_0_300 bl_0_301 br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303
+ bl_0_304 br_0_304 bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307
+ br_0_307 bl_0_308 br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310
+ bl_0_311 br_0_311 bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314
+ br_0_314 bl_0_315 br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317
+ bl_0_318 br_0_318 bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321
+ br_0_321 bl_0_322 br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324
+ bl_0_325 br_0_325 bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328
+ br_0_328 bl_0_329 br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331
+ bl_0_332 br_0_332 bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335
+ br_0_335 bl_0_336 br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338
+ bl_0_339 br_0_339 bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342
+ br_0_342 bl_0_343 br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345
+ bl_0_346 br_0_346 bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349
+ br_0_349 bl_0_350 br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352
+ bl_0_353 br_0_353 bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356
+ br_0_356 bl_0_357 br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359
+ bl_0_360 br_0_360 bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363
+ br_0_363 bl_0_364 br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366
+ bl_0_367 br_0_367 bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370
+ br_0_370 bl_0_371 br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373
+ bl_0_374 br_0_374 bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377
+ br_0_377 bl_0_378 br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380
+ bl_0_381 br_0_381 bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384
+ br_0_384 bl_0_385 br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387
+ bl_0_388 br_0_388 bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391
+ br_0_391 bl_0_392 br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394
+ bl_0_395 br_0_395 bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398
+ br_0_398 bl_0_399 br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401
+ bl_0_402 br_0_402 bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405
+ br_0_405 bl_0_406 br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408
+ bl_0_409 br_0_409 bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412
+ br_0_412 bl_0_413 br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415
+ bl_0_416 br_0_416 bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419
+ br_0_419 bl_0_420 br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422
+ bl_0_423 br_0_423 bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426
+ br_0_426 bl_0_427 br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429
+ bl_0_430 br_0_430 bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433
+ br_0_433 bl_0_434 br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436
+ bl_0_437 br_0_437 bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440
+ br_0_440 bl_0_441 br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443
+ bl_0_444 br_0_444 bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447
+ br_0_447 bl_0_448 br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450
+ bl_0_451 br_0_451 bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454
+ br_0_454 bl_0_455 br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457
+ bl_0_458 br_0_458 bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461
+ br_0_461 bl_0_462 br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464
+ bl_0_465 br_0_465 bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468
+ br_0_468 bl_0_469 br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471
+ bl_0_472 br_0_472 bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475
+ br_0_475 bl_0_476 br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478
+ bl_0_479 br_0_479 bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482
+ br_0_482 bl_0_483 br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485
+ bl_0_486 br_0_486 bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489
+ br_0_489 bl_0_490 br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492
+ bl_0_493 br_0_493 bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496
+ br_0_496 bl_0_497 br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499
+ bl_0_500 br_0_500 bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503
+ br_0_503 bl_0_504 br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506
+ bl_0_507 br_0_507 bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510
+ br_0_510 bl_0_511 br_0_511 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3
+ wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12
+ wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20
+ wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28
+ wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36
+ wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 vdd
+ gnd
+ freepdk45_sram_1rw0r_45x512_replica_bitcell_array
Xdummy_row_bot
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258
+ br_0_258 bl_0_259 br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261
+ bl_0_262 br_0_262 bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265
+ br_0_265 bl_0_266 br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268
+ bl_0_269 br_0_269 bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272
+ br_0_272 bl_0_273 br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275
+ bl_0_276 br_0_276 bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279
+ br_0_279 bl_0_280 br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282
+ bl_0_283 br_0_283 bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286
+ br_0_286 bl_0_287 br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289
+ bl_0_290 br_0_290 bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293
+ br_0_293 bl_0_294 br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296
+ bl_0_297 br_0_297 bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300
+ br_0_300 bl_0_301 br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303
+ bl_0_304 br_0_304 bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307
+ br_0_307 bl_0_308 br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310
+ bl_0_311 br_0_311 bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314
+ br_0_314 bl_0_315 br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317
+ bl_0_318 br_0_318 bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321
+ br_0_321 bl_0_322 br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324
+ bl_0_325 br_0_325 bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328
+ br_0_328 bl_0_329 br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331
+ bl_0_332 br_0_332 bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335
+ br_0_335 bl_0_336 br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338
+ bl_0_339 br_0_339 bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342
+ br_0_342 bl_0_343 br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345
+ bl_0_346 br_0_346 bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349
+ br_0_349 bl_0_350 br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352
+ bl_0_353 br_0_353 bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356
+ br_0_356 bl_0_357 br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359
+ bl_0_360 br_0_360 bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363
+ br_0_363 bl_0_364 br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366
+ bl_0_367 br_0_367 bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370
+ br_0_370 bl_0_371 br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373
+ bl_0_374 br_0_374 bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377
+ br_0_377 bl_0_378 br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380
+ bl_0_381 br_0_381 bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384
+ br_0_384 bl_0_385 br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387
+ bl_0_388 br_0_388 bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391
+ br_0_391 bl_0_392 br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394
+ bl_0_395 br_0_395 bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398
+ br_0_398 bl_0_399 br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401
+ bl_0_402 br_0_402 bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405
+ br_0_405 bl_0_406 br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408
+ bl_0_409 br_0_409 bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412
+ br_0_412 bl_0_413 br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415
+ bl_0_416 br_0_416 bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419
+ br_0_419 bl_0_420 br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422
+ bl_0_423 br_0_423 bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426
+ br_0_426 bl_0_427 br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429
+ bl_0_430 br_0_430 bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433
+ br_0_433 bl_0_434 br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436
+ bl_0_437 br_0_437 bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440
+ br_0_440 bl_0_441 br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443
+ bl_0_444 br_0_444 bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447
+ br_0_447 bl_0_448 br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450
+ bl_0_451 br_0_451 bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454
+ br_0_454 bl_0_455 br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457
+ bl_0_458 br_0_458 bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461
+ br_0_461 bl_0_462 br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464
+ bl_0_465 br_0_465 bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468
+ br_0_468 bl_0_469 br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471
+ bl_0_472 br_0_472 bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475
+ br_0_475 bl_0_476 br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478
+ bl_0_479 br_0_479 bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482
+ br_0_482 bl_0_483 br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485
+ bl_0_486 br_0_486 bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489
+ br_0_489 bl_0_490 br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492
+ bl_0_493 br_0_493 bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496
+ br_0_496 bl_0_497 br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499
+ bl_0_500 br_0_500 bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503
+ br_0_503 bl_0_504 br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506
+ bl_0_507 br_0_507 bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510
+ br_0_510 bl_0_511 br_0_511 gnd vdd gnd
+ freepdk45_sram_1rw0r_45x512_dummy_array_1
Xdummy_row_top
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258
+ br_0_258 bl_0_259 br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261
+ bl_0_262 br_0_262 bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265
+ br_0_265 bl_0_266 br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268
+ bl_0_269 br_0_269 bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272
+ br_0_272 bl_0_273 br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275
+ bl_0_276 br_0_276 bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279
+ br_0_279 bl_0_280 br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282
+ bl_0_283 br_0_283 bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286
+ br_0_286 bl_0_287 br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289
+ bl_0_290 br_0_290 bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293
+ br_0_293 bl_0_294 br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296
+ bl_0_297 br_0_297 bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300
+ br_0_300 bl_0_301 br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303
+ bl_0_304 br_0_304 bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307
+ br_0_307 bl_0_308 br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310
+ bl_0_311 br_0_311 bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314
+ br_0_314 bl_0_315 br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317
+ bl_0_318 br_0_318 bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321
+ br_0_321 bl_0_322 br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324
+ bl_0_325 br_0_325 bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328
+ br_0_328 bl_0_329 br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331
+ bl_0_332 br_0_332 bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335
+ br_0_335 bl_0_336 br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338
+ bl_0_339 br_0_339 bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342
+ br_0_342 bl_0_343 br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345
+ bl_0_346 br_0_346 bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349
+ br_0_349 bl_0_350 br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352
+ bl_0_353 br_0_353 bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356
+ br_0_356 bl_0_357 br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359
+ bl_0_360 br_0_360 bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363
+ br_0_363 bl_0_364 br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366
+ bl_0_367 br_0_367 bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370
+ br_0_370 bl_0_371 br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373
+ bl_0_374 br_0_374 bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377
+ br_0_377 bl_0_378 br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380
+ bl_0_381 br_0_381 bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384
+ br_0_384 bl_0_385 br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387
+ bl_0_388 br_0_388 bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391
+ br_0_391 bl_0_392 br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394
+ bl_0_395 br_0_395 bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398
+ br_0_398 bl_0_399 br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401
+ bl_0_402 br_0_402 bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405
+ br_0_405 bl_0_406 br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408
+ bl_0_409 br_0_409 bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412
+ br_0_412 bl_0_413 br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415
+ bl_0_416 br_0_416 bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419
+ br_0_419 bl_0_420 br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422
+ bl_0_423 br_0_423 bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426
+ br_0_426 bl_0_427 br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429
+ bl_0_430 br_0_430 bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433
+ br_0_433 bl_0_434 br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436
+ bl_0_437 br_0_437 bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440
+ br_0_440 bl_0_441 br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443
+ bl_0_444 br_0_444 bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447
+ br_0_447 bl_0_448 br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450
+ bl_0_451 br_0_451 bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454
+ br_0_454 bl_0_455 br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457
+ bl_0_458 br_0_458 bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461
+ br_0_461 bl_0_462 br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464
+ bl_0_465 br_0_465 bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468
+ br_0_468 bl_0_469 br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471
+ bl_0_472 br_0_472 bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475
+ br_0_475 bl_0_476 br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478
+ bl_0_479 br_0_479 bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482
+ br_0_482 bl_0_483 br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485
+ bl_0_486 br_0_486 bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489
+ br_0_489 bl_0_490 br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492
+ bl_0_493 br_0_493 bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496
+ br_0_496 bl_0_497 br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499
+ bl_0_500 br_0_500 bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503
+ br_0_503 bl_0_504 br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506
+ bl_0_507 br_0_507 bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510
+ br_0_510 bl_0_511 br_0_511 gnd vdd gnd
+ freepdk45_sram_1rw0r_45x512_dummy_array_0
Xdummy_col_left
+ dummy_left_bl_0_0 dummy_left_br_0_0 gnd rbl_wl_0_0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 gnd vdd gnd
+ freepdk45_sram_1rw0r_45x512_dummy_array_2
Xdummy_col_right
+ dummy_right_bl_0_0 dummy_right_br_0_0 gnd rbl_wl_0_0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 gnd vdd gnd
+ freepdk45_sram_1rw0r_45x512_dummy_array_3
.ENDS freepdk45_sram_1rw0r_45x512_capped_replica_bitcell_array

.SUBCKT freepdk45_sram_1rw0r_45x512_bank
+ dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7
+ dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15
+ dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22
+ dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29
+ dout0_30 dout0_31 dout0_32 dout0_33 dout0_34 dout0_35 dout0_36
+ dout0_37 dout0_38 dout0_39 dout0_40 dout0_41 dout0_42 dout0_43
+ dout0_44 dout0_45 dout0_46 dout0_47 dout0_48 dout0_49 dout0_50
+ dout0_51 dout0_52 dout0_53 dout0_54 dout0_55 dout0_56 dout0_57
+ dout0_58 dout0_59 dout0_60 dout0_61 dout0_62 dout0_63 dout0_64
+ dout0_65 dout0_66 dout0_67 dout0_68 dout0_69 dout0_70 dout0_71
+ dout0_72 dout0_73 dout0_74 dout0_75 dout0_76 dout0_77 dout0_78
+ dout0_79 dout0_80 dout0_81 dout0_82 dout0_83 dout0_84 dout0_85
+ dout0_86 dout0_87 dout0_88 dout0_89 dout0_90 dout0_91 dout0_92
+ dout0_93 dout0_94 dout0_95 dout0_96 dout0_97 dout0_98 dout0_99
+ dout0_100 dout0_101 dout0_102 dout0_103 dout0_104 dout0_105 dout0_106
+ dout0_107 dout0_108 dout0_109 dout0_110 dout0_111 dout0_112 dout0_113
+ dout0_114 dout0_115 dout0_116 dout0_117 dout0_118 dout0_119 dout0_120
+ dout0_121 dout0_122 dout0_123 dout0_124 dout0_125 dout0_126 dout0_127
+ dout0_128 dout0_129 dout0_130 dout0_131 dout0_132 dout0_133 dout0_134
+ dout0_135 dout0_136 dout0_137 dout0_138 dout0_139 dout0_140 dout0_141
+ dout0_142 dout0_143 dout0_144 dout0_145 dout0_146 dout0_147 dout0_148
+ dout0_149 dout0_150 dout0_151 dout0_152 dout0_153 dout0_154 dout0_155
+ dout0_156 dout0_157 dout0_158 dout0_159 dout0_160 dout0_161 dout0_162
+ dout0_163 dout0_164 dout0_165 dout0_166 dout0_167 dout0_168 dout0_169
+ dout0_170 dout0_171 dout0_172 dout0_173 dout0_174 dout0_175 dout0_176
+ dout0_177 dout0_178 dout0_179 dout0_180 dout0_181 dout0_182 dout0_183
+ dout0_184 dout0_185 dout0_186 dout0_187 dout0_188 dout0_189 dout0_190
+ dout0_191 dout0_192 dout0_193 dout0_194 dout0_195 dout0_196 dout0_197
+ dout0_198 dout0_199 dout0_200 dout0_201 dout0_202 dout0_203 dout0_204
+ dout0_205 dout0_206 dout0_207 dout0_208 dout0_209 dout0_210 dout0_211
+ dout0_212 dout0_213 dout0_214 dout0_215 dout0_216 dout0_217 dout0_218
+ dout0_219 dout0_220 dout0_221 dout0_222 dout0_223 dout0_224 dout0_225
+ dout0_226 dout0_227 dout0_228 dout0_229 dout0_230 dout0_231 dout0_232
+ dout0_233 dout0_234 dout0_235 dout0_236 dout0_237 dout0_238 dout0_239
+ dout0_240 dout0_241 dout0_242 dout0_243 dout0_244 dout0_245 dout0_246
+ dout0_247 dout0_248 dout0_249 dout0_250 dout0_251 dout0_252 dout0_253
+ dout0_254 dout0_255 dout0_256 dout0_257 dout0_258 dout0_259 dout0_260
+ dout0_261 dout0_262 dout0_263 dout0_264 dout0_265 dout0_266 dout0_267
+ dout0_268 dout0_269 dout0_270 dout0_271 dout0_272 dout0_273 dout0_274
+ dout0_275 dout0_276 dout0_277 dout0_278 dout0_279 dout0_280 dout0_281
+ dout0_282 dout0_283 dout0_284 dout0_285 dout0_286 dout0_287 dout0_288
+ dout0_289 dout0_290 dout0_291 dout0_292 dout0_293 dout0_294 dout0_295
+ dout0_296 dout0_297 dout0_298 dout0_299 dout0_300 dout0_301 dout0_302
+ dout0_303 dout0_304 dout0_305 dout0_306 dout0_307 dout0_308 dout0_309
+ dout0_310 dout0_311 dout0_312 dout0_313 dout0_314 dout0_315 dout0_316
+ dout0_317 dout0_318 dout0_319 dout0_320 dout0_321 dout0_322 dout0_323
+ dout0_324 dout0_325 dout0_326 dout0_327 dout0_328 dout0_329 dout0_330
+ dout0_331 dout0_332 dout0_333 dout0_334 dout0_335 dout0_336 dout0_337
+ dout0_338 dout0_339 dout0_340 dout0_341 dout0_342 dout0_343 dout0_344
+ dout0_345 dout0_346 dout0_347 dout0_348 dout0_349 dout0_350 dout0_351
+ dout0_352 dout0_353 dout0_354 dout0_355 dout0_356 dout0_357 dout0_358
+ dout0_359 dout0_360 dout0_361 dout0_362 dout0_363 dout0_364 dout0_365
+ dout0_366 dout0_367 dout0_368 dout0_369 dout0_370 dout0_371 dout0_372
+ dout0_373 dout0_374 dout0_375 dout0_376 dout0_377 dout0_378 dout0_379
+ dout0_380 dout0_381 dout0_382 dout0_383 dout0_384 dout0_385 dout0_386
+ dout0_387 dout0_388 dout0_389 dout0_390 dout0_391 dout0_392 dout0_393
+ dout0_394 dout0_395 dout0_396 dout0_397 dout0_398 dout0_399 dout0_400
+ dout0_401 dout0_402 dout0_403 dout0_404 dout0_405 dout0_406 dout0_407
+ dout0_408 dout0_409 dout0_410 dout0_411 dout0_412 dout0_413 dout0_414
+ dout0_415 dout0_416 dout0_417 dout0_418 dout0_419 dout0_420 dout0_421
+ dout0_422 dout0_423 dout0_424 dout0_425 dout0_426 dout0_427 dout0_428
+ dout0_429 dout0_430 dout0_431 dout0_432 dout0_433 dout0_434 dout0_435
+ dout0_436 dout0_437 dout0_438 dout0_439 dout0_440 dout0_441 dout0_442
+ dout0_443 dout0_444 dout0_445 dout0_446 dout0_447 dout0_448 dout0_449
+ dout0_450 dout0_451 dout0_452 dout0_453 dout0_454 dout0_455 dout0_456
+ dout0_457 dout0_458 dout0_459 dout0_460 dout0_461 dout0_462 dout0_463
+ dout0_464 dout0_465 dout0_466 dout0_467 dout0_468 dout0_469 dout0_470
+ dout0_471 dout0_472 dout0_473 dout0_474 dout0_475 dout0_476 dout0_477
+ dout0_478 dout0_479 dout0_480 dout0_481 dout0_482 dout0_483 dout0_484
+ dout0_485 dout0_486 dout0_487 dout0_488 dout0_489 dout0_490 dout0_491
+ dout0_492 dout0_493 dout0_494 dout0_495 dout0_496 dout0_497 dout0_498
+ dout0_499 dout0_500 dout0_501 dout0_502 dout0_503 dout0_504 dout0_505
+ dout0_506 dout0_507 dout0_508 dout0_509 dout0_510 dout0_511 rbl_bl_0_0
+ din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9
+ din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17
+ din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25
+ din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 din0_32 din0_33
+ din0_34 din0_35 din0_36 din0_37 din0_38 din0_39 din0_40 din0_41
+ din0_42 din0_43 din0_44 din0_45 din0_46 din0_47 din0_48 din0_49
+ din0_50 din0_51 din0_52 din0_53 din0_54 din0_55 din0_56 din0_57
+ din0_58 din0_59 din0_60 din0_61 din0_62 din0_63 din0_64 din0_65
+ din0_66 din0_67 din0_68 din0_69 din0_70 din0_71 din0_72 din0_73
+ din0_74 din0_75 din0_76 din0_77 din0_78 din0_79 din0_80 din0_81
+ din0_82 din0_83 din0_84 din0_85 din0_86 din0_87 din0_88 din0_89
+ din0_90 din0_91 din0_92 din0_93 din0_94 din0_95 din0_96 din0_97
+ din0_98 din0_99 din0_100 din0_101 din0_102 din0_103 din0_104 din0_105
+ din0_106 din0_107 din0_108 din0_109 din0_110 din0_111 din0_112
+ din0_113 din0_114 din0_115 din0_116 din0_117 din0_118 din0_119
+ din0_120 din0_121 din0_122 din0_123 din0_124 din0_125 din0_126
+ din0_127 din0_128 din0_129 din0_130 din0_131 din0_132 din0_133
+ din0_134 din0_135 din0_136 din0_137 din0_138 din0_139 din0_140
+ din0_141 din0_142 din0_143 din0_144 din0_145 din0_146 din0_147
+ din0_148 din0_149 din0_150 din0_151 din0_152 din0_153 din0_154
+ din0_155 din0_156 din0_157 din0_158 din0_159 din0_160 din0_161
+ din0_162 din0_163 din0_164 din0_165 din0_166 din0_167 din0_168
+ din0_169 din0_170 din0_171 din0_172 din0_173 din0_174 din0_175
+ din0_176 din0_177 din0_178 din0_179 din0_180 din0_181 din0_182
+ din0_183 din0_184 din0_185 din0_186 din0_187 din0_188 din0_189
+ din0_190 din0_191 din0_192 din0_193 din0_194 din0_195 din0_196
+ din0_197 din0_198 din0_199 din0_200 din0_201 din0_202 din0_203
+ din0_204 din0_205 din0_206 din0_207 din0_208 din0_209 din0_210
+ din0_211 din0_212 din0_213 din0_214 din0_215 din0_216 din0_217
+ din0_218 din0_219 din0_220 din0_221 din0_222 din0_223 din0_224
+ din0_225 din0_226 din0_227 din0_228 din0_229 din0_230 din0_231
+ din0_232 din0_233 din0_234 din0_235 din0_236 din0_237 din0_238
+ din0_239 din0_240 din0_241 din0_242 din0_243 din0_244 din0_245
+ din0_246 din0_247 din0_248 din0_249 din0_250 din0_251 din0_252
+ din0_253 din0_254 din0_255 din0_256 din0_257 din0_258 din0_259
+ din0_260 din0_261 din0_262 din0_263 din0_264 din0_265 din0_266
+ din0_267 din0_268 din0_269 din0_270 din0_271 din0_272 din0_273
+ din0_274 din0_275 din0_276 din0_277 din0_278 din0_279 din0_280
+ din0_281 din0_282 din0_283 din0_284 din0_285 din0_286 din0_287
+ din0_288 din0_289 din0_290 din0_291 din0_292 din0_293 din0_294
+ din0_295 din0_296 din0_297 din0_298 din0_299 din0_300 din0_301
+ din0_302 din0_303 din0_304 din0_305 din0_306 din0_307 din0_308
+ din0_309 din0_310 din0_311 din0_312 din0_313 din0_314 din0_315
+ din0_316 din0_317 din0_318 din0_319 din0_320 din0_321 din0_322
+ din0_323 din0_324 din0_325 din0_326 din0_327 din0_328 din0_329
+ din0_330 din0_331 din0_332 din0_333 din0_334 din0_335 din0_336
+ din0_337 din0_338 din0_339 din0_340 din0_341 din0_342 din0_343
+ din0_344 din0_345 din0_346 din0_347 din0_348 din0_349 din0_350
+ din0_351 din0_352 din0_353 din0_354 din0_355 din0_356 din0_357
+ din0_358 din0_359 din0_360 din0_361 din0_362 din0_363 din0_364
+ din0_365 din0_366 din0_367 din0_368 din0_369 din0_370 din0_371
+ din0_372 din0_373 din0_374 din0_375 din0_376 din0_377 din0_378
+ din0_379 din0_380 din0_381 din0_382 din0_383 din0_384 din0_385
+ din0_386 din0_387 din0_388 din0_389 din0_390 din0_391 din0_392
+ din0_393 din0_394 din0_395 din0_396 din0_397 din0_398 din0_399
+ din0_400 din0_401 din0_402 din0_403 din0_404 din0_405 din0_406
+ din0_407 din0_408 din0_409 din0_410 din0_411 din0_412 din0_413
+ din0_414 din0_415 din0_416 din0_417 din0_418 din0_419 din0_420
+ din0_421 din0_422 din0_423 din0_424 din0_425 din0_426 din0_427
+ din0_428 din0_429 din0_430 din0_431 din0_432 din0_433 din0_434
+ din0_435 din0_436 din0_437 din0_438 din0_439 din0_440 din0_441
+ din0_442 din0_443 din0_444 din0_445 din0_446 din0_447 din0_448
+ din0_449 din0_450 din0_451 din0_452 din0_453 din0_454 din0_455
+ din0_456 din0_457 din0_458 din0_459 din0_460 din0_461 din0_462
+ din0_463 din0_464 din0_465 din0_466 din0_467 din0_468 din0_469
+ din0_470 din0_471 din0_472 din0_473 din0_474 din0_475 din0_476
+ din0_477 din0_478 din0_479 din0_480 din0_481 din0_482 din0_483
+ din0_484 din0_485 din0_486 din0_487 din0_488 din0_489 din0_490
+ din0_491 din0_492 din0_493 din0_494 din0_495 din0_496 din0_497
+ din0_498 din0_499 din0_500 din0_501 din0_502 din0_503 din0_504
+ din0_505 din0_506 din0_507 din0_508 din0_509 din0_510 din0_511 addr0_0
+ addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 s_en0 p_en_bar0 w_en0 wl_en0
+ vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: dout0_32 
* OUTPUT: dout0_33 
* OUTPUT: dout0_34 
* OUTPUT: dout0_35 
* OUTPUT: dout0_36 
* OUTPUT: dout0_37 
* OUTPUT: dout0_38 
* OUTPUT: dout0_39 
* OUTPUT: dout0_40 
* OUTPUT: dout0_41 
* OUTPUT: dout0_42 
* OUTPUT: dout0_43 
* OUTPUT: dout0_44 
* OUTPUT: dout0_45 
* OUTPUT: dout0_46 
* OUTPUT: dout0_47 
* OUTPUT: dout0_48 
* OUTPUT: dout0_49 
* OUTPUT: dout0_50 
* OUTPUT: dout0_51 
* OUTPUT: dout0_52 
* OUTPUT: dout0_53 
* OUTPUT: dout0_54 
* OUTPUT: dout0_55 
* OUTPUT: dout0_56 
* OUTPUT: dout0_57 
* OUTPUT: dout0_58 
* OUTPUT: dout0_59 
* OUTPUT: dout0_60 
* OUTPUT: dout0_61 
* OUTPUT: dout0_62 
* OUTPUT: dout0_63 
* OUTPUT: dout0_64 
* OUTPUT: dout0_65 
* OUTPUT: dout0_66 
* OUTPUT: dout0_67 
* OUTPUT: dout0_68 
* OUTPUT: dout0_69 
* OUTPUT: dout0_70 
* OUTPUT: dout0_71 
* OUTPUT: dout0_72 
* OUTPUT: dout0_73 
* OUTPUT: dout0_74 
* OUTPUT: dout0_75 
* OUTPUT: dout0_76 
* OUTPUT: dout0_77 
* OUTPUT: dout0_78 
* OUTPUT: dout0_79 
* OUTPUT: dout0_80 
* OUTPUT: dout0_81 
* OUTPUT: dout0_82 
* OUTPUT: dout0_83 
* OUTPUT: dout0_84 
* OUTPUT: dout0_85 
* OUTPUT: dout0_86 
* OUTPUT: dout0_87 
* OUTPUT: dout0_88 
* OUTPUT: dout0_89 
* OUTPUT: dout0_90 
* OUTPUT: dout0_91 
* OUTPUT: dout0_92 
* OUTPUT: dout0_93 
* OUTPUT: dout0_94 
* OUTPUT: dout0_95 
* OUTPUT: dout0_96 
* OUTPUT: dout0_97 
* OUTPUT: dout0_98 
* OUTPUT: dout0_99 
* OUTPUT: dout0_100 
* OUTPUT: dout0_101 
* OUTPUT: dout0_102 
* OUTPUT: dout0_103 
* OUTPUT: dout0_104 
* OUTPUT: dout0_105 
* OUTPUT: dout0_106 
* OUTPUT: dout0_107 
* OUTPUT: dout0_108 
* OUTPUT: dout0_109 
* OUTPUT: dout0_110 
* OUTPUT: dout0_111 
* OUTPUT: dout0_112 
* OUTPUT: dout0_113 
* OUTPUT: dout0_114 
* OUTPUT: dout0_115 
* OUTPUT: dout0_116 
* OUTPUT: dout0_117 
* OUTPUT: dout0_118 
* OUTPUT: dout0_119 
* OUTPUT: dout0_120 
* OUTPUT: dout0_121 
* OUTPUT: dout0_122 
* OUTPUT: dout0_123 
* OUTPUT: dout0_124 
* OUTPUT: dout0_125 
* OUTPUT: dout0_126 
* OUTPUT: dout0_127 
* OUTPUT: dout0_128 
* OUTPUT: dout0_129 
* OUTPUT: dout0_130 
* OUTPUT: dout0_131 
* OUTPUT: dout0_132 
* OUTPUT: dout0_133 
* OUTPUT: dout0_134 
* OUTPUT: dout0_135 
* OUTPUT: dout0_136 
* OUTPUT: dout0_137 
* OUTPUT: dout0_138 
* OUTPUT: dout0_139 
* OUTPUT: dout0_140 
* OUTPUT: dout0_141 
* OUTPUT: dout0_142 
* OUTPUT: dout0_143 
* OUTPUT: dout0_144 
* OUTPUT: dout0_145 
* OUTPUT: dout0_146 
* OUTPUT: dout0_147 
* OUTPUT: dout0_148 
* OUTPUT: dout0_149 
* OUTPUT: dout0_150 
* OUTPUT: dout0_151 
* OUTPUT: dout0_152 
* OUTPUT: dout0_153 
* OUTPUT: dout0_154 
* OUTPUT: dout0_155 
* OUTPUT: dout0_156 
* OUTPUT: dout0_157 
* OUTPUT: dout0_158 
* OUTPUT: dout0_159 
* OUTPUT: dout0_160 
* OUTPUT: dout0_161 
* OUTPUT: dout0_162 
* OUTPUT: dout0_163 
* OUTPUT: dout0_164 
* OUTPUT: dout0_165 
* OUTPUT: dout0_166 
* OUTPUT: dout0_167 
* OUTPUT: dout0_168 
* OUTPUT: dout0_169 
* OUTPUT: dout0_170 
* OUTPUT: dout0_171 
* OUTPUT: dout0_172 
* OUTPUT: dout0_173 
* OUTPUT: dout0_174 
* OUTPUT: dout0_175 
* OUTPUT: dout0_176 
* OUTPUT: dout0_177 
* OUTPUT: dout0_178 
* OUTPUT: dout0_179 
* OUTPUT: dout0_180 
* OUTPUT: dout0_181 
* OUTPUT: dout0_182 
* OUTPUT: dout0_183 
* OUTPUT: dout0_184 
* OUTPUT: dout0_185 
* OUTPUT: dout0_186 
* OUTPUT: dout0_187 
* OUTPUT: dout0_188 
* OUTPUT: dout0_189 
* OUTPUT: dout0_190 
* OUTPUT: dout0_191 
* OUTPUT: dout0_192 
* OUTPUT: dout0_193 
* OUTPUT: dout0_194 
* OUTPUT: dout0_195 
* OUTPUT: dout0_196 
* OUTPUT: dout0_197 
* OUTPUT: dout0_198 
* OUTPUT: dout0_199 
* OUTPUT: dout0_200 
* OUTPUT: dout0_201 
* OUTPUT: dout0_202 
* OUTPUT: dout0_203 
* OUTPUT: dout0_204 
* OUTPUT: dout0_205 
* OUTPUT: dout0_206 
* OUTPUT: dout0_207 
* OUTPUT: dout0_208 
* OUTPUT: dout0_209 
* OUTPUT: dout0_210 
* OUTPUT: dout0_211 
* OUTPUT: dout0_212 
* OUTPUT: dout0_213 
* OUTPUT: dout0_214 
* OUTPUT: dout0_215 
* OUTPUT: dout0_216 
* OUTPUT: dout0_217 
* OUTPUT: dout0_218 
* OUTPUT: dout0_219 
* OUTPUT: dout0_220 
* OUTPUT: dout0_221 
* OUTPUT: dout0_222 
* OUTPUT: dout0_223 
* OUTPUT: dout0_224 
* OUTPUT: dout0_225 
* OUTPUT: dout0_226 
* OUTPUT: dout0_227 
* OUTPUT: dout0_228 
* OUTPUT: dout0_229 
* OUTPUT: dout0_230 
* OUTPUT: dout0_231 
* OUTPUT: dout0_232 
* OUTPUT: dout0_233 
* OUTPUT: dout0_234 
* OUTPUT: dout0_235 
* OUTPUT: dout0_236 
* OUTPUT: dout0_237 
* OUTPUT: dout0_238 
* OUTPUT: dout0_239 
* OUTPUT: dout0_240 
* OUTPUT: dout0_241 
* OUTPUT: dout0_242 
* OUTPUT: dout0_243 
* OUTPUT: dout0_244 
* OUTPUT: dout0_245 
* OUTPUT: dout0_246 
* OUTPUT: dout0_247 
* OUTPUT: dout0_248 
* OUTPUT: dout0_249 
* OUTPUT: dout0_250 
* OUTPUT: dout0_251 
* OUTPUT: dout0_252 
* OUTPUT: dout0_253 
* OUTPUT: dout0_254 
* OUTPUT: dout0_255 
* OUTPUT: dout0_256 
* OUTPUT: dout0_257 
* OUTPUT: dout0_258 
* OUTPUT: dout0_259 
* OUTPUT: dout0_260 
* OUTPUT: dout0_261 
* OUTPUT: dout0_262 
* OUTPUT: dout0_263 
* OUTPUT: dout0_264 
* OUTPUT: dout0_265 
* OUTPUT: dout0_266 
* OUTPUT: dout0_267 
* OUTPUT: dout0_268 
* OUTPUT: dout0_269 
* OUTPUT: dout0_270 
* OUTPUT: dout0_271 
* OUTPUT: dout0_272 
* OUTPUT: dout0_273 
* OUTPUT: dout0_274 
* OUTPUT: dout0_275 
* OUTPUT: dout0_276 
* OUTPUT: dout0_277 
* OUTPUT: dout0_278 
* OUTPUT: dout0_279 
* OUTPUT: dout0_280 
* OUTPUT: dout0_281 
* OUTPUT: dout0_282 
* OUTPUT: dout0_283 
* OUTPUT: dout0_284 
* OUTPUT: dout0_285 
* OUTPUT: dout0_286 
* OUTPUT: dout0_287 
* OUTPUT: dout0_288 
* OUTPUT: dout0_289 
* OUTPUT: dout0_290 
* OUTPUT: dout0_291 
* OUTPUT: dout0_292 
* OUTPUT: dout0_293 
* OUTPUT: dout0_294 
* OUTPUT: dout0_295 
* OUTPUT: dout0_296 
* OUTPUT: dout0_297 
* OUTPUT: dout0_298 
* OUTPUT: dout0_299 
* OUTPUT: dout0_300 
* OUTPUT: dout0_301 
* OUTPUT: dout0_302 
* OUTPUT: dout0_303 
* OUTPUT: dout0_304 
* OUTPUT: dout0_305 
* OUTPUT: dout0_306 
* OUTPUT: dout0_307 
* OUTPUT: dout0_308 
* OUTPUT: dout0_309 
* OUTPUT: dout0_310 
* OUTPUT: dout0_311 
* OUTPUT: dout0_312 
* OUTPUT: dout0_313 
* OUTPUT: dout0_314 
* OUTPUT: dout0_315 
* OUTPUT: dout0_316 
* OUTPUT: dout0_317 
* OUTPUT: dout0_318 
* OUTPUT: dout0_319 
* OUTPUT: dout0_320 
* OUTPUT: dout0_321 
* OUTPUT: dout0_322 
* OUTPUT: dout0_323 
* OUTPUT: dout0_324 
* OUTPUT: dout0_325 
* OUTPUT: dout0_326 
* OUTPUT: dout0_327 
* OUTPUT: dout0_328 
* OUTPUT: dout0_329 
* OUTPUT: dout0_330 
* OUTPUT: dout0_331 
* OUTPUT: dout0_332 
* OUTPUT: dout0_333 
* OUTPUT: dout0_334 
* OUTPUT: dout0_335 
* OUTPUT: dout0_336 
* OUTPUT: dout0_337 
* OUTPUT: dout0_338 
* OUTPUT: dout0_339 
* OUTPUT: dout0_340 
* OUTPUT: dout0_341 
* OUTPUT: dout0_342 
* OUTPUT: dout0_343 
* OUTPUT: dout0_344 
* OUTPUT: dout0_345 
* OUTPUT: dout0_346 
* OUTPUT: dout0_347 
* OUTPUT: dout0_348 
* OUTPUT: dout0_349 
* OUTPUT: dout0_350 
* OUTPUT: dout0_351 
* OUTPUT: dout0_352 
* OUTPUT: dout0_353 
* OUTPUT: dout0_354 
* OUTPUT: dout0_355 
* OUTPUT: dout0_356 
* OUTPUT: dout0_357 
* OUTPUT: dout0_358 
* OUTPUT: dout0_359 
* OUTPUT: dout0_360 
* OUTPUT: dout0_361 
* OUTPUT: dout0_362 
* OUTPUT: dout0_363 
* OUTPUT: dout0_364 
* OUTPUT: dout0_365 
* OUTPUT: dout0_366 
* OUTPUT: dout0_367 
* OUTPUT: dout0_368 
* OUTPUT: dout0_369 
* OUTPUT: dout0_370 
* OUTPUT: dout0_371 
* OUTPUT: dout0_372 
* OUTPUT: dout0_373 
* OUTPUT: dout0_374 
* OUTPUT: dout0_375 
* OUTPUT: dout0_376 
* OUTPUT: dout0_377 
* OUTPUT: dout0_378 
* OUTPUT: dout0_379 
* OUTPUT: dout0_380 
* OUTPUT: dout0_381 
* OUTPUT: dout0_382 
* OUTPUT: dout0_383 
* OUTPUT: dout0_384 
* OUTPUT: dout0_385 
* OUTPUT: dout0_386 
* OUTPUT: dout0_387 
* OUTPUT: dout0_388 
* OUTPUT: dout0_389 
* OUTPUT: dout0_390 
* OUTPUT: dout0_391 
* OUTPUT: dout0_392 
* OUTPUT: dout0_393 
* OUTPUT: dout0_394 
* OUTPUT: dout0_395 
* OUTPUT: dout0_396 
* OUTPUT: dout0_397 
* OUTPUT: dout0_398 
* OUTPUT: dout0_399 
* OUTPUT: dout0_400 
* OUTPUT: dout0_401 
* OUTPUT: dout0_402 
* OUTPUT: dout0_403 
* OUTPUT: dout0_404 
* OUTPUT: dout0_405 
* OUTPUT: dout0_406 
* OUTPUT: dout0_407 
* OUTPUT: dout0_408 
* OUTPUT: dout0_409 
* OUTPUT: dout0_410 
* OUTPUT: dout0_411 
* OUTPUT: dout0_412 
* OUTPUT: dout0_413 
* OUTPUT: dout0_414 
* OUTPUT: dout0_415 
* OUTPUT: dout0_416 
* OUTPUT: dout0_417 
* OUTPUT: dout0_418 
* OUTPUT: dout0_419 
* OUTPUT: dout0_420 
* OUTPUT: dout0_421 
* OUTPUT: dout0_422 
* OUTPUT: dout0_423 
* OUTPUT: dout0_424 
* OUTPUT: dout0_425 
* OUTPUT: dout0_426 
* OUTPUT: dout0_427 
* OUTPUT: dout0_428 
* OUTPUT: dout0_429 
* OUTPUT: dout0_430 
* OUTPUT: dout0_431 
* OUTPUT: dout0_432 
* OUTPUT: dout0_433 
* OUTPUT: dout0_434 
* OUTPUT: dout0_435 
* OUTPUT: dout0_436 
* OUTPUT: dout0_437 
* OUTPUT: dout0_438 
* OUTPUT: dout0_439 
* OUTPUT: dout0_440 
* OUTPUT: dout0_441 
* OUTPUT: dout0_442 
* OUTPUT: dout0_443 
* OUTPUT: dout0_444 
* OUTPUT: dout0_445 
* OUTPUT: dout0_446 
* OUTPUT: dout0_447 
* OUTPUT: dout0_448 
* OUTPUT: dout0_449 
* OUTPUT: dout0_450 
* OUTPUT: dout0_451 
* OUTPUT: dout0_452 
* OUTPUT: dout0_453 
* OUTPUT: dout0_454 
* OUTPUT: dout0_455 
* OUTPUT: dout0_456 
* OUTPUT: dout0_457 
* OUTPUT: dout0_458 
* OUTPUT: dout0_459 
* OUTPUT: dout0_460 
* OUTPUT: dout0_461 
* OUTPUT: dout0_462 
* OUTPUT: dout0_463 
* OUTPUT: dout0_464 
* OUTPUT: dout0_465 
* OUTPUT: dout0_466 
* OUTPUT: dout0_467 
* OUTPUT: dout0_468 
* OUTPUT: dout0_469 
* OUTPUT: dout0_470 
* OUTPUT: dout0_471 
* OUTPUT: dout0_472 
* OUTPUT: dout0_473 
* OUTPUT: dout0_474 
* OUTPUT: dout0_475 
* OUTPUT: dout0_476 
* OUTPUT: dout0_477 
* OUTPUT: dout0_478 
* OUTPUT: dout0_479 
* OUTPUT: dout0_480 
* OUTPUT: dout0_481 
* OUTPUT: dout0_482 
* OUTPUT: dout0_483 
* OUTPUT: dout0_484 
* OUTPUT: dout0_485 
* OUTPUT: dout0_486 
* OUTPUT: dout0_487 
* OUTPUT: dout0_488 
* OUTPUT: dout0_489 
* OUTPUT: dout0_490 
* OUTPUT: dout0_491 
* OUTPUT: dout0_492 
* OUTPUT: dout0_493 
* OUTPUT: dout0_494 
* OUTPUT: dout0_495 
* OUTPUT: dout0_496 
* OUTPUT: dout0_497 
* OUTPUT: dout0_498 
* OUTPUT: dout0_499 
* OUTPUT: dout0_500 
* OUTPUT: dout0_501 
* OUTPUT: dout0_502 
* OUTPUT: dout0_503 
* OUTPUT: dout0_504 
* OUTPUT: dout0_505 
* OUTPUT: dout0_506 
* OUTPUT: dout0_507 
* OUTPUT: dout0_508 
* OUTPUT: dout0_509 
* OUTPUT: dout0_510 
* OUTPUT: dout0_511 
* OUTPUT: rbl_bl_0_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : din0_32 
* INPUT : din0_33 
* INPUT : din0_34 
* INPUT : din0_35 
* INPUT : din0_36 
* INPUT : din0_37 
* INPUT : din0_38 
* INPUT : din0_39 
* INPUT : din0_40 
* INPUT : din0_41 
* INPUT : din0_42 
* INPUT : din0_43 
* INPUT : din0_44 
* INPUT : din0_45 
* INPUT : din0_46 
* INPUT : din0_47 
* INPUT : din0_48 
* INPUT : din0_49 
* INPUT : din0_50 
* INPUT : din0_51 
* INPUT : din0_52 
* INPUT : din0_53 
* INPUT : din0_54 
* INPUT : din0_55 
* INPUT : din0_56 
* INPUT : din0_57 
* INPUT : din0_58 
* INPUT : din0_59 
* INPUT : din0_60 
* INPUT : din0_61 
* INPUT : din0_62 
* INPUT : din0_63 
* INPUT : din0_64 
* INPUT : din0_65 
* INPUT : din0_66 
* INPUT : din0_67 
* INPUT : din0_68 
* INPUT : din0_69 
* INPUT : din0_70 
* INPUT : din0_71 
* INPUT : din0_72 
* INPUT : din0_73 
* INPUT : din0_74 
* INPUT : din0_75 
* INPUT : din0_76 
* INPUT : din0_77 
* INPUT : din0_78 
* INPUT : din0_79 
* INPUT : din0_80 
* INPUT : din0_81 
* INPUT : din0_82 
* INPUT : din0_83 
* INPUT : din0_84 
* INPUT : din0_85 
* INPUT : din0_86 
* INPUT : din0_87 
* INPUT : din0_88 
* INPUT : din0_89 
* INPUT : din0_90 
* INPUT : din0_91 
* INPUT : din0_92 
* INPUT : din0_93 
* INPUT : din0_94 
* INPUT : din0_95 
* INPUT : din0_96 
* INPUT : din0_97 
* INPUT : din0_98 
* INPUT : din0_99 
* INPUT : din0_100 
* INPUT : din0_101 
* INPUT : din0_102 
* INPUT : din0_103 
* INPUT : din0_104 
* INPUT : din0_105 
* INPUT : din0_106 
* INPUT : din0_107 
* INPUT : din0_108 
* INPUT : din0_109 
* INPUT : din0_110 
* INPUT : din0_111 
* INPUT : din0_112 
* INPUT : din0_113 
* INPUT : din0_114 
* INPUT : din0_115 
* INPUT : din0_116 
* INPUT : din0_117 
* INPUT : din0_118 
* INPUT : din0_119 
* INPUT : din0_120 
* INPUT : din0_121 
* INPUT : din0_122 
* INPUT : din0_123 
* INPUT : din0_124 
* INPUT : din0_125 
* INPUT : din0_126 
* INPUT : din0_127 
* INPUT : din0_128 
* INPUT : din0_129 
* INPUT : din0_130 
* INPUT : din0_131 
* INPUT : din0_132 
* INPUT : din0_133 
* INPUT : din0_134 
* INPUT : din0_135 
* INPUT : din0_136 
* INPUT : din0_137 
* INPUT : din0_138 
* INPUT : din0_139 
* INPUT : din0_140 
* INPUT : din0_141 
* INPUT : din0_142 
* INPUT : din0_143 
* INPUT : din0_144 
* INPUT : din0_145 
* INPUT : din0_146 
* INPUT : din0_147 
* INPUT : din0_148 
* INPUT : din0_149 
* INPUT : din0_150 
* INPUT : din0_151 
* INPUT : din0_152 
* INPUT : din0_153 
* INPUT : din0_154 
* INPUT : din0_155 
* INPUT : din0_156 
* INPUT : din0_157 
* INPUT : din0_158 
* INPUT : din0_159 
* INPUT : din0_160 
* INPUT : din0_161 
* INPUT : din0_162 
* INPUT : din0_163 
* INPUT : din0_164 
* INPUT : din0_165 
* INPUT : din0_166 
* INPUT : din0_167 
* INPUT : din0_168 
* INPUT : din0_169 
* INPUT : din0_170 
* INPUT : din0_171 
* INPUT : din0_172 
* INPUT : din0_173 
* INPUT : din0_174 
* INPUT : din0_175 
* INPUT : din0_176 
* INPUT : din0_177 
* INPUT : din0_178 
* INPUT : din0_179 
* INPUT : din0_180 
* INPUT : din0_181 
* INPUT : din0_182 
* INPUT : din0_183 
* INPUT : din0_184 
* INPUT : din0_185 
* INPUT : din0_186 
* INPUT : din0_187 
* INPUT : din0_188 
* INPUT : din0_189 
* INPUT : din0_190 
* INPUT : din0_191 
* INPUT : din0_192 
* INPUT : din0_193 
* INPUT : din0_194 
* INPUT : din0_195 
* INPUT : din0_196 
* INPUT : din0_197 
* INPUT : din0_198 
* INPUT : din0_199 
* INPUT : din0_200 
* INPUT : din0_201 
* INPUT : din0_202 
* INPUT : din0_203 
* INPUT : din0_204 
* INPUT : din0_205 
* INPUT : din0_206 
* INPUT : din0_207 
* INPUT : din0_208 
* INPUT : din0_209 
* INPUT : din0_210 
* INPUT : din0_211 
* INPUT : din0_212 
* INPUT : din0_213 
* INPUT : din0_214 
* INPUT : din0_215 
* INPUT : din0_216 
* INPUT : din0_217 
* INPUT : din0_218 
* INPUT : din0_219 
* INPUT : din0_220 
* INPUT : din0_221 
* INPUT : din0_222 
* INPUT : din0_223 
* INPUT : din0_224 
* INPUT : din0_225 
* INPUT : din0_226 
* INPUT : din0_227 
* INPUT : din0_228 
* INPUT : din0_229 
* INPUT : din0_230 
* INPUT : din0_231 
* INPUT : din0_232 
* INPUT : din0_233 
* INPUT : din0_234 
* INPUT : din0_235 
* INPUT : din0_236 
* INPUT : din0_237 
* INPUT : din0_238 
* INPUT : din0_239 
* INPUT : din0_240 
* INPUT : din0_241 
* INPUT : din0_242 
* INPUT : din0_243 
* INPUT : din0_244 
* INPUT : din0_245 
* INPUT : din0_246 
* INPUT : din0_247 
* INPUT : din0_248 
* INPUT : din0_249 
* INPUT : din0_250 
* INPUT : din0_251 
* INPUT : din0_252 
* INPUT : din0_253 
* INPUT : din0_254 
* INPUT : din0_255 
* INPUT : din0_256 
* INPUT : din0_257 
* INPUT : din0_258 
* INPUT : din0_259 
* INPUT : din0_260 
* INPUT : din0_261 
* INPUT : din0_262 
* INPUT : din0_263 
* INPUT : din0_264 
* INPUT : din0_265 
* INPUT : din0_266 
* INPUT : din0_267 
* INPUT : din0_268 
* INPUT : din0_269 
* INPUT : din0_270 
* INPUT : din0_271 
* INPUT : din0_272 
* INPUT : din0_273 
* INPUT : din0_274 
* INPUT : din0_275 
* INPUT : din0_276 
* INPUT : din0_277 
* INPUT : din0_278 
* INPUT : din0_279 
* INPUT : din0_280 
* INPUT : din0_281 
* INPUT : din0_282 
* INPUT : din0_283 
* INPUT : din0_284 
* INPUT : din0_285 
* INPUT : din0_286 
* INPUT : din0_287 
* INPUT : din0_288 
* INPUT : din0_289 
* INPUT : din0_290 
* INPUT : din0_291 
* INPUT : din0_292 
* INPUT : din0_293 
* INPUT : din0_294 
* INPUT : din0_295 
* INPUT : din0_296 
* INPUT : din0_297 
* INPUT : din0_298 
* INPUT : din0_299 
* INPUT : din0_300 
* INPUT : din0_301 
* INPUT : din0_302 
* INPUT : din0_303 
* INPUT : din0_304 
* INPUT : din0_305 
* INPUT : din0_306 
* INPUT : din0_307 
* INPUT : din0_308 
* INPUT : din0_309 
* INPUT : din0_310 
* INPUT : din0_311 
* INPUT : din0_312 
* INPUT : din0_313 
* INPUT : din0_314 
* INPUT : din0_315 
* INPUT : din0_316 
* INPUT : din0_317 
* INPUT : din0_318 
* INPUT : din0_319 
* INPUT : din0_320 
* INPUT : din0_321 
* INPUT : din0_322 
* INPUT : din0_323 
* INPUT : din0_324 
* INPUT : din0_325 
* INPUT : din0_326 
* INPUT : din0_327 
* INPUT : din0_328 
* INPUT : din0_329 
* INPUT : din0_330 
* INPUT : din0_331 
* INPUT : din0_332 
* INPUT : din0_333 
* INPUT : din0_334 
* INPUT : din0_335 
* INPUT : din0_336 
* INPUT : din0_337 
* INPUT : din0_338 
* INPUT : din0_339 
* INPUT : din0_340 
* INPUT : din0_341 
* INPUT : din0_342 
* INPUT : din0_343 
* INPUT : din0_344 
* INPUT : din0_345 
* INPUT : din0_346 
* INPUT : din0_347 
* INPUT : din0_348 
* INPUT : din0_349 
* INPUT : din0_350 
* INPUT : din0_351 
* INPUT : din0_352 
* INPUT : din0_353 
* INPUT : din0_354 
* INPUT : din0_355 
* INPUT : din0_356 
* INPUT : din0_357 
* INPUT : din0_358 
* INPUT : din0_359 
* INPUT : din0_360 
* INPUT : din0_361 
* INPUT : din0_362 
* INPUT : din0_363 
* INPUT : din0_364 
* INPUT : din0_365 
* INPUT : din0_366 
* INPUT : din0_367 
* INPUT : din0_368 
* INPUT : din0_369 
* INPUT : din0_370 
* INPUT : din0_371 
* INPUT : din0_372 
* INPUT : din0_373 
* INPUT : din0_374 
* INPUT : din0_375 
* INPUT : din0_376 
* INPUT : din0_377 
* INPUT : din0_378 
* INPUT : din0_379 
* INPUT : din0_380 
* INPUT : din0_381 
* INPUT : din0_382 
* INPUT : din0_383 
* INPUT : din0_384 
* INPUT : din0_385 
* INPUT : din0_386 
* INPUT : din0_387 
* INPUT : din0_388 
* INPUT : din0_389 
* INPUT : din0_390 
* INPUT : din0_391 
* INPUT : din0_392 
* INPUT : din0_393 
* INPUT : din0_394 
* INPUT : din0_395 
* INPUT : din0_396 
* INPUT : din0_397 
* INPUT : din0_398 
* INPUT : din0_399 
* INPUT : din0_400 
* INPUT : din0_401 
* INPUT : din0_402 
* INPUT : din0_403 
* INPUT : din0_404 
* INPUT : din0_405 
* INPUT : din0_406 
* INPUT : din0_407 
* INPUT : din0_408 
* INPUT : din0_409 
* INPUT : din0_410 
* INPUT : din0_411 
* INPUT : din0_412 
* INPUT : din0_413 
* INPUT : din0_414 
* INPUT : din0_415 
* INPUT : din0_416 
* INPUT : din0_417 
* INPUT : din0_418 
* INPUT : din0_419 
* INPUT : din0_420 
* INPUT : din0_421 
* INPUT : din0_422 
* INPUT : din0_423 
* INPUT : din0_424 
* INPUT : din0_425 
* INPUT : din0_426 
* INPUT : din0_427 
* INPUT : din0_428 
* INPUT : din0_429 
* INPUT : din0_430 
* INPUT : din0_431 
* INPUT : din0_432 
* INPUT : din0_433 
* INPUT : din0_434 
* INPUT : din0_435 
* INPUT : din0_436 
* INPUT : din0_437 
* INPUT : din0_438 
* INPUT : din0_439 
* INPUT : din0_440 
* INPUT : din0_441 
* INPUT : din0_442 
* INPUT : din0_443 
* INPUT : din0_444 
* INPUT : din0_445 
* INPUT : din0_446 
* INPUT : din0_447 
* INPUT : din0_448 
* INPUT : din0_449 
* INPUT : din0_450 
* INPUT : din0_451 
* INPUT : din0_452 
* INPUT : din0_453 
* INPUT : din0_454 
* INPUT : din0_455 
* INPUT : din0_456 
* INPUT : din0_457 
* INPUT : din0_458 
* INPUT : din0_459 
* INPUT : din0_460 
* INPUT : din0_461 
* INPUT : din0_462 
* INPUT : din0_463 
* INPUT : din0_464 
* INPUT : din0_465 
* INPUT : din0_466 
* INPUT : din0_467 
* INPUT : din0_468 
* INPUT : din0_469 
* INPUT : din0_470 
* INPUT : din0_471 
* INPUT : din0_472 
* INPUT : din0_473 
* INPUT : din0_474 
* INPUT : din0_475 
* INPUT : din0_476 
* INPUT : din0_477 
* INPUT : din0_478 
* INPUT : din0_479 
* INPUT : din0_480 
* INPUT : din0_481 
* INPUT : din0_482 
* INPUT : din0_483 
* INPUT : din0_484 
* INPUT : din0_485 
* INPUT : din0_486 
* INPUT : din0_487 
* INPUT : din0_488 
* INPUT : din0_489 
* INPUT : din0_490 
* INPUT : din0_491 
* INPUT : din0_492 
* INPUT : din0_493 
* INPUT : din0_494 
* INPUT : din0_495 
* INPUT : din0_496 
* INPUT : din0_497 
* INPUT : din0_498 
* INPUT : din0_499 
* INPUT : din0_500 
* INPUT : din0_501 
* INPUT : din0_502 
* INPUT : din0_503 
* INPUT : din0_504 
* INPUT : din0_505 
* INPUT : din0_506 
* INPUT : din0_507 
* INPUT : din0_508 
* INPUT : din0_509 
* INPUT : din0_510 
* INPUT : din0_511 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xbitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258
+ br_0_258 bl_0_259 br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261
+ bl_0_262 br_0_262 bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265
+ br_0_265 bl_0_266 br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268
+ bl_0_269 br_0_269 bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272
+ br_0_272 bl_0_273 br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275
+ bl_0_276 br_0_276 bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279
+ br_0_279 bl_0_280 br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282
+ bl_0_283 br_0_283 bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286
+ br_0_286 bl_0_287 br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289
+ bl_0_290 br_0_290 bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293
+ br_0_293 bl_0_294 br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296
+ bl_0_297 br_0_297 bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300
+ br_0_300 bl_0_301 br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303
+ bl_0_304 br_0_304 bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307
+ br_0_307 bl_0_308 br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310
+ bl_0_311 br_0_311 bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314
+ br_0_314 bl_0_315 br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317
+ bl_0_318 br_0_318 bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321
+ br_0_321 bl_0_322 br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324
+ bl_0_325 br_0_325 bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328
+ br_0_328 bl_0_329 br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331
+ bl_0_332 br_0_332 bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335
+ br_0_335 bl_0_336 br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338
+ bl_0_339 br_0_339 bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342
+ br_0_342 bl_0_343 br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345
+ bl_0_346 br_0_346 bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349
+ br_0_349 bl_0_350 br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352
+ bl_0_353 br_0_353 bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356
+ br_0_356 bl_0_357 br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359
+ bl_0_360 br_0_360 bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363
+ br_0_363 bl_0_364 br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366
+ bl_0_367 br_0_367 bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370
+ br_0_370 bl_0_371 br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373
+ bl_0_374 br_0_374 bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377
+ br_0_377 bl_0_378 br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380
+ bl_0_381 br_0_381 bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384
+ br_0_384 bl_0_385 br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387
+ bl_0_388 br_0_388 bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391
+ br_0_391 bl_0_392 br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394
+ bl_0_395 br_0_395 bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398
+ br_0_398 bl_0_399 br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401
+ bl_0_402 br_0_402 bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405
+ br_0_405 bl_0_406 br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408
+ bl_0_409 br_0_409 bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412
+ br_0_412 bl_0_413 br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415
+ bl_0_416 br_0_416 bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419
+ br_0_419 bl_0_420 br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422
+ bl_0_423 br_0_423 bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426
+ br_0_426 bl_0_427 br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429
+ bl_0_430 br_0_430 bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433
+ br_0_433 bl_0_434 br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436
+ bl_0_437 br_0_437 bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440
+ br_0_440 bl_0_441 br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443
+ bl_0_444 br_0_444 bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447
+ br_0_447 bl_0_448 br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450
+ bl_0_451 br_0_451 bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454
+ br_0_454 bl_0_455 br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457
+ bl_0_458 br_0_458 bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461
+ br_0_461 bl_0_462 br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464
+ bl_0_465 br_0_465 bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468
+ br_0_468 bl_0_469 br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471
+ bl_0_472 br_0_472 bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475
+ br_0_475 bl_0_476 br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478
+ bl_0_479 br_0_479 bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482
+ br_0_482 bl_0_483 br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485
+ bl_0_486 br_0_486 bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489
+ br_0_489 bl_0_490 br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492
+ bl_0_493 br_0_493 bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496
+ br_0_496 bl_0_497 br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499
+ bl_0_500 br_0_500 bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503
+ br_0_503 bl_0_504 br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506
+ bl_0_507 br_0_507 bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510
+ br_0_510 bl_0_511 br_0_511 rbl_wl0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4
+ wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13
+ wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21
+ wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37
+ wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 vdd gnd
+ freepdk45_sram_1rw0r_45x512_capped_replica_bitcell_array
Xport_data0
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 bl_0_256 br_0_256 bl_0_257 br_0_257 bl_0_258
+ br_0_258 bl_0_259 br_0_259 bl_0_260 br_0_260 bl_0_261 br_0_261
+ bl_0_262 br_0_262 bl_0_263 br_0_263 bl_0_264 br_0_264 bl_0_265
+ br_0_265 bl_0_266 br_0_266 bl_0_267 br_0_267 bl_0_268 br_0_268
+ bl_0_269 br_0_269 bl_0_270 br_0_270 bl_0_271 br_0_271 bl_0_272
+ br_0_272 bl_0_273 br_0_273 bl_0_274 br_0_274 bl_0_275 br_0_275
+ bl_0_276 br_0_276 bl_0_277 br_0_277 bl_0_278 br_0_278 bl_0_279
+ br_0_279 bl_0_280 br_0_280 bl_0_281 br_0_281 bl_0_282 br_0_282
+ bl_0_283 br_0_283 bl_0_284 br_0_284 bl_0_285 br_0_285 bl_0_286
+ br_0_286 bl_0_287 br_0_287 bl_0_288 br_0_288 bl_0_289 br_0_289
+ bl_0_290 br_0_290 bl_0_291 br_0_291 bl_0_292 br_0_292 bl_0_293
+ br_0_293 bl_0_294 br_0_294 bl_0_295 br_0_295 bl_0_296 br_0_296
+ bl_0_297 br_0_297 bl_0_298 br_0_298 bl_0_299 br_0_299 bl_0_300
+ br_0_300 bl_0_301 br_0_301 bl_0_302 br_0_302 bl_0_303 br_0_303
+ bl_0_304 br_0_304 bl_0_305 br_0_305 bl_0_306 br_0_306 bl_0_307
+ br_0_307 bl_0_308 br_0_308 bl_0_309 br_0_309 bl_0_310 br_0_310
+ bl_0_311 br_0_311 bl_0_312 br_0_312 bl_0_313 br_0_313 bl_0_314
+ br_0_314 bl_0_315 br_0_315 bl_0_316 br_0_316 bl_0_317 br_0_317
+ bl_0_318 br_0_318 bl_0_319 br_0_319 bl_0_320 br_0_320 bl_0_321
+ br_0_321 bl_0_322 br_0_322 bl_0_323 br_0_323 bl_0_324 br_0_324
+ bl_0_325 br_0_325 bl_0_326 br_0_326 bl_0_327 br_0_327 bl_0_328
+ br_0_328 bl_0_329 br_0_329 bl_0_330 br_0_330 bl_0_331 br_0_331
+ bl_0_332 br_0_332 bl_0_333 br_0_333 bl_0_334 br_0_334 bl_0_335
+ br_0_335 bl_0_336 br_0_336 bl_0_337 br_0_337 bl_0_338 br_0_338
+ bl_0_339 br_0_339 bl_0_340 br_0_340 bl_0_341 br_0_341 bl_0_342
+ br_0_342 bl_0_343 br_0_343 bl_0_344 br_0_344 bl_0_345 br_0_345
+ bl_0_346 br_0_346 bl_0_347 br_0_347 bl_0_348 br_0_348 bl_0_349
+ br_0_349 bl_0_350 br_0_350 bl_0_351 br_0_351 bl_0_352 br_0_352
+ bl_0_353 br_0_353 bl_0_354 br_0_354 bl_0_355 br_0_355 bl_0_356
+ br_0_356 bl_0_357 br_0_357 bl_0_358 br_0_358 bl_0_359 br_0_359
+ bl_0_360 br_0_360 bl_0_361 br_0_361 bl_0_362 br_0_362 bl_0_363
+ br_0_363 bl_0_364 br_0_364 bl_0_365 br_0_365 bl_0_366 br_0_366
+ bl_0_367 br_0_367 bl_0_368 br_0_368 bl_0_369 br_0_369 bl_0_370
+ br_0_370 bl_0_371 br_0_371 bl_0_372 br_0_372 bl_0_373 br_0_373
+ bl_0_374 br_0_374 bl_0_375 br_0_375 bl_0_376 br_0_376 bl_0_377
+ br_0_377 bl_0_378 br_0_378 bl_0_379 br_0_379 bl_0_380 br_0_380
+ bl_0_381 br_0_381 bl_0_382 br_0_382 bl_0_383 br_0_383 bl_0_384
+ br_0_384 bl_0_385 br_0_385 bl_0_386 br_0_386 bl_0_387 br_0_387
+ bl_0_388 br_0_388 bl_0_389 br_0_389 bl_0_390 br_0_390 bl_0_391
+ br_0_391 bl_0_392 br_0_392 bl_0_393 br_0_393 bl_0_394 br_0_394
+ bl_0_395 br_0_395 bl_0_396 br_0_396 bl_0_397 br_0_397 bl_0_398
+ br_0_398 bl_0_399 br_0_399 bl_0_400 br_0_400 bl_0_401 br_0_401
+ bl_0_402 br_0_402 bl_0_403 br_0_403 bl_0_404 br_0_404 bl_0_405
+ br_0_405 bl_0_406 br_0_406 bl_0_407 br_0_407 bl_0_408 br_0_408
+ bl_0_409 br_0_409 bl_0_410 br_0_410 bl_0_411 br_0_411 bl_0_412
+ br_0_412 bl_0_413 br_0_413 bl_0_414 br_0_414 bl_0_415 br_0_415
+ bl_0_416 br_0_416 bl_0_417 br_0_417 bl_0_418 br_0_418 bl_0_419
+ br_0_419 bl_0_420 br_0_420 bl_0_421 br_0_421 bl_0_422 br_0_422
+ bl_0_423 br_0_423 bl_0_424 br_0_424 bl_0_425 br_0_425 bl_0_426
+ br_0_426 bl_0_427 br_0_427 bl_0_428 br_0_428 bl_0_429 br_0_429
+ bl_0_430 br_0_430 bl_0_431 br_0_431 bl_0_432 br_0_432 bl_0_433
+ br_0_433 bl_0_434 br_0_434 bl_0_435 br_0_435 bl_0_436 br_0_436
+ bl_0_437 br_0_437 bl_0_438 br_0_438 bl_0_439 br_0_439 bl_0_440
+ br_0_440 bl_0_441 br_0_441 bl_0_442 br_0_442 bl_0_443 br_0_443
+ bl_0_444 br_0_444 bl_0_445 br_0_445 bl_0_446 br_0_446 bl_0_447
+ br_0_447 bl_0_448 br_0_448 bl_0_449 br_0_449 bl_0_450 br_0_450
+ bl_0_451 br_0_451 bl_0_452 br_0_452 bl_0_453 br_0_453 bl_0_454
+ br_0_454 bl_0_455 br_0_455 bl_0_456 br_0_456 bl_0_457 br_0_457
+ bl_0_458 br_0_458 bl_0_459 br_0_459 bl_0_460 br_0_460 bl_0_461
+ br_0_461 bl_0_462 br_0_462 bl_0_463 br_0_463 bl_0_464 br_0_464
+ bl_0_465 br_0_465 bl_0_466 br_0_466 bl_0_467 br_0_467 bl_0_468
+ br_0_468 bl_0_469 br_0_469 bl_0_470 br_0_470 bl_0_471 br_0_471
+ bl_0_472 br_0_472 bl_0_473 br_0_473 bl_0_474 br_0_474 bl_0_475
+ br_0_475 bl_0_476 br_0_476 bl_0_477 br_0_477 bl_0_478 br_0_478
+ bl_0_479 br_0_479 bl_0_480 br_0_480 bl_0_481 br_0_481 bl_0_482
+ br_0_482 bl_0_483 br_0_483 bl_0_484 br_0_484 bl_0_485 br_0_485
+ bl_0_486 br_0_486 bl_0_487 br_0_487 bl_0_488 br_0_488 bl_0_489
+ br_0_489 bl_0_490 br_0_490 bl_0_491 br_0_491 bl_0_492 br_0_492
+ bl_0_493 br_0_493 bl_0_494 br_0_494 bl_0_495 br_0_495 bl_0_496
+ br_0_496 bl_0_497 br_0_497 bl_0_498 br_0_498 bl_0_499 br_0_499
+ bl_0_500 br_0_500 bl_0_501 br_0_501 bl_0_502 br_0_502 bl_0_503
+ br_0_503 bl_0_504 br_0_504 bl_0_505 br_0_505 bl_0_506 br_0_506
+ bl_0_507 br_0_507 bl_0_508 br_0_508 bl_0_509 br_0_509 bl_0_510
+ br_0_510 bl_0_511 br_0_511 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4
+ dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12
+ dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19
+ dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26
+ dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout0_32 dout0_33
+ dout0_34 dout0_35 dout0_36 dout0_37 dout0_38 dout0_39 dout0_40
+ dout0_41 dout0_42 dout0_43 dout0_44 dout0_45 dout0_46 dout0_47
+ dout0_48 dout0_49 dout0_50 dout0_51 dout0_52 dout0_53 dout0_54
+ dout0_55 dout0_56 dout0_57 dout0_58 dout0_59 dout0_60 dout0_61
+ dout0_62 dout0_63 dout0_64 dout0_65 dout0_66 dout0_67 dout0_68
+ dout0_69 dout0_70 dout0_71 dout0_72 dout0_73 dout0_74 dout0_75
+ dout0_76 dout0_77 dout0_78 dout0_79 dout0_80 dout0_81 dout0_82
+ dout0_83 dout0_84 dout0_85 dout0_86 dout0_87 dout0_88 dout0_89
+ dout0_90 dout0_91 dout0_92 dout0_93 dout0_94 dout0_95 dout0_96
+ dout0_97 dout0_98 dout0_99 dout0_100 dout0_101 dout0_102 dout0_103
+ dout0_104 dout0_105 dout0_106 dout0_107 dout0_108 dout0_109 dout0_110
+ dout0_111 dout0_112 dout0_113 dout0_114 dout0_115 dout0_116 dout0_117
+ dout0_118 dout0_119 dout0_120 dout0_121 dout0_122 dout0_123 dout0_124
+ dout0_125 dout0_126 dout0_127 dout0_128 dout0_129 dout0_130 dout0_131
+ dout0_132 dout0_133 dout0_134 dout0_135 dout0_136 dout0_137 dout0_138
+ dout0_139 dout0_140 dout0_141 dout0_142 dout0_143 dout0_144 dout0_145
+ dout0_146 dout0_147 dout0_148 dout0_149 dout0_150 dout0_151 dout0_152
+ dout0_153 dout0_154 dout0_155 dout0_156 dout0_157 dout0_158 dout0_159
+ dout0_160 dout0_161 dout0_162 dout0_163 dout0_164 dout0_165 dout0_166
+ dout0_167 dout0_168 dout0_169 dout0_170 dout0_171 dout0_172 dout0_173
+ dout0_174 dout0_175 dout0_176 dout0_177 dout0_178 dout0_179 dout0_180
+ dout0_181 dout0_182 dout0_183 dout0_184 dout0_185 dout0_186 dout0_187
+ dout0_188 dout0_189 dout0_190 dout0_191 dout0_192 dout0_193 dout0_194
+ dout0_195 dout0_196 dout0_197 dout0_198 dout0_199 dout0_200 dout0_201
+ dout0_202 dout0_203 dout0_204 dout0_205 dout0_206 dout0_207 dout0_208
+ dout0_209 dout0_210 dout0_211 dout0_212 dout0_213 dout0_214 dout0_215
+ dout0_216 dout0_217 dout0_218 dout0_219 dout0_220 dout0_221 dout0_222
+ dout0_223 dout0_224 dout0_225 dout0_226 dout0_227 dout0_228 dout0_229
+ dout0_230 dout0_231 dout0_232 dout0_233 dout0_234 dout0_235 dout0_236
+ dout0_237 dout0_238 dout0_239 dout0_240 dout0_241 dout0_242 dout0_243
+ dout0_244 dout0_245 dout0_246 dout0_247 dout0_248 dout0_249 dout0_250
+ dout0_251 dout0_252 dout0_253 dout0_254 dout0_255 dout0_256 dout0_257
+ dout0_258 dout0_259 dout0_260 dout0_261 dout0_262 dout0_263 dout0_264
+ dout0_265 dout0_266 dout0_267 dout0_268 dout0_269 dout0_270 dout0_271
+ dout0_272 dout0_273 dout0_274 dout0_275 dout0_276 dout0_277 dout0_278
+ dout0_279 dout0_280 dout0_281 dout0_282 dout0_283 dout0_284 dout0_285
+ dout0_286 dout0_287 dout0_288 dout0_289 dout0_290 dout0_291 dout0_292
+ dout0_293 dout0_294 dout0_295 dout0_296 dout0_297 dout0_298 dout0_299
+ dout0_300 dout0_301 dout0_302 dout0_303 dout0_304 dout0_305 dout0_306
+ dout0_307 dout0_308 dout0_309 dout0_310 dout0_311 dout0_312 dout0_313
+ dout0_314 dout0_315 dout0_316 dout0_317 dout0_318 dout0_319 dout0_320
+ dout0_321 dout0_322 dout0_323 dout0_324 dout0_325 dout0_326 dout0_327
+ dout0_328 dout0_329 dout0_330 dout0_331 dout0_332 dout0_333 dout0_334
+ dout0_335 dout0_336 dout0_337 dout0_338 dout0_339 dout0_340 dout0_341
+ dout0_342 dout0_343 dout0_344 dout0_345 dout0_346 dout0_347 dout0_348
+ dout0_349 dout0_350 dout0_351 dout0_352 dout0_353 dout0_354 dout0_355
+ dout0_356 dout0_357 dout0_358 dout0_359 dout0_360 dout0_361 dout0_362
+ dout0_363 dout0_364 dout0_365 dout0_366 dout0_367 dout0_368 dout0_369
+ dout0_370 dout0_371 dout0_372 dout0_373 dout0_374 dout0_375 dout0_376
+ dout0_377 dout0_378 dout0_379 dout0_380 dout0_381 dout0_382 dout0_383
+ dout0_384 dout0_385 dout0_386 dout0_387 dout0_388 dout0_389 dout0_390
+ dout0_391 dout0_392 dout0_393 dout0_394 dout0_395 dout0_396 dout0_397
+ dout0_398 dout0_399 dout0_400 dout0_401 dout0_402 dout0_403 dout0_404
+ dout0_405 dout0_406 dout0_407 dout0_408 dout0_409 dout0_410 dout0_411
+ dout0_412 dout0_413 dout0_414 dout0_415 dout0_416 dout0_417 dout0_418
+ dout0_419 dout0_420 dout0_421 dout0_422 dout0_423 dout0_424 dout0_425
+ dout0_426 dout0_427 dout0_428 dout0_429 dout0_430 dout0_431 dout0_432
+ dout0_433 dout0_434 dout0_435 dout0_436 dout0_437 dout0_438 dout0_439
+ dout0_440 dout0_441 dout0_442 dout0_443 dout0_444 dout0_445 dout0_446
+ dout0_447 dout0_448 dout0_449 dout0_450 dout0_451 dout0_452 dout0_453
+ dout0_454 dout0_455 dout0_456 dout0_457 dout0_458 dout0_459 dout0_460
+ dout0_461 dout0_462 dout0_463 dout0_464 dout0_465 dout0_466 dout0_467
+ dout0_468 dout0_469 dout0_470 dout0_471 dout0_472 dout0_473 dout0_474
+ dout0_475 dout0_476 dout0_477 dout0_478 dout0_479 dout0_480 dout0_481
+ dout0_482 dout0_483 dout0_484 dout0_485 dout0_486 dout0_487 dout0_488
+ dout0_489 dout0_490 dout0_491 dout0_492 dout0_493 dout0_494 dout0_495
+ dout0_496 dout0_497 dout0_498 dout0_499 dout0_500 dout0_501 dout0_502
+ dout0_503 dout0_504 dout0_505 dout0_506 dout0_507 dout0_508 dout0_509
+ dout0_510 dout0_511 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6
+ din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15
+ din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23
+ din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31
+ din0_32 din0_33 din0_34 din0_35 din0_36 din0_37 din0_38 din0_39
+ din0_40 din0_41 din0_42 din0_43 din0_44 din0_45 din0_46 din0_47
+ din0_48 din0_49 din0_50 din0_51 din0_52 din0_53 din0_54 din0_55
+ din0_56 din0_57 din0_58 din0_59 din0_60 din0_61 din0_62 din0_63
+ din0_64 din0_65 din0_66 din0_67 din0_68 din0_69 din0_70 din0_71
+ din0_72 din0_73 din0_74 din0_75 din0_76 din0_77 din0_78 din0_79
+ din0_80 din0_81 din0_82 din0_83 din0_84 din0_85 din0_86 din0_87
+ din0_88 din0_89 din0_90 din0_91 din0_92 din0_93 din0_94 din0_95
+ din0_96 din0_97 din0_98 din0_99 din0_100 din0_101 din0_102 din0_103
+ din0_104 din0_105 din0_106 din0_107 din0_108 din0_109 din0_110
+ din0_111 din0_112 din0_113 din0_114 din0_115 din0_116 din0_117
+ din0_118 din0_119 din0_120 din0_121 din0_122 din0_123 din0_124
+ din0_125 din0_126 din0_127 din0_128 din0_129 din0_130 din0_131
+ din0_132 din0_133 din0_134 din0_135 din0_136 din0_137 din0_138
+ din0_139 din0_140 din0_141 din0_142 din0_143 din0_144 din0_145
+ din0_146 din0_147 din0_148 din0_149 din0_150 din0_151 din0_152
+ din0_153 din0_154 din0_155 din0_156 din0_157 din0_158 din0_159
+ din0_160 din0_161 din0_162 din0_163 din0_164 din0_165 din0_166
+ din0_167 din0_168 din0_169 din0_170 din0_171 din0_172 din0_173
+ din0_174 din0_175 din0_176 din0_177 din0_178 din0_179 din0_180
+ din0_181 din0_182 din0_183 din0_184 din0_185 din0_186 din0_187
+ din0_188 din0_189 din0_190 din0_191 din0_192 din0_193 din0_194
+ din0_195 din0_196 din0_197 din0_198 din0_199 din0_200 din0_201
+ din0_202 din0_203 din0_204 din0_205 din0_206 din0_207 din0_208
+ din0_209 din0_210 din0_211 din0_212 din0_213 din0_214 din0_215
+ din0_216 din0_217 din0_218 din0_219 din0_220 din0_221 din0_222
+ din0_223 din0_224 din0_225 din0_226 din0_227 din0_228 din0_229
+ din0_230 din0_231 din0_232 din0_233 din0_234 din0_235 din0_236
+ din0_237 din0_238 din0_239 din0_240 din0_241 din0_242 din0_243
+ din0_244 din0_245 din0_246 din0_247 din0_248 din0_249 din0_250
+ din0_251 din0_252 din0_253 din0_254 din0_255 din0_256 din0_257
+ din0_258 din0_259 din0_260 din0_261 din0_262 din0_263 din0_264
+ din0_265 din0_266 din0_267 din0_268 din0_269 din0_270 din0_271
+ din0_272 din0_273 din0_274 din0_275 din0_276 din0_277 din0_278
+ din0_279 din0_280 din0_281 din0_282 din0_283 din0_284 din0_285
+ din0_286 din0_287 din0_288 din0_289 din0_290 din0_291 din0_292
+ din0_293 din0_294 din0_295 din0_296 din0_297 din0_298 din0_299
+ din0_300 din0_301 din0_302 din0_303 din0_304 din0_305 din0_306
+ din0_307 din0_308 din0_309 din0_310 din0_311 din0_312 din0_313
+ din0_314 din0_315 din0_316 din0_317 din0_318 din0_319 din0_320
+ din0_321 din0_322 din0_323 din0_324 din0_325 din0_326 din0_327
+ din0_328 din0_329 din0_330 din0_331 din0_332 din0_333 din0_334
+ din0_335 din0_336 din0_337 din0_338 din0_339 din0_340 din0_341
+ din0_342 din0_343 din0_344 din0_345 din0_346 din0_347 din0_348
+ din0_349 din0_350 din0_351 din0_352 din0_353 din0_354 din0_355
+ din0_356 din0_357 din0_358 din0_359 din0_360 din0_361 din0_362
+ din0_363 din0_364 din0_365 din0_366 din0_367 din0_368 din0_369
+ din0_370 din0_371 din0_372 din0_373 din0_374 din0_375 din0_376
+ din0_377 din0_378 din0_379 din0_380 din0_381 din0_382 din0_383
+ din0_384 din0_385 din0_386 din0_387 din0_388 din0_389 din0_390
+ din0_391 din0_392 din0_393 din0_394 din0_395 din0_396 din0_397
+ din0_398 din0_399 din0_400 din0_401 din0_402 din0_403 din0_404
+ din0_405 din0_406 din0_407 din0_408 din0_409 din0_410 din0_411
+ din0_412 din0_413 din0_414 din0_415 din0_416 din0_417 din0_418
+ din0_419 din0_420 din0_421 din0_422 din0_423 din0_424 din0_425
+ din0_426 din0_427 din0_428 din0_429 din0_430 din0_431 din0_432
+ din0_433 din0_434 din0_435 din0_436 din0_437 din0_438 din0_439
+ din0_440 din0_441 din0_442 din0_443 din0_444 din0_445 din0_446
+ din0_447 din0_448 din0_449 din0_450 din0_451 din0_452 din0_453
+ din0_454 din0_455 din0_456 din0_457 din0_458 din0_459 din0_460
+ din0_461 din0_462 din0_463 din0_464 din0_465 din0_466 din0_467
+ din0_468 din0_469 din0_470 din0_471 din0_472 din0_473 din0_474
+ din0_475 din0_476 din0_477 din0_478 din0_479 din0_480 din0_481
+ din0_482 din0_483 din0_484 din0_485 din0_486 din0_487 din0_488
+ din0_489 din0_490 din0_491 din0_492 din0_493 din0_494 din0_495
+ din0_496 din0_497 din0_498 din0_499 din0_500 din0_501 din0_502
+ din0_503 din0_504 din0_505 din0_506 din0_507 din0_508 din0_509
+ din0_510 din0_511 s_en0 p_en_bar0 w_en0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_port_data
Xport_address0
+ addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 wl_en0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 rbl_wl0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_port_address
.ENDS freepdk45_sram_1rw0r_45x512_bank

.SUBCKT freepdk45_sram_1rw0r_45x512
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22]
+ din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29]
+ din0[30] din0[31] din0[32] din0[33] din0[34] din0[35] din0[36]
+ din0[37] din0[38] din0[39] din0[40] din0[41] din0[42] din0[43]
+ din0[44] din0[45] din0[46] din0[47] din0[48] din0[49] din0[50]
+ din0[51] din0[52] din0[53] din0[54] din0[55] din0[56] din0[57]
+ din0[58] din0[59] din0[60] din0[61] din0[62] din0[63] din0[64]
+ din0[65] din0[66] din0[67] din0[68] din0[69] din0[70] din0[71]
+ din0[72] din0[73] din0[74] din0[75] din0[76] din0[77] din0[78]
+ din0[79] din0[80] din0[81] din0[82] din0[83] din0[84] din0[85]
+ din0[86] din0[87] din0[88] din0[89] din0[90] din0[91] din0[92]
+ din0[93] din0[94] din0[95] din0[96] din0[97] din0[98] din0[99]
+ din0[100] din0[101] din0[102] din0[103] din0[104] din0[105] din0[106]
+ din0[107] din0[108] din0[109] din0[110] din0[111] din0[112] din0[113]
+ din0[114] din0[115] din0[116] din0[117] din0[118] din0[119] din0[120]
+ din0[121] din0[122] din0[123] din0[124] din0[125] din0[126] din0[127]
+ din0[128] din0[129] din0[130] din0[131] din0[132] din0[133] din0[134]
+ din0[135] din0[136] din0[137] din0[138] din0[139] din0[140] din0[141]
+ din0[142] din0[143] din0[144] din0[145] din0[146] din0[147] din0[148]
+ din0[149] din0[150] din0[151] din0[152] din0[153] din0[154] din0[155]
+ din0[156] din0[157] din0[158] din0[159] din0[160] din0[161] din0[162]
+ din0[163] din0[164] din0[165] din0[166] din0[167] din0[168] din0[169]
+ din0[170] din0[171] din0[172] din0[173] din0[174] din0[175] din0[176]
+ din0[177] din0[178] din0[179] din0[180] din0[181] din0[182] din0[183]
+ din0[184] din0[185] din0[186] din0[187] din0[188] din0[189] din0[190]
+ din0[191] din0[192] din0[193] din0[194] din0[195] din0[196] din0[197]
+ din0[198] din0[199] din0[200] din0[201] din0[202] din0[203] din0[204]
+ din0[205] din0[206] din0[207] din0[208] din0[209] din0[210] din0[211]
+ din0[212] din0[213] din0[214] din0[215] din0[216] din0[217] din0[218]
+ din0[219] din0[220] din0[221] din0[222] din0[223] din0[224] din0[225]
+ din0[226] din0[227] din0[228] din0[229] din0[230] din0[231] din0[232]
+ din0[233] din0[234] din0[235] din0[236] din0[237] din0[238] din0[239]
+ din0[240] din0[241] din0[242] din0[243] din0[244] din0[245] din0[246]
+ din0[247] din0[248] din0[249] din0[250] din0[251] din0[252] din0[253]
+ din0[254] din0[255] din0[256] din0[257] din0[258] din0[259] din0[260]
+ din0[261] din0[262] din0[263] din0[264] din0[265] din0[266] din0[267]
+ din0[268] din0[269] din0[270] din0[271] din0[272] din0[273] din0[274]
+ din0[275] din0[276] din0[277] din0[278] din0[279] din0[280] din0[281]
+ din0[282] din0[283] din0[284] din0[285] din0[286] din0[287] din0[288]
+ din0[289] din0[290] din0[291] din0[292] din0[293] din0[294] din0[295]
+ din0[296] din0[297] din0[298] din0[299] din0[300] din0[301] din0[302]
+ din0[303] din0[304] din0[305] din0[306] din0[307] din0[308] din0[309]
+ din0[310] din0[311] din0[312] din0[313] din0[314] din0[315] din0[316]
+ din0[317] din0[318] din0[319] din0[320] din0[321] din0[322] din0[323]
+ din0[324] din0[325] din0[326] din0[327] din0[328] din0[329] din0[330]
+ din0[331] din0[332] din0[333] din0[334] din0[335] din0[336] din0[337]
+ din0[338] din0[339] din0[340] din0[341] din0[342] din0[343] din0[344]
+ din0[345] din0[346] din0[347] din0[348] din0[349] din0[350] din0[351]
+ din0[352] din0[353] din0[354] din0[355] din0[356] din0[357] din0[358]
+ din0[359] din0[360] din0[361] din0[362] din0[363] din0[364] din0[365]
+ din0[366] din0[367] din0[368] din0[369] din0[370] din0[371] din0[372]
+ din0[373] din0[374] din0[375] din0[376] din0[377] din0[378] din0[379]
+ din0[380] din0[381] din0[382] din0[383] din0[384] din0[385] din0[386]
+ din0[387] din0[388] din0[389] din0[390] din0[391] din0[392] din0[393]
+ din0[394] din0[395] din0[396] din0[397] din0[398] din0[399] din0[400]
+ din0[401] din0[402] din0[403] din0[404] din0[405] din0[406] din0[407]
+ din0[408] din0[409] din0[410] din0[411] din0[412] din0[413] din0[414]
+ din0[415] din0[416] din0[417] din0[418] din0[419] din0[420] din0[421]
+ din0[422] din0[423] din0[424] din0[425] din0[426] din0[427] din0[428]
+ din0[429] din0[430] din0[431] din0[432] din0[433] din0[434] din0[435]
+ din0[436] din0[437] din0[438] din0[439] din0[440] din0[441] din0[442]
+ din0[443] din0[444] din0[445] din0[446] din0[447] din0[448] din0[449]
+ din0[450] din0[451] din0[452] din0[453] din0[454] din0[455] din0[456]
+ din0[457] din0[458] din0[459] din0[460] din0[461] din0[462] din0[463]
+ din0[464] din0[465] din0[466] din0[467] din0[468] din0[469] din0[470]
+ din0[471] din0[472] din0[473] din0[474] din0[475] din0[476] din0[477]
+ din0[478] din0[479] din0[480] din0[481] din0[482] din0[483] din0[484]
+ din0[485] din0[486] din0[487] din0[488] din0[489] din0[490] din0[491]
+ din0[492] din0[493] din0[494] din0[495] din0[496] din0[497] din0[498]
+ din0[499] din0[500] din0[501] din0[502] din0[503] din0[504] din0[505]
+ din0[506] din0[507] din0[508] din0[509] din0[510] din0[511] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] csb0 web0 clk0 dout0[0]
+ dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7]
+ dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14]
+ dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21]
+ dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28]
+ dout0[29] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35]
+ dout0[36] dout0[37] dout0[38] dout0[39] dout0[40] dout0[41] dout0[42]
+ dout0[43] dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49]
+ dout0[50] dout0[51] dout0[52] dout0[53] dout0[54] dout0[55] dout0[56]
+ dout0[57] dout0[58] dout0[59] dout0[60] dout0[61] dout0[62] dout0[63]
+ dout0[64] dout0[65] dout0[66] dout0[67] dout0[68] dout0[69] dout0[70]
+ dout0[71] dout0[72] dout0[73] dout0[74] dout0[75] dout0[76] dout0[77]
+ dout0[78] dout0[79] dout0[80] dout0[81] dout0[82] dout0[83] dout0[84]
+ dout0[85] dout0[86] dout0[87] dout0[88] dout0[89] dout0[90] dout0[91]
+ dout0[92] dout0[93] dout0[94] dout0[95] dout0[96] dout0[97] dout0[98]
+ dout0[99] dout0[100] dout0[101] dout0[102] dout0[103] dout0[104]
+ dout0[105] dout0[106] dout0[107] dout0[108] dout0[109] dout0[110]
+ dout0[111] dout0[112] dout0[113] dout0[114] dout0[115] dout0[116]
+ dout0[117] dout0[118] dout0[119] dout0[120] dout0[121] dout0[122]
+ dout0[123] dout0[124] dout0[125] dout0[126] dout0[127] dout0[128]
+ dout0[129] dout0[130] dout0[131] dout0[132] dout0[133] dout0[134]
+ dout0[135] dout0[136] dout0[137] dout0[138] dout0[139] dout0[140]
+ dout0[141] dout0[142] dout0[143] dout0[144] dout0[145] dout0[146]
+ dout0[147] dout0[148] dout0[149] dout0[150] dout0[151] dout0[152]
+ dout0[153] dout0[154] dout0[155] dout0[156] dout0[157] dout0[158]
+ dout0[159] dout0[160] dout0[161] dout0[162] dout0[163] dout0[164]
+ dout0[165] dout0[166] dout0[167] dout0[168] dout0[169] dout0[170]
+ dout0[171] dout0[172] dout0[173] dout0[174] dout0[175] dout0[176]
+ dout0[177] dout0[178] dout0[179] dout0[180] dout0[181] dout0[182]
+ dout0[183] dout0[184] dout0[185] dout0[186] dout0[187] dout0[188]
+ dout0[189] dout0[190] dout0[191] dout0[192] dout0[193] dout0[194]
+ dout0[195] dout0[196] dout0[197] dout0[198] dout0[199] dout0[200]
+ dout0[201] dout0[202] dout0[203] dout0[204] dout0[205] dout0[206]
+ dout0[207] dout0[208] dout0[209] dout0[210] dout0[211] dout0[212]
+ dout0[213] dout0[214] dout0[215] dout0[216] dout0[217] dout0[218]
+ dout0[219] dout0[220] dout0[221] dout0[222] dout0[223] dout0[224]
+ dout0[225] dout0[226] dout0[227] dout0[228] dout0[229] dout0[230]
+ dout0[231] dout0[232] dout0[233] dout0[234] dout0[235] dout0[236]
+ dout0[237] dout0[238] dout0[239] dout0[240] dout0[241] dout0[242]
+ dout0[243] dout0[244] dout0[245] dout0[246] dout0[247] dout0[248]
+ dout0[249] dout0[250] dout0[251] dout0[252] dout0[253] dout0[254]
+ dout0[255] dout0[256] dout0[257] dout0[258] dout0[259] dout0[260]
+ dout0[261] dout0[262] dout0[263] dout0[264] dout0[265] dout0[266]
+ dout0[267] dout0[268] dout0[269] dout0[270] dout0[271] dout0[272]
+ dout0[273] dout0[274] dout0[275] dout0[276] dout0[277] dout0[278]
+ dout0[279] dout0[280] dout0[281] dout0[282] dout0[283] dout0[284]
+ dout0[285] dout0[286] dout0[287] dout0[288] dout0[289] dout0[290]
+ dout0[291] dout0[292] dout0[293] dout0[294] dout0[295] dout0[296]
+ dout0[297] dout0[298] dout0[299] dout0[300] dout0[301] dout0[302]
+ dout0[303] dout0[304] dout0[305] dout0[306] dout0[307] dout0[308]
+ dout0[309] dout0[310] dout0[311] dout0[312] dout0[313] dout0[314]
+ dout0[315] dout0[316] dout0[317] dout0[318] dout0[319] dout0[320]
+ dout0[321] dout0[322] dout0[323] dout0[324] dout0[325] dout0[326]
+ dout0[327] dout0[328] dout0[329] dout0[330] dout0[331] dout0[332]
+ dout0[333] dout0[334] dout0[335] dout0[336] dout0[337] dout0[338]
+ dout0[339] dout0[340] dout0[341] dout0[342] dout0[343] dout0[344]
+ dout0[345] dout0[346] dout0[347] dout0[348] dout0[349] dout0[350]
+ dout0[351] dout0[352] dout0[353] dout0[354] dout0[355] dout0[356]
+ dout0[357] dout0[358] dout0[359] dout0[360] dout0[361] dout0[362]
+ dout0[363] dout0[364] dout0[365] dout0[366] dout0[367] dout0[368]
+ dout0[369] dout0[370] dout0[371] dout0[372] dout0[373] dout0[374]
+ dout0[375] dout0[376] dout0[377] dout0[378] dout0[379] dout0[380]
+ dout0[381] dout0[382] dout0[383] dout0[384] dout0[385] dout0[386]
+ dout0[387] dout0[388] dout0[389] dout0[390] dout0[391] dout0[392]
+ dout0[393] dout0[394] dout0[395] dout0[396] dout0[397] dout0[398]
+ dout0[399] dout0[400] dout0[401] dout0[402] dout0[403] dout0[404]
+ dout0[405] dout0[406] dout0[407] dout0[408] dout0[409] dout0[410]
+ dout0[411] dout0[412] dout0[413] dout0[414] dout0[415] dout0[416]
+ dout0[417] dout0[418] dout0[419] dout0[420] dout0[421] dout0[422]
+ dout0[423] dout0[424] dout0[425] dout0[426] dout0[427] dout0[428]
+ dout0[429] dout0[430] dout0[431] dout0[432] dout0[433] dout0[434]
+ dout0[435] dout0[436] dout0[437] dout0[438] dout0[439] dout0[440]
+ dout0[441] dout0[442] dout0[443] dout0[444] dout0[445] dout0[446]
+ dout0[447] dout0[448] dout0[449] dout0[450] dout0[451] dout0[452]
+ dout0[453] dout0[454] dout0[455] dout0[456] dout0[457] dout0[458]
+ dout0[459] dout0[460] dout0[461] dout0[462] dout0[463] dout0[464]
+ dout0[465] dout0[466] dout0[467] dout0[468] dout0[469] dout0[470]
+ dout0[471] dout0[472] dout0[473] dout0[474] dout0[475] dout0[476]
+ dout0[477] dout0[478] dout0[479] dout0[480] dout0[481] dout0[482]
+ dout0[483] dout0[484] dout0[485] dout0[486] dout0[487] dout0[488]
+ dout0[489] dout0[490] dout0[491] dout0[492] dout0[493] dout0[494]
+ dout0[495] dout0[496] dout0[497] dout0[498] dout0[499] dout0[500]
+ dout0[501] dout0[502] dout0[503] dout0[504] dout0[505] dout0[506]
+ dout0[507] dout0[508] dout0[509] dout0[510] dout0[511] vdd gnd
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : din0[32] 
* INPUT : din0[33] 
* INPUT : din0[34] 
* INPUT : din0[35] 
* INPUT : din0[36] 
* INPUT : din0[37] 
* INPUT : din0[38] 
* INPUT : din0[39] 
* INPUT : din0[40] 
* INPUT : din0[41] 
* INPUT : din0[42] 
* INPUT : din0[43] 
* INPUT : din0[44] 
* INPUT : din0[45] 
* INPUT : din0[46] 
* INPUT : din0[47] 
* INPUT : din0[48] 
* INPUT : din0[49] 
* INPUT : din0[50] 
* INPUT : din0[51] 
* INPUT : din0[52] 
* INPUT : din0[53] 
* INPUT : din0[54] 
* INPUT : din0[55] 
* INPUT : din0[56] 
* INPUT : din0[57] 
* INPUT : din0[58] 
* INPUT : din0[59] 
* INPUT : din0[60] 
* INPUT : din0[61] 
* INPUT : din0[62] 
* INPUT : din0[63] 
* INPUT : din0[64] 
* INPUT : din0[65] 
* INPUT : din0[66] 
* INPUT : din0[67] 
* INPUT : din0[68] 
* INPUT : din0[69] 
* INPUT : din0[70] 
* INPUT : din0[71] 
* INPUT : din0[72] 
* INPUT : din0[73] 
* INPUT : din0[74] 
* INPUT : din0[75] 
* INPUT : din0[76] 
* INPUT : din0[77] 
* INPUT : din0[78] 
* INPUT : din0[79] 
* INPUT : din0[80] 
* INPUT : din0[81] 
* INPUT : din0[82] 
* INPUT : din0[83] 
* INPUT : din0[84] 
* INPUT : din0[85] 
* INPUT : din0[86] 
* INPUT : din0[87] 
* INPUT : din0[88] 
* INPUT : din0[89] 
* INPUT : din0[90] 
* INPUT : din0[91] 
* INPUT : din0[92] 
* INPUT : din0[93] 
* INPUT : din0[94] 
* INPUT : din0[95] 
* INPUT : din0[96] 
* INPUT : din0[97] 
* INPUT : din0[98] 
* INPUT : din0[99] 
* INPUT : din0[100] 
* INPUT : din0[101] 
* INPUT : din0[102] 
* INPUT : din0[103] 
* INPUT : din0[104] 
* INPUT : din0[105] 
* INPUT : din0[106] 
* INPUT : din0[107] 
* INPUT : din0[108] 
* INPUT : din0[109] 
* INPUT : din0[110] 
* INPUT : din0[111] 
* INPUT : din0[112] 
* INPUT : din0[113] 
* INPUT : din0[114] 
* INPUT : din0[115] 
* INPUT : din0[116] 
* INPUT : din0[117] 
* INPUT : din0[118] 
* INPUT : din0[119] 
* INPUT : din0[120] 
* INPUT : din0[121] 
* INPUT : din0[122] 
* INPUT : din0[123] 
* INPUT : din0[124] 
* INPUT : din0[125] 
* INPUT : din0[126] 
* INPUT : din0[127] 
* INPUT : din0[128] 
* INPUT : din0[129] 
* INPUT : din0[130] 
* INPUT : din0[131] 
* INPUT : din0[132] 
* INPUT : din0[133] 
* INPUT : din0[134] 
* INPUT : din0[135] 
* INPUT : din0[136] 
* INPUT : din0[137] 
* INPUT : din0[138] 
* INPUT : din0[139] 
* INPUT : din0[140] 
* INPUT : din0[141] 
* INPUT : din0[142] 
* INPUT : din0[143] 
* INPUT : din0[144] 
* INPUT : din0[145] 
* INPUT : din0[146] 
* INPUT : din0[147] 
* INPUT : din0[148] 
* INPUT : din0[149] 
* INPUT : din0[150] 
* INPUT : din0[151] 
* INPUT : din0[152] 
* INPUT : din0[153] 
* INPUT : din0[154] 
* INPUT : din0[155] 
* INPUT : din0[156] 
* INPUT : din0[157] 
* INPUT : din0[158] 
* INPUT : din0[159] 
* INPUT : din0[160] 
* INPUT : din0[161] 
* INPUT : din0[162] 
* INPUT : din0[163] 
* INPUT : din0[164] 
* INPUT : din0[165] 
* INPUT : din0[166] 
* INPUT : din0[167] 
* INPUT : din0[168] 
* INPUT : din0[169] 
* INPUT : din0[170] 
* INPUT : din0[171] 
* INPUT : din0[172] 
* INPUT : din0[173] 
* INPUT : din0[174] 
* INPUT : din0[175] 
* INPUT : din0[176] 
* INPUT : din0[177] 
* INPUT : din0[178] 
* INPUT : din0[179] 
* INPUT : din0[180] 
* INPUT : din0[181] 
* INPUT : din0[182] 
* INPUT : din0[183] 
* INPUT : din0[184] 
* INPUT : din0[185] 
* INPUT : din0[186] 
* INPUT : din0[187] 
* INPUT : din0[188] 
* INPUT : din0[189] 
* INPUT : din0[190] 
* INPUT : din0[191] 
* INPUT : din0[192] 
* INPUT : din0[193] 
* INPUT : din0[194] 
* INPUT : din0[195] 
* INPUT : din0[196] 
* INPUT : din0[197] 
* INPUT : din0[198] 
* INPUT : din0[199] 
* INPUT : din0[200] 
* INPUT : din0[201] 
* INPUT : din0[202] 
* INPUT : din0[203] 
* INPUT : din0[204] 
* INPUT : din0[205] 
* INPUT : din0[206] 
* INPUT : din0[207] 
* INPUT : din0[208] 
* INPUT : din0[209] 
* INPUT : din0[210] 
* INPUT : din0[211] 
* INPUT : din0[212] 
* INPUT : din0[213] 
* INPUT : din0[214] 
* INPUT : din0[215] 
* INPUT : din0[216] 
* INPUT : din0[217] 
* INPUT : din0[218] 
* INPUT : din0[219] 
* INPUT : din0[220] 
* INPUT : din0[221] 
* INPUT : din0[222] 
* INPUT : din0[223] 
* INPUT : din0[224] 
* INPUT : din0[225] 
* INPUT : din0[226] 
* INPUT : din0[227] 
* INPUT : din0[228] 
* INPUT : din0[229] 
* INPUT : din0[230] 
* INPUT : din0[231] 
* INPUT : din0[232] 
* INPUT : din0[233] 
* INPUT : din0[234] 
* INPUT : din0[235] 
* INPUT : din0[236] 
* INPUT : din0[237] 
* INPUT : din0[238] 
* INPUT : din0[239] 
* INPUT : din0[240] 
* INPUT : din0[241] 
* INPUT : din0[242] 
* INPUT : din0[243] 
* INPUT : din0[244] 
* INPUT : din0[245] 
* INPUT : din0[246] 
* INPUT : din0[247] 
* INPUT : din0[248] 
* INPUT : din0[249] 
* INPUT : din0[250] 
* INPUT : din0[251] 
* INPUT : din0[252] 
* INPUT : din0[253] 
* INPUT : din0[254] 
* INPUT : din0[255] 
* INPUT : din0[256] 
* INPUT : din0[257] 
* INPUT : din0[258] 
* INPUT : din0[259] 
* INPUT : din0[260] 
* INPUT : din0[261] 
* INPUT : din0[262] 
* INPUT : din0[263] 
* INPUT : din0[264] 
* INPUT : din0[265] 
* INPUT : din0[266] 
* INPUT : din0[267] 
* INPUT : din0[268] 
* INPUT : din0[269] 
* INPUT : din0[270] 
* INPUT : din0[271] 
* INPUT : din0[272] 
* INPUT : din0[273] 
* INPUT : din0[274] 
* INPUT : din0[275] 
* INPUT : din0[276] 
* INPUT : din0[277] 
* INPUT : din0[278] 
* INPUT : din0[279] 
* INPUT : din0[280] 
* INPUT : din0[281] 
* INPUT : din0[282] 
* INPUT : din0[283] 
* INPUT : din0[284] 
* INPUT : din0[285] 
* INPUT : din0[286] 
* INPUT : din0[287] 
* INPUT : din0[288] 
* INPUT : din0[289] 
* INPUT : din0[290] 
* INPUT : din0[291] 
* INPUT : din0[292] 
* INPUT : din0[293] 
* INPUT : din0[294] 
* INPUT : din0[295] 
* INPUT : din0[296] 
* INPUT : din0[297] 
* INPUT : din0[298] 
* INPUT : din0[299] 
* INPUT : din0[300] 
* INPUT : din0[301] 
* INPUT : din0[302] 
* INPUT : din0[303] 
* INPUT : din0[304] 
* INPUT : din0[305] 
* INPUT : din0[306] 
* INPUT : din0[307] 
* INPUT : din0[308] 
* INPUT : din0[309] 
* INPUT : din0[310] 
* INPUT : din0[311] 
* INPUT : din0[312] 
* INPUT : din0[313] 
* INPUT : din0[314] 
* INPUT : din0[315] 
* INPUT : din0[316] 
* INPUT : din0[317] 
* INPUT : din0[318] 
* INPUT : din0[319] 
* INPUT : din0[320] 
* INPUT : din0[321] 
* INPUT : din0[322] 
* INPUT : din0[323] 
* INPUT : din0[324] 
* INPUT : din0[325] 
* INPUT : din0[326] 
* INPUT : din0[327] 
* INPUT : din0[328] 
* INPUT : din0[329] 
* INPUT : din0[330] 
* INPUT : din0[331] 
* INPUT : din0[332] 
* INPUT : din0[333] 
* INPUT : din0[334] 
* INPUT : din0[335] 
* INPUT : din0[336] 
* INPUT : din0[337] 
* INPUT : din0[338] 
* INPUT : din0[339] 
* INPUT : din0[340] 
* INPUT : din0[341] 
* INPUT : din0[342] 
* INPUT : din0[343] 
* INPUT : din0[344] 
* INPUT : din0[345] 
* INPUT : din0[346] 
* INPUT : din0[347] 
* INPUT : din0[348] 
* INPUT : din0[349] 
* INPUT : din0[350] 
* INPUT : din0[351] 
* INPUT : din0[352] 
* INPUT : din0[353] 
* INPUT : din0[354] 
* INPUT : din0[355] 
* INPUT : din0[356] 
* INPUT : din0[357] 
* INPUT : din0[358] 
* INPUT : din0[359] 
* INPUT : din0[360] 
* INPUT : din0[361] 
* INPUT : din0[362] 
* INPUT : din0[363] 
* INPUT : din0[364] 
* INPUT : din0[365] 
* INPUT : din0[366] 
* INPUT : din0[367] 
* INPUT : din0[368] 
* INPUT : din0[369] 
* INPUT : din0[370] 
* INPUT : din0[371] 
* INPUT : din0[372] 
* INPUT : din0[373] 
* INPUT : din0[374] 
* INPUT : din0[375] 
* INPUT : din0[376] 
* INPUT : din0[377] 
* INPUT : din0[378] 
* INPUT : din0[379] 
* INPUT : din0[380] 
* INPUT : din0[381] 
* INPUT : din0[382] 
* INPUT : din0[383] 
* INPUT : din0[384] 
* INPUT : din0[385] 
* INPUT : din0[386] 
* INPUT : din0[387] 
* INPUT : din0[388] 
* INPUT : din0[389] 
* INPUT : din0[390] 
* INPUT : din0[391] 
* INPUT : din0[392] 
* INPUT : din0[393] 
* INPUT : din0[394] 
* INPUT : din0[395] 
* INPUT : din0[396] 
* INPUT : din0[397] 
* INPUT : din0[398] 
* INPUT : din0[399] 
* INPUT : din0[400] 
* INPUT : din0[401] 
* INPUT : din0[402] 
* INPUT : din0[403] 
* INPUT : din0[404] 
* INPUT : din0[405] 
* INPUT : din0[406] 
* INPUT : din0[407] 
* INPUT : din0[408] 
* INPUT : din0[409] 
* INPUT : din0[410] 
* INPUT : din0[411] 
* INPUT : din0[412] 
* INPUT : din0[413] 
* INPUT : din0[414] 
* INPUT : din0[415] 
* INPUT : din0[416] 
* INPUT : din0[417] 
* INPUT : din0[418] 
* INPUT : din0[419] 
* INPUT : din0[420] 
* INPUT : din0[421] 
* INPUT : din0[422] 
* INPUT : din0[423] 
* INPUT : din0[424] 
* INPUT : din0[425] 
* INPUT : din0[426] 
* INPUT : din0[427] 
* INPUT : din0[428] 
* INPUT : din0[429] 
* INPUT : din0[430] 
* INPUT : din0[431] 
* INPUT : din0[432] 
* INPUT : din0[433] 
* INPUT : din0[434] 
* INPUT : din0[435] 
* INPUT : din0[436] 
* INPUT : din0[437] 
* INPUT : din0[438] 
* INPUT : din0[439] 
* INPUT : din0[440] 
* INPUT : din0[441] 
* INPUT : din0[442] 
* INPUT : din0[443] 
* INPUT : din0[444] 
* INPUT : din0[445] 
* INPUT : din0[446] 
* INPUT : din0[447] 
* INPUT : din0[448] 
* INPUT : din0[449] 
* INPUT : din0[450] 
* INPUT : din0[451] 
* INPUT : din0[452] 
* INPUT : din0[453] 
* INPUT : din0[454] 
* INPUT : din0[455] 
* INPUT : din0[456] 
* INPUT : din0[457] 
* INPUT : din0[458] 
* INPUT : din0[459] 
* INPUT : din0[460] 
* INPUT : din0[461] 
* INPUT : din0[462] 
* INPUT : din0[463] 
* INPUT : din0[464] 
* INPUT : din0[465] 
* INPUT : din0[466] 
* INPUT : din0[467] 
* INPUT : din0[468] 
* INPUT : din0[469] 
* INPUT : din0[470] 
* INPUT : din0[471] 
* INPUT : din0[472] 
* INPUT : din0[473] 
* INPUT : din0[474] 
* INPUT : din0[475] 
* INPUT : din0[476] 
* INPUT : din0[477] 
* INPUT : din0[478] 
* INPUT : din0[479] 
* INPUT : din0[480] 
* INPUT : din0[481] 
* INPUT : din0[482] 
* INPUT : din0[483] 
* INPUT : din0[484] 
* INPUT : din0[485] 
* INPUT : din0[486] 
* INPUT : din0[487] 
* INPUT : din0[488] 
* INPUT : din0[489] 
* INPUT : din0[490] 
* INPUT : din0[491] 
* INPUT : din0[492] 
* INPUT : din0[493] 
* INPUT : din0[494] 
* INPUT : din0[495] 
* INPUT : din0[496] 
* INPUT : din0[497] 
* INPUT : din0[498] 
* INPUT : din0[499] 
* INPUT : din0[500] 
* INPUT : din0[501] 
* INPUT : din0[502] 
* INPUT : din0[503] 
* INPUT : din0[504] 
* INPUT : din0[505] 
* INPUT : din0[506] 
* INPUT : din0[507] 
* INPUT : din0[508] 
* INPUT : din0[509] 
* INPUT : din0[510] 
* INPUT : din0[511] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* OUTPUT: dout0[32] 
* OUTPUT: dout0[33] 
* OUTPUT: dout0[34] 
* OUTPUT: dout0[35] 
* OUTPUT: dout0[36] 
* OUTPUT: dout0[37] 
* OUTPUT: dout0[38] 
* OUTPUT: dout0[39] 
* OUTPUT: dout0[40] 
* OUTPUT: dout0[41] 
* OUTPUT: dout0[42] 
* OUTPUT: dout0[43] 
* OUTPUT: dout0[44] 
* OUTPUT: dout0[45] 
* OUTPUT: dout0[46] 
* OUTPUT: dout0[47] 
* OUTPUT: dout0[48] 
* OUTPUT: dout0[49] 
* OUTPUT: dout0[50] 
* OUTPUT: dout0[51] 
* OUTPUT: dout0[52] 
* OUTPUT: dout0[53] 
* OUTPUT: dout0[54] 
* OUTPUT: dout0[55] 
* OUTPUT: dout0[56] 
* OUTPUT: dout0[57] 
* OUTPUT: dout0[58] 
* OUTPUT: dout0[59] 
* OUTPUT: dout0[60] 
* OUTPUT: dout0[61] 
* OUTPUT: dout0[62] 
* OUTPUT: dout0[63] 
* OUTPUT: dout0[64] 
* OUTPUT: dout0[65] 
* OUTPUT: dout0[66] 
* OUTPUT: dout0[67] 
* OUTPUT: dout0[68] 
* OUTPUT: dout0[69] 
* OUTPUT: dout0[70] 
* OUTPUT: dout0[71] 
* OUTPUT: dout0[72] 
* OUTPUT: dout0[73] 
* OUTPUT: dout0[74] 
* OUTPUT: dout0[75] 
* OUTPUT: dout0[76] 
* OUTPUT: dout0[77] 
* OUTPUT: dout0[78] 
* OUTPUT: dout0[79] 
* OUTPUT: dout0[80] 
* OUTPUT: dout0[81] 
* OUTPUT: dout0[82] 
* OUTPUT: dout0[83] 
* OUTPUT: dout0[84] 
* OUTPUT: dout0[85] 
* OUTPUT: dout0[86] 
* OUTPUT: dout0[87] 
* OUTPUT: dout0[88] 
* OUTPUT: dout0[89] 
* OUTPUT: dout0[90] 
* OUTPUT: dout0[91] 
* OUTPUT: dout0[92] 
* OUTPUT: dout0[93] 
* OUTPUT: dout0[94] 
* OUTPUT: dout0[95] 
* OUTPUT: dout0[96] 
* OUTPUT: dout0[97] 
* OUTPUT: dout0[98] 
* OUTPUT: dout0[99] 
* OUTPUT: dout0[100] 
* OUTPUT: dout0[101] 
* OUTPUT: dout0[102] 
* OUTPUT: dout0[103] 
* OUTPUT: dout0[104] 
* OUTPUT: dout0[105] 
* OUTPUT: dout0[106] 
* OUTPUT: dout0[107] 
* OUTPUT: dout0[108] 
* OUTPUT: dout0[109] 
* OUTPUT: dout0[110] 
* OUTPUT: dout0[111] 
* OUTPUT: dout0[112] 
* OUTPUT: dout0[113] 
* OUTPUT: dout0[114] 
* OUTPUT: dout0[115] 
* OUTPUT: dout0[116] 
* OUTPUT: dout0[117] 
* OUTPUT: dout0[118] 
* OUTPUT: dout0[119] 
* OUTPUT: dout0[120] 
* OUTPUT: dout0[121] 
* OUTPUT: dout0[122] 
* OUTPUT: dout0[123] 
* OUTPUT: dout0[124] 
* OUTPUT: dout0[125] 
* OUTPUT: dout0[126] 
* OUTPUT: dout0[127] 
* OUTPUT: dout0[128] 
* OUTPUT: dout0[129] 
* OUTPUT: dout0[130] 
* OUTPUT: dout0[131] 
* OUTPUT: dout0[132] 
* OUTPUT: dout0[133] 
* OUTPUT: dout0[134] 
* OUTPUT: dout0[135] 
* OUTPUT: dout0[136] 
* OUTPUT: dout0[137] 
* OUTPUT: dout0[138] 
* OUTPUT: dout0[139] 
* OUTPUT: dout0[140] 
* OUTPUT: dout0[141] 
* OUTPUT: dout0[142] 
* OUTPUT: dout0[143] 
* OUTPUT: dout0[144] 
* OUTPUT: dout0[145] 
* OUTPUT: dout0[146] 
* OUTPUT: dout0[147] 
* OUTPUT: dout0[148] 
* OUTPUT: dout0[149] 
* OUTPUT: dout0[150] 
* OUTPUT: dout0[151] 
* OUTPUT: dout0[152] 
* OUTPUT: dout0[153] 
* OUTPUT: dout0[154] 
* OUTPUT: dout0[155] 
* OUTPUT: dout0[156] 
* OUTPUT: dout0[157] 
* OUTPUT: dout0[158] 
* OUTPUT: dout0[159] 
* OUTPUT: dout0[160] 
* OUTPUT: dout0[161] 
* OUTPUT: dout0[162] 
* OUTPUT: dout0[163] 
* OUTPUT: dout0[164] 
* OUTPUT: dout0[165] 
* OUTPUT: dout0[166] 
* OUTPUT: dout0[167] 
* OUTPUT: dout0[168] 
* OUTPUT: dout0[169] 
* OUTPUT: dout0[170] 
* OUTPUT: dout0[171] 
* OUTPUT: dout0[172] 
* OUTPUT: dout0[173] 
* OUTPUT: dout0[174] 
* OUTPUT: dout0[175] 
* OUTPUT: dout0[176] 
* OUTPUT: dout0[177] 
* OUTPUT: dout0[178] 
* OUTPUT: dout0[179] 
* OUTPUT: dout0[180] 
* OUTPUT: dout0[181] 
* OUTPUT: dout0[182] 
* OUTPUT: dout0[183] 
* OUTPUT: dout0[184] 
* OUTPUT: dout0[185] 
* OUTPUT: dout0[186] 
* OUTPUT: dout0[187] 
* OUTPUT: dout0[188] 
* OUTPUT: dout0[189] 
* OUTPUT: dout0[190] 
* OUTPUT: dout0[191] 
* OUTPUT: dout0[192] 
* OUTPUT: dout0[193] 
* OUTPUT: dout0[194] 
* OUTPUT: dout0[195] 
* OUTPUT: dout0[196] 
* OUTPUT: dout0[197] 
* OUTPUT: dout0[198] 
* OUTPUT: dout0[199] 
* OUTPUT: dout0[200] 
* OUTPUT: dout0[201] 
* OUTPUT: dout0[202] 
* OUTPUT: dout0[203] 
* OUTPUT: dout0[204] 
* OUTPUT: dout0[205] 
* OUTPUT: dout0[206] 
* OUTPUT: dout0[207] 
* OUTPUT: dout0[208] 
* OUTPUT: dout0[209] 
* OUTPUT: dout0[210] 
* OUTPUT: dout0[211] 
* OUTPUT: dout0[212] 
* OUTPUT: dout0[213] 
* OUTPUT: dout0[214] 
* OUTPUT: dout0[215] 
* OUTPUT: dout0[216] 
* OUTPUT: dout0[217] 
* OUTPUT: dout0[218] 
* OUTPUT: dout0[219] 
* OUTPUT: dout0[220] 
* OUTPUT: dout0[221] 
* OUTPUT: dout0[222] 
* OUTPUT: dout0[223] 
* OUTPUT: dout0[224] 
* OUTPUT: dout0[225] 
* OUTPUT: dout0[226] 
* OUTPUT: dout0[227] 
* OUTPUT: dout0[228] 
* OUTPUT: dout0[229] 
* OUTPUT: dout0[230] 
* OUTPUT: dout0[231] 
* OUTPUT: dout0[232] 
* OUTPUT: dout0[233] 
* OUTPUT: dout0[234] 
* OUTPUT: dout0[235] 
* OUTPUT: dout0[236] 
* OUTPUT: dout0[237] 
* OUTPUT: dout0[238] 
* OUTPUT: dout0[239] 
* OUTPUT: dout0[240] 
* OUTPUT: dout0[241] 
* OUTPUT: dout0[242] 
* OUTPUT: dout0[243] 
* OUTPUT: dout0[244] 
* OUTPUT: dout0[245] 
* OUTPUT: dout0[246] 
* OUTPUT: dout0[247] 
* OUTPUT: dout0[248] 
* OUTPUT: dout0[249] 
* OUTPUT: dout0[250] 
* OUTPUT: dout0[251] 
* OUTPUT: dout0[252] 
* OUTPUT: dout0[253] 
* OUTPUT: dout0[254] 
* OUTPUT: dout0[255] 
* OUTPUT: dout0[256] 
* OUTPUT: dout0[257] 
* OUTPUT: dout0[258] 
* OUTPUT: dout0[259] 
* OUTPUT: dout0[260] 
* OUTPUT: dout0[261] 
* OUTPUT: dout0[262] 
* OUTPUT: dout0[263] 
* OUTPUT: dout0[264] 
* OUTPUT: dout0[265] 
* OUTPUT: dout0[266] 
* OUTPUT: dout0[267] 
* OUTPUT: dout0[268] 
* OUTPUT: dout0[269] 
* OUTPUT: dout0[270] 
* OUTPUT: dout0[271] 
* OUTPUT: dout0[272] 
* OUTPUT: dout0[273] 
* OUTPUT: dout0[274] 
* OUTPUT: dout0[275] 
* OUTPUT: dout0[276] 
* OUTPUT: dout0[277] 
* OUTPUT: dout0[278] 
* OUTPUT: dout0[279] 
* OUTPUT: dout0[280] 
* OUTPUT: dout0[281] 
* OUTPUT: dout0[282] 
* OUTPUT: dout0[283] 
* OUTPUT: dout0[284] 
* OUTPUT: dout0[285] 
* OUTPUT: dout0[286] 
* OUTPUT: dout0[287] 
* OUTPUT: dout0[288] 
* OUTPUT: dout0[289] 
* OUTPUT: dout0[290] 
* OUTPUT: dout0[291] 
* OUTPUT: dout0[292] 
* OUTPUT: dout0[293] 
* OUTPUT: dout0[294] 
* OUTPUT: dout0[295] 
* OUTPUT: dout0[296] 
* OUTPUT: dout0[297] 
* OUTPUT: dout0[298] 
* OUTPUT: dout0[299] 
* OUTPUT: dout0[300] 
* OUTPUT: dout0[301] 
* OUTPUT: dout0[302] 
* OUTPUT: dout0[303] 
* OUTPUT: dout0[304] 
* OUTPUT: dout0[305] 
* OUTPUT: dout0[306] 
* OUTPUT: dout0[307] 
* OUTPUT: dout0[308] 
* OUTPUT: dout0[309] 
* OUTPUT: dout0[310] 
* OUTPUT: dout0[311] 
* OUTPUT: dout0[312] 
* OUTPUT: dout0[313] 
* OUTPUT: dout0[314] 
* OUTPUT: dout0[315] 
* OUTPUT: dout0[316] 
* OUTPUT: dout0[317] 
* OUTPUT: dout0[318] 
* OUTPUT: dout0[319] 
* OUTPUT: dout0[320] 
* OUTPUT: dout0[321] 
* OUTPUT: dout0[322] 
* OUTPUT: dout0[323] 
* OUTPUT: dout0[324] 
* OUTPUT: dout0[325] 
* OUTPUT: dout0[326] 
* OUTPUT: dout0[327] 
* OUTPUT: dout0[328] 
* OUTPUT: dout0[329] 
* OUTPUT: dout0[330] 
* OUTPUT: dout0[331] 
* OUTPUT: dout0[332] 
* OUTPUT: dout0[333] 
* OUTPUT: dout0[334] 
* OUTPUT: dout0[335] 
* OUTPUT: dout0[336] 
* OUTPUT: dout0[337] 
* OUTPUT: dout0[338] 
* OUTPUT: dout0[339] 
* OUTPUT: dout0[340] 
* OUTPUT: dout0[341] 
* OUTPUT: dout0[342] 
* OUTPUT: dout0[343] 
* OUTPUT: dout0[344] 
* OUTPUT: dout0[345] 
* OUTPUT: dout0[346] 
* OUTPUT: dout0[347] 
* OUTPUT: dout0[348] 
* OUTPUT: dout0[349] 
* OUTPUT: dout0[350] 
* OUTPUT: dout0[351] 
* OUTPUT: dout0[352] 
* OUTPUT: dout0[353] 
* OUTPUT: dout0[354] 
* OUTPUT: dout0[355] 
* OUTPUT: dout0[356] 
* OUTPUT: dout0[357] 
* OUTPUT: dout0[358] 
* OUTPUT: dout0[359] 
* OUTPUT: dout0[360] 
* OUTPUT: dout0[361] 
* OUTPUT: dout0[362] 
* OUTPUT: dout0[363] 
* OUTPUT: dout0[364] 
* OUTPUT: dout0[365] 
* OUTPUT: dout0[366] 
* OUTPUT: dout0[367] 
* OUTPUT: dout0[368] 
* OUTPUT: dout0[369] 
* OUTPUT: dout0[370] 
* OUTPUT: dout0[371] 
* OUTPUT: dout0[372] 
* OUTPUT: dout0[373] 
* OUTPUT: dout0[374] 
* OUTPUT: dout0[375] 
* OUTPUT: dout0[376] 
* OUTPUT: dout0[377] 
* OUTPUT: dout0[378] 
* OUTPUT: dout0[379] 
* OUTPUT: dout0[380] 
* OUTPUT: dout0[381] 
* OUTPUT: dout0[382] 
* OUTPUT: dout0[383] 
* OUTPUT: dout0[384] 
* OUTPUT: dout0[385] 
* OUTPUT: dout0[386] 
* OUTPUT: dout0[387] 
* OUTPUT: dout0[388] 
* OUTPUT: dout0[389] 
* OUTPUT: dout0[390] 
* OUTPUT: dout0[391] 
* OUTPUT: dout0[392] 
* OUTPUT: dout0[393] 
* OUTPUT: dout0[394] 
* OUTPUT: dout0[395] 
* OUTPUT: dout0[396] 
* OUTPUT: dout0[397] 
* OUTPUT: dout0[398] 
* OUTPUT: dout0[399] 
* OUTPUT: dout0[400] 
* OUTPUT: dout0[401] 
* OUTPUT: dout0[402] 
* OUTPUT: dout0[403] 
* OUTPUT: dout0[404] 
* OUTPUT: dout0[405] 
* OUTPUT: dout0[406] 
* OUTPUT: dout0[407] 
* OUTPUT: dout0[408] 
* OUTPUT: dout0[409] 
* OUTPUT: dout0[410] 
* OUTPUT: dout0[411] 
* OUTPUT: dout0[412] 
* OUTPUT: dout0[413] 
* OUTPUT: dout0[414] 
* OUTPUT: dout0[415] 
* OUTPUT: dout0[416] 
* OUTPUT: dout0[417] 
* OUTPUT: dout0[418] 
* OUTPUT: dout0[419] 
* OUTPUT: dout0[420] 
* OUTPUT: dout0[421] 
* OUTPUT: dout0[422] 
* OUTPUT: dout0[423] 
* OUTPUT: dout0[424] 
* OUTPUT: dout0[425] 
* OUTPUT: dout0[426] 
* OUTPUT: dout0[427] 
* OUTPUT: dout0[428] 
* OUTPUT: dout0[429] 
* OUTPUT: dout0[430] 
* OUTPUT: dout0[431] 
* OUTPUT: dout0[432] 
* OUTPUT: dout0[433] 
* OUTPUT: dout0[434] 
* OUTPUT: dout0[435] 
* OUTPUT: dout0[436] 
* OUTPUT: dout0[437] 
* OUTPUT: dout0[438] 
* OUTPUT: dout0[439] 
* OUTPUT: dout0[440] 
* OUTPUT: dout0[441] 
* OUTPUT: dout0[442] 
* OUTPUT: dout0[443] 
* OUTPUT: dout0[444] 
* OUTPUT: dout0[445] 
* OUTPUT: dout0[446] 
* OUTPUT: dout0[447] 
* OUTPUT: dout0[448] 
* OUTPUT: dout0[449] 
* OUTPUT: dout0[450] 
* OUTPUT: dout0[451] 
* OUTPUT: dout0[452] 
* OUTPUT: dout0[453] 
* OUTPUT: dout0[454] 
* OUTPUT: dout0[455] 
* OUTPUT: dout0[456] 
* OUTPUT: dout0[457] 
* OUTPUT: dout0[458] 
* OUTPUT: dout0[459] 
* OUTPUT: dout0[460] 
* OUTPUT: dout0[461] 
* OUTPUT: dout0[462] 
* OUTPUT: dout0[463] 
* OUTPUT: dout0[464] 
* OUTPUT: dout0[465] 
* OUTPUT: dout0[466] 
* OUTPUT: dout0[467] 
* OUTPUT: dout0[468] 
* OUTPUT: dout0[469] 
* OUTPUT: dout0[470] 
* OUTPUT: dout0[471] 
* OUTPUT: dout0[472] 
* OUTPUT: dout0[473] 
* OUTPUT: dout0[474] 
* OUTPUT: dout0[475] 
* OUTPUT: dout0[476] 
* OUTPUT: dout0[477] 
* OUTPUT: dout0[478] 
* OUTPUT: dout0[479] 
* OUTPUT: dout0[480] 
* OUTPUT: dout0[481] 
* OUTPUT: dout0[482] 
* OUTPUT: dout0[483] 
* OUTPUT: dout0[484] 
* OUTPUT: dout0[485] 
* OUTPUT: dout0[486] 
* OUTPUT: dout0[487] 
* OUTPUT: dout0[488] 
* OUTPUT: dout0[489] 
* OUTPUT: dout0[490] 
* OUTPUT: dout0[491] 
* OUTPUT: dout0[492] 
* OUTPUT: dout0[493] 
* OUTPUT: dout0[494] 
* OUTPUT: dout0[495] 
* OUTPUT: dout0[496] 
* OUTPUT: dout0[497] 
* OUTPUT: dout0[498] 
* OUTPUT: dout0[499] 
* OUTPUT: dout0[500] 
* OUTPUT: dout0[501] 
* OUTPUT: dout0[502] 
* OUTPUT: dout0[503] 
* OUTPUT: dout0[504] 
* OUTPUT: dout0[505] 
* OUTPUT: dout0[506] 
* OUTPUT: dout0[507] 
* OUTPUT: dout0[508] 
* OUTPUT: dout0[509] 
* OUTPUT: dout0[510] 
* OUTPUT: dout0[511] 
* POWER : vdd 
* GROUND: gnd 
Xbank0
+ dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6]
+ dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13]
+ dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20]
+ dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34]
+ dout0[35] dout0[36] dout0[37] dout0[38] dout0[39] dout0[40] dout0[41]
+ dout0[42] dout0[43] dout0[44] dout0[45] dout0[46] dout0[47] dout0[48]
+ dout0[49] dout0[50] dout0[51] dout0[52] dout0[53] dout0[54] dout0[55]
+ dout0[56] dout0[57] dout0[58] dout0[59] dout0[60] dout0[61] dout0[62]
+ dout0[63] dout0[64] dout0[65] dout0[66] dout0[67] dout0[68] dout0[69]
+ dout0[70] dout0[71] dout0[72] dout0[73] dout0[74] dout0[75] dout0[76]
+ dout0[77] dout0[78] dout0[79] dout0[80] dout0[81] dout0[82] dout0[83]
+ dout0[84] dout0[85] dout0[86] dout0[87] dout0[88] dout0[89] dout0[90]
+ dout0[91] dout0[92] dout0[93] dout0[94] dout0[95] dout0[96] dout0[97]
+ dout0[98] dout0[99] dout0[100] dout0[101] dout0[102] dout0[103]
+ dout0[104] dout0[105] dout0[106] dout0[107] dout0[108] dout0[109]
+ dout0[110] dout0[111] dout0[112] dout0[113] dout0[114] dout0[115]
+ dout0[116] dout0[117] dout0[118] dout0[119] dout0[120] dout0[121]
+ dout0[122] dout0[123] dout0[124] dout0[125] dout0[126] dout0[127]
+ dout0[128] dout0[129] dout0[130] dout0[131] dout0[132] dout0[133]
+ dout0[134] dout0[135] dout0[136] dout0[137] dout0[138] dout0[139]
+ dout0[140] dout0[141] dout0[142] dout0[143] dout0[144] dout0[145]
+ dout0[146] dout0[147] dout0[148] dout0[149] dout0[150] dout0[151]
+ dout0[152] dout0[153] dout0[154] dout0[155] dout0[156] dout0[157]
+ dout0[158] dout0[159] dout0[160] dout0[161] dout0[162] dout0[163]
+ dout0[164] dout0[165] dout0[166] dout0[167] dout0[168] dout0[169]
+ dout0[170] dout0[171] dout0[172] dout0[173] dout0[174] dout0[175]
+ dout0[176] dout0[177] dout0[178] dout0[179] dout0[180] dout0[181]
+ dout0[182] dout0[183] dout0[184] dout0[185] dout0[186] dout0[187]
+ dout0[188] dout0[189] dout0[190] dout0[191] dout0[192] dout0[193]
+ dout0[194] dout0[195] dout0[196] dout0[197] dout0[198] dout0[199]
+ dout0[200] dout0[201] dout0[202] dout0[203] dout0[204] dout0[205]
+ dout0[206] dout0[207] dout0[208] dout0[209] dout0[210] dout0[211]
+ dout0[212] dout0[213] dout0[214] dout0[215] dout0[216] dout0[217]
+ dout0[218] dout0[219] dout0[220] dout0[221] dout0[222] dout0[223]
+ dout0[224] dout0[225] dout0[226] dout0[227] dout0[228] dout0[229]
+ dout0[230] dout0[231] dout0[232] dout0[233] dout0[234] dout0[235]
+ dout0[236] dout0[237] dout0[238] dout0[239] dout0[240] dout0[241]
+ dout0[242] dout0[243] dout0[244] dout0[245] dout0[246] dout0[247]
+ dout0[248] dout0[249] dout0[250] dout0[251] dout0[252] dout0[253]
+ dout0[254] dout0[255] dout0[256] dout0[257] dout0[258] dout0[259]
+ dout0[260] dout0[261] dout0[262] dout0[263] dout0[264] dout0[265]
+ dout0[266] dout0[267] dout0[268] dout0[269] dout0[270] dout0[271]
+ dout0[272] dout0[273] dout0[274] dout0[275] dout0[276] dout0[277]
+ dout0[278] dout0[279] dout0[280] dout0[281] dout0[282] dout0[283]
+ dout0[284] dout0[285] dout0[286] dout0[287] dout0[288] dout0[289]
+ dout0[290] dout0[291] dout0[292] dout0[293] dout0[294] dout0[295]
+ dout0[296] dout0[297] dout0[298] dout0[299] dout0[300] dout0[301]
+ dout0[302] dout0[303] dout0[304] dout0[305] dout0[306] dout0[307]
+ dout0[308] dout0[309] dout0[310] dout0[311] dout0[312] dout0[313]
+ dout0[314] dout0[315] dout0[316] dout0[317] dout0[318] dout0[319]
+ dout0[320] dout0[321] dout0[322] dout0[323] dout0[324] dout0[325]
+ dout0[326] dout0[327] dout0[328] dout0[329] dout0[330] dout0[331]
+ dout0[332] dout0[333] dout0[334] dout0[335] dout0[336] dout0[337]
+ dout0[338] dout0[339] dout0[340] dout0[341] dout0[342] dout0[343]
+ dout0[344] dout0[345] dout0[346] dout0[347] dout0[348] dout0[349]
+ dout0[350] dout0[351] dout0[352] dout0[353] dout0[354] dout0[355]
+ dout0[356] dout0[357] dout0[358] dout0[359] dout0[360] dout0[361]
+ dout0[362] dout0[363] dout0[364] dout0[365] dout0[366] dout0[367]
+ dout0[368] dout0[369] dout0[370] dout0[371] dout0[372] dout0[373]
+ dout0[374] dout0[375] dout0[376] dout0[377] dout0[378] dout0[379]
+ dout0[380] dout0[381] dout0[382] dout0[383] dout0[384] dout0[385]
+ dout0[386] dout0[387] dout0[388] dout0[389] dout0[390] dout0[391]
+ dout0[392] dout0[393] dout0[394] dout0[395] dout0[396] dout0[397]
+ dout0[398] dout0[399] dout0[400] dout0[401] dout0[402] dout0[403]
+ dout0[404] dout0[405] dout0[406] dout0[407] dout0[408] dout0[409]
+ dout0[410] dout0[411] dout0[412] dout0[413] dout0[414] dout0[415]
+ dout0[416] dout0[417] dout0[418] dout0[419] dout0[420] dout0[421]
+ dout0[422] dout0[423] dout0[424] dout0[425] dout0[426] dout0[427]
+ dout0[428] dout0[429] dout0[430] dout0[431] dout0[432] dout0[433]
+ dout0[434] dout0[435] dout0[436] dout0[437] dout0[438] dout0[439]
+ dout0[440] dout0[441] dout0[442] dout0[443] dout0[444] dout0[445]
+ dout0[446] dout0[447] dout0[448] dout0[449] dout0[450] dout0[451]
+ dout0[452] dout0[453] dout0[454] dout0[455] dout0[456] dout0[457]
+ dout0[458] dout0[459] dout0[460] dout0[461] dout0[462] dout0[463]
+ dout0[464] dout0[465] dout0[466] dout0[467] dout0[468] dout0[469]
+ dout0[470] dout0[471] dout0[472] dout0[473] dout0[474] dout0[475]
+ dout0[476] dout0[477] dout0[478] dout0[479] dout0[480] dout0[481]
+ dout0[482] dout0[483] dout0[484] dout0[485] dout0[486] dout0[487]
+ dout0[488] dout0[489] dout0[490] dout0[491] dout0[492] dout0[493]
+ dout0[494] dout0[495] dout0[496] dout0[497] dout0[498] dout0[499]
+ dout0[500] dout0[501] dout0[502] dout0[503] dout0[504] dout0[505]
+ dout0[506] dout0[507] dout0[508] dout0[509] dout0[510] dout0[511]
+ rbl_bl0 bank_din0_0 bank_din0_1 bank_din0_2 bank_din0_3 bank_din0_4
+ bank_din0_5 bank_din0_6 bank_din0_7 bank_din0_8 bank_din0_9
+ bank_din0_10 bank_din0_11 bank_din0_12 bank_din0_13 bank_din0_14
+ bank_din0_15 bank_din0_16 bank_din0_17 bank_din0_18 bank_din0_19
+ bank_din0_20 bank_din0_21 bank_din0_22 bank_din0_23 bank_din0_24
+ bank_din0_25 bank_din0_26 bank_din0_27 bank_din0_28 bank_din0_29
+ bank_din0_30 bank_din0_31 bank_din0_32 bank_din0_33 bank_din0_34
+ bank_din0_35 bank_din0_36 bank_din0_37 bank_din0_38 bank_din0_39
+ bank_din0_40 bank_din0_41 bank_din0_42 bank_din0_43 bank_din0_44
+ bank_din0_45 bank_din0_46 bank_din0_47 bank_din0_48 bank_din0_49
+ bank_din0_50 bank_din0_51 bank_din0_52 bank_din0_53 bank_din0_54
+ bank_din0_55 bank_din0_56 bank_din0_57 bank_din0_58 bank_din0_59
+ bank_din0_60 bank_din0_61 bank_din0_62 bank_din0_63 bank_din0_64
+ bank_din0_65 bank_din0_66 bank_din0_67 bank_din0_68 bank_din0_69
+ bank_din0_70 bank_din0_71 bank_din0_72 bank_din0_73 bank_din0_74
+ bank_din0_75 bank_din0_76 bank_din0_77 bank_din0_78 bank_din0_79
+ bank_din0_80 bank_din0_81 bank_din0_82 bank_din0_83 bank_din0_84
+ bank_din0_85 bank_din0_86 bank_din0_87 bank_din0_88 bank_din0_89
+ bank_din0_90 bank_din0_91 bank_din0_92 bank_din0_93 bank_din0_94
+ bank_din0_95 bank_din0_96 bank_din0_97 bank_din0_98 bank_din0_99
+ bank_din0_100 bank_din0_101 bank_din0_102 bank_din0_103 bank_din0_104
+ bank_din0_105 bank_din0_106 bank_din0_107 bank_din0_108 bank_din0_109
+ bank_din0_110 bank_din0_111 bank_din0_112 bank_din0_113 bank_din0_114
+ bank_din0_115 bank_din0_116 bank_din0_117 bank_din0_118 bank_din0_119
+ bank_din0_120 bank_din0_121 bank_din0_122 bank_din0_123 bank_din0_124
+ bank_din0_125 bank_din0_126 bank_din0_127 bank_din0_128 bank_din0_129
+ bank_din0_130 bank_din0_131 bank_din0_132 bank_din0_133 bank_din0_134
+ bank_din0_135 bank_din0_136 bank_din0_137 bank_din0_138 bank_din0_139
+ bank_din0_140 bank_din0_141 bank_din0_142 bank_din0_143 bank_din0_144
+ bank_din0_145 bank_din0_146 bank_din0_147 bank_din0_148 bank_din0_149
+ bank_din0_150 bank_din0_151 bank_din0_152 bank_din0_153 bank_din0_154
+ bank_din0_155 bank_din0_156 bank_din0_157 bank_din0_158 bank_din0_159
+ bank_din0_160 bank_din0_161 bank_din0_162 bank_din0_163 bank_din0_164
+ bank_din0_165 bank_din0_166 bank_din0_167 bank_din0_168 bank_din0_169
+ bank_din0_170 bank_din0_171 bank_din0_172 bank_din0_173 bank_din0_174
+ bank_din0_175 bank_din0_176 bank_din0_177 bank_din0_178 bank_din0_179
+ bank_din0_180 bank_din0_181 bank_din0_182 bank_din0_183 bank_din0_184
+ bank_din0_185 bank_din0_186 bank_din0_187 bank_din0_188 bank_din0_189
+ bank_din0_190 bank_din0_191 bank_din0_192 bank_din0_193 bank_din0_194
+ bank_din0_195 bank_din0_196 bank_din0_197 bank_din0_198 bank_din0_199
+ bank_din0_200 bank_din0_201 bank_din0_202 bank_din0_203 bank_din0_204
+ bank_din0_205 bank_din0_206 bank_din0_207 bank_din0_208 bank_din0_209
+ bank_din0_210 bank_din0_211 bank_din0_212 bank_din0_213 bank_din0_214
+ bank_din0_215 bank_din0_216 bank_din0_217 bank_din0_218 bank_din0_219
+ bank_din0_220 bank_din0_221 bank_din0_222 bank_din0_223 bank_din0_224
+ bank_din0_225 bank_din0_226 bank_din0_227 bank_din0_228 bank_din0_229
+ bank_din0_230 bank_din0_231 bank_din0_232 bank_din0_233 bank_din0_234
+ bank_din0_235 bank_din0_236 bank_din0_237 bank_din0_238 bank_din0_239
+ bank_din0_240 bank_din0_241 bank_din0_242 bank_din0_243 bank_din0_244
+ bank_din0_245 bank_din0_246 bank_din0_247 bank_din0_248 bank_din0_249
+ bank_din0_250 bank_din0_251 bank_din0_252 bank_din0_253 bank_din0_254
+ bank_din0_255 bank_din0_256 bank_din0_257 bank_din0_258 bank_din0_259
+ bank_din0_260 bank_din0_261 bank_din0_262 bank_din0_263 bank_din0_264
+ bank_din0_265 bank_din0_266 bank_din0_267 bank_din0_268 bank_din0_269
+ bank_din0_270 bank_din0_271 bank_din0_272 bank_din0_273 bank_din0_274
+ bank_din0_275 bank_din0_276 bank_din0_277 bank_din0_278 bank_din0_279
+ bank_din0_280 bank_din0_281 bank_din0_282 bank_din0_283 bank_din0_284
+ bank_din0_285 bank_din0_286 bank_din0_287 bank_din0_288 bank_din0_289
+ bank_din0_290 bank_din0_291 bank_din0_292 bank_din0_293 bank_din0_294
+ bank_din0_295 bank_din0_296 bank_din0_297 bank_din0_298 bank_din0_299
+ bank_din0_300 bank_din0_301 bank_din0_302 bank_din0_303 bank_din0_304
+ bank_din0_305 bank_din0_306 bank_din0_307 bank_din0_308 bank_din0_309
+ bank_din0_310 bank_din0_311 bank_din0_312 bank_din0_313 bank_din0_314
+ bank_din0_315 bank_din0_316 bank_din0_317 bank_din0_318 bank_din0_319
+ bank_din0_320 bank_din0_321 bank_din0_322 bank_din0_323 bank_din0_324
+ bank_din0_325 bank_din0_326 bank_din0_327 bank_din0_328 bank_din0_329
+ bank_din0_330 bank_din0_331 bank_din0_332 bank_din0_333 bank_din0_334
+ bank_din0_335 bank_din0_336 bank_din0_337 bank_din0_338 bank_din0_339
+ bank_din0_340 bank_din0_341 bank_din0_342 bank_din0_343 bank_din0_344
+ bank_din0_345 bank_din0_346 bank_din0_347 bank_din0_348 bank_din0_349
+ bank_din0_350 bank_din0_351 bank_din0_352 bank_din0_353 bank_din0_354
+ bank_din0_355 bank_din0_356 bank_din0_357 bank_din0_358 bank_din0_359
+ bank_din0_360 bank_din0_361 bank_din0_362 bank_din0_363 bank_din0_364
+ bank_din0_365 bank_din0_366 bank_din0_367 bank_din0_368 bank_din0_369
+ bank_din0_370 bank_din0_371 bank_din0_372 bank_din0_373 bank_din0_374
+ bank_din0_375 bank_din0_376 bank_din0_377 bank_din0_378 bank_din0_379
+ bank_din0_380 bank_din0_381 bank_din0_382 bank_din0_383 bank_din0_384
+ bank_din0_385 bank_din0_386 bank_din0_387 bank_din0_388 bank_din0_389
+ bank_din0_390 bank_din0_391 bank_din0_392 bank_din0_393 bank_din0_394
+ bank_din0_395 bank_din0_396 bank_din0_397 bank_din0_398 bank_din0_399
+ bank_din0_400 bank_din0_401 bank_din0_402 bank_din0_403 bank_din0_404
+ bank_din0_405 bank_din0_406 bank_din0_407 bank_din0_408 bank_din0_409
+ bank_din0_410 bank_din0_411 bank_din0_412 bank_din0_413 bank_din0_414
+ bank_din0_415 bank_din0_416 bank_din0_417 bank_din0_418 bank_din0_419
+ bank_din0_420 bank_din0_421 bank_din0_422 bank_din0_423 bank_din0_424
+ bank_din0_425 bank_din0_426 bank_din0_427 bank_din0_428 bank_din0_429
+ bank_din0_430 bank_din0_431 bank_din0_432 bank_din0_433 bank_din0_434
+ bank_din0_435 bank_din0_436 bank_din0_437 bank_din0_438 bank_din0_439
+ bank_din0_440 bank_din0_441 bank_din0_442 bank_din0_443 bank_din0_444
+ bank_din0_445 bank_din0_446 bank_din0_447 bank_din0_448 bank_din0_449
+ bank_din0_450 bank_din0_451 bank_din0_452 bank_din0_453 bank_din0_454
+ bank_din0_455 bank_din0_456 bank_din0_457 bank_din0_458 bank_din0_459
+ bank_din0_460 bank_din0_461 bank_din0_462 bank_din0_463 bank_din0_464
+ bank_din0_465 bank_din0_466 bank_din0_467 bank_din0_468 bank_din0_469
+ bank_din0_470 bank_din0_471 bank_din0_472 bank_din0_473 bank_din0_474
+ bank_din0_475 bank_din0_476 bank_din0_477 bank_din0_478 bank_din0_479
+ bank_din0_480 bank_din0_481 bank_din0_482 bank_din0_483 bank_din0_484
+ bank_din0_485 bank_din0_486 bank_din0_487 bank_din0_488 bank_din0_489
+ bank_din0_490 bank_din0_491 bank_din0_492 bank_din0_493 bank_din0_494
+ bank_din0_495 bank_din0_496 bank_din0_497 bank_din0_498 bank_din0_499
+ bank_din0_500 bank_din0_501 bank_din0_502 bank_din0_503 bank_din0_504
+ bank_din0_505 bank_din0_506 bank_din0_507 bank_din0_508 bank_din0_509
+ bank_din0_510 bank_din0_511 a0_0 a0_1 a0_2 a0_3 a0_4 a0_5 s_en0
+ p_en_bar0 w_en0 wl_en0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_bank
Xcontrol0
+ csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_control_logic_rw
Xrow_address0
+ addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] a0_0 a0_1 a0_2
+ a0_3 a0_4 a0_5 clk_buf0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_row_addr_dff
Xdata_dff0
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22]
+ din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29]
+ din0[30] din0[31] din0[32] din0[33] din0[34] din0[35] din0[36]
+ din0[37] din0[38] din0[39] din0[40] din0[41] din0[42] din0[43]
+ din0[44] din0[45] din0[46] din0[47] din0[48] din0[49] din0[50]
+ din0[51] din0[52] din0[53] din0[54] din0[55] din0[56] din0[57]
+ din0[58] din0[59] din0[60] din0[61] din0[62] din0[63] din0[64]
+ din0[65] din0[66] din0[67] din0[68] din0[69] din0[70] din0[71]
+ din0[72] din0[73] din0[74] din0[75] din0[76] din0[77] din0[78]
+ din0[79] din0[80] din0[81] din0[82] din0[83] din0[84] din0[85]
+ din0[86] din0[87] din0[88] din0[89] din0[90] din0[91] din0[92]
+ din0[93] din0[94] din0[95] din0[96] din0[97] din0[98] din0[99]
+ din0[100] din0[101] din0[102] din0[103] din0[104] din0[105] din0[106]
+ din0[107] din0[108] din0[109] din0[110] din0[111] din0[112] din0[113]
+ din0[114] din0[115] din0[116] din0[117] din0[118] din0[119] din0[120]
+ din0[121] din0[122] din0[123] din0[124] din0[125] din0[126] din0[127]
+ din0[128] din0[129] din0[130] din0[131] din0[132] din0[133] din0[134]
+ din0[135] din0[136] din0[137] din0[138] din0[139] din0[140] din0[141]
+ din0[142] din0[143] din0[144] din0[145] din0[146] din0[147] din0[148]
+ din0[149] din0[150] din0[151] din0[152] din0[153] din0[154] din0[155]
+ din0[156] din0[157] din0[158] din0[159] din0[160] din0[161] din0[162]
+ din0[163] din0[164] din0[165] din0[166] din0[167] din0[168] din0[169]
+ din0[170] din0[171] din0[172] din0[173] din0[174] din0[175] din0[176]
+ din0[177] din0[178] din0[179] din0[180] din0[181] din0[182] din0[183]
+ din0[184] din0[185] din0[186] din0[187] din0[188] din0[189] din0[190]
+ din0[191] din0[192] din0[193] din0[194] din0[195] din0[196] din0[197]
+ din0[198] din0[199] din0[200] din0[201] din0[202] din0[203] din0[204]
+ din0[205] din0[206] din0[207] din0[208] din0[209] din0[210] din0[211]
+ din0[212] din0[213] din0[214] din0[215] din0[216] din0[217] din0[218]
+ din0[219] din0[220] din0[221] din0[222] din0[223] din0[224] din0[225]
+ din0[226] din0[227] din0[228] din0[229] din0[230] din0[231] din0[232]
+ din0[233] din0[234] din0[235] din0[236] din0[237] din0[238] din0[239]
+ din0[240] din0[241] din0[242] din0[243] din0[244] din0[245] din0[246]
+ din0[247] din0[248] din0[249] din0[250] din0[251] din0[252] din0[253]
+ din0[254] din0[255] din0[256] din0[257] din0[258] din0[259] din0[260]
+ din0[261] din0[262] din0[263] din0[264] din0[265] din0[266] din0[267]
+ din0[268] din0[269] din0[270] din0[271] din0[272] din0[273] din0[274]
+ din0[275] din0[276] din0[277] din0[278] din0[279] din0[280] din0[281]
+ din0[282] din0[283] din0[284] din0[285] din0[286] din0[287] din0[288]
+ din0[289] din0[290] din0[291] din0[292] din0[293] din0[294] din0[295]
+ din0[296] din0[297] din0[298] din0[299] din0[300] din0[301] din0[302]
+ din0[303] din0[304] din0[305] din0[306] din0[307] din0[308] din0[309]
+ din0[310] din0[311] din0[312] din0[313] din0[314] din0[315] din0[316]
+ din0[317] din0[318] din0[319] din0[320] din0[321] din0[322] din0[323]
+ din0[324] din0[325] din0[326] din0[327] din0[328] din0[329] din0[330]
+ din0[331] din0[332] din0[333] din0[334] din0[335] din0[336] din0[337]
+ din0[338] din0[339] din0[340] din0[341] din0[342] din0[343] din0[344]
+ din0[345] din0[346] din0[347] din0[348] din0[349] din0[350] din0[351]
+ din0[352] din0[353] din0[354] din0[355] din0[356] din0[357] din0[358]
+ din0[359] din0[360] din0[361] din0[362] din0[363] din0[364] din0[365]
+ din0[366] din0[367] din0[368] din0[369] din0[370] din0[371] din0[372]
+ din0[373] din0[374] din0[375] din0[376] din0[377] din0[378] din0[379]
+ din0[380] din0[381] din0[382] din0[383] din0[384] din0[385] din0[386]
+ din0[387] din0[388] din0[389] din0[390] din0[391] din0[392] din0[393]
+ din0[394] din0[395] din0[396] din0[397] din0[398] din0[399] din0[400]
+ din0[401] din0[402] din0[403] din0[404] din0[405] din0[406] din0[407]
+ din0[408] din0[409] din0[410] din0[411] din0[412] din0[413] din0[414]
+ din0[415] din0[416] din0[417] din0[418] din0[419] din0[420] din0[421]
+ din0[422] din0[423] din0[424] din0[425] din0[426] din0[427] din0[428]
+ din0[429] din0[430] din0[431] din0[432] din0[433] din0[434] din0[435]
+ din0[436] din0[437] din0[438] din0[439] din0[440] din0[441] din0[442]
+ din0[443] din0[444] din0[445] din0[446] din0[447] din0[448] din0[449]
+ din0[450] din0[451] din0[452] din0[453] din0[454] din0[455] din0[456]
+ din0[457] din0[458] din0[459] din0[460] din0[461] din0[462] din0[463]
+ din0[464] din0[465] din0[466] din0[467] din0[468] din0[469] din0[470]
+ din0[471] din0[472] din0[473] din0[474] din0[475] din0[476] din0[477]
+ din0[478] din0[479] din0[480] din0[481] din0[482] din0[483] din0[484]
+ din0[485] din0[486] din0[487] din0[488] din0[489] din0[490] din0[491]
+ din0[492] din0[493] din0[494] din0[495] din0[496] din0[497] din0[498]
+ din0[499] din0[500] din0[501] din0[502] din0[503] din0[504] din0[505]
+ din0[506] din0[507] din0[508] din0[509] din0[510] din0[511]
+ bank_din0_0 bank_din0_1 bank_din0_2 bank_din0_3 bank_din0_4
+ bank_din0_5 bank_din0_6 bank_din0_7 bank_din0_8 bank_din0_9
+ bank_din0_10 bank_din0_11 bank_din0_12 bank_din0_13 bank_din0_14
+ bank_din0_15 bank_din0_16 bank_din0_17 bank_din0_18 bank_din0_19
+ bank_din0_20 bank_din0_21 bank_din0_22 bank_din0_23 bank_din0_24
+ bank_din0_25 bank_din0_26 bank_din0_27 bank_din0_28 bank_din0_29
+ bank_din0_30 bank_din0_31 bank_din0_32 bank_din0_33 bank_din0_34
+ bank_din0_35 bank_din0_36 bank_din0_37 bank_din0_38 bank_din0_39
+ bank_din0_40 bank_din0_41 bank_din0_42 bank_din0_43 bank_din0_44
+ bank_din0_45 bank_din0_46 bank_din0_47 bank_din0_48 bank_din0_49
+ bank_din0_50 bank_din0_51 bank_din0_52 bank_din0_53 bank_din0_54
+ bank_din0_55 bank_din0_56 bank_din0_57 bank_din0_58 bank_din0_59
+ bank_din0_60 bank_din0_61 bank_din0_62 bank_din0_63 bank_din0_64
+ bank_din0_65 bank_din0_66 bank_din0_67 bank_din0_68 bank_din0_69
+ bank_din0_70 bank_din0_71 bank_din0_72 bank_din0_73 bank_din0_74
+ bank_din0_75 bank_din0_76 bank_din0_77 bank_din0_78 bank_din0_79
+ bank_din0_80 bank_din0_81 bank_din0_82 bank_din0_83 bank_din0_84
+ bank_din0_85 bank_din0_86 bank_din0_87 bank_din0_88 bank_din0_89
+ bank_din0_90 bank_din0_91 bank_din0_92 bank_din0_93 bank_din0_94
+ bank_din0_95 bank_din0_96 bank_din0_97 bank_din0_98 bank_din0_99
+ bank_din0_100 bank_din0_101 bank_din0_102 bank_din0_103 bank_din0_104
+ bank_din0_105 bank_din0_106 bank_din0_107 bank_din0_108 bank_din0_109
+ bank_din0_110 bank_din0_111 bank_din0_112 bank_din0_113 bank_din0_114
+ bank_din0_115 bank_din0_116 bank_din0_117 bank_din0_118 bank_din0_119
+ bank_din0_120 bank_din0_121 bank_din0_122 bank_din0_123 bank_din0_124
+ bank_din0_125 bank_din0_126 bank_din0_127 bank_din0_128 bank_din0_129
+ bank_din0_130 bank_din0_131 bank_din0_132 bank_din0_133 bank_din0_134
+ bank_din0_135 bank_din0_136 bank_din0_137 bank_din0_138 bank_din0_139
+ bank_din0_140 bank_din0_141 bank_din0_142 bank_din0_143 bank_din0_144
+ bank_din0_145 bank_din0_146 bank_din0_147 bank_din0_148 bank_din0_149
+ bank_din0_150 bank_din0_151 bank_din0_152 bank_din0_153 bank_din0_154
+ bank_din0_155 bank_din0_156 bank_din0_157 bank_din0_158 bank_din0_159
+ bank_din0_160 bank_din0_161 bank_din0_162 bank_din0_163 bank_din0_164
+ bank_din0_165 bank_din0_166 bank_din0_167 bank_din0_168 bank_din0_169
+ bank_din0_170 bank_din0_171 bank_din0_172 bank_din0_173 bank_din0_174
+ bank_din0_175 bank_din0_176 bank_din0_177 bank_din0_178 bank_din0_179
+ bank_din0_180 bank_din0_181 bank_din0_182 bank_din0_183 bank_din0_184
+ bank_din0_185 bank_din0_186 bank_din0_187 bank_din0_188 bank_din0_189
+ bank_din0_190 bank_din0_191 bank_din0_192 bank_din0_193 bank_din0_194
+ bank_din0_195 bank_din0_196 bank_din0_197 bank_din0_198 bank_din0_199
+ bank_din0_200 bank_din0_201 bank_din0_202 bank_din0_203 bank_din0_204
+ bank_din0_205 bank_din0_206 bank_din0_207 bank_din0_208 bank_din0_209
+ bank_din0_210 bank_din0_211 bank_din0_212 bank_din0_213 bank_din0_214
+ bank_din0_215 bank_din0_216 bank_din0_217 bank_din0_218 bank_din0_219
+ bank_din0_220 bank_din0_221 bank_din0_222 bank_din0_223 bank_din0_224
+ bank_din0_225 bank_din0_226 bank_din0_227 bank_din0_228 bank_din0_229
+ bank_din0_230 bank_din0_231 bank_din0_232 bank_din0_233 bank_din0_234
+ bank_din0_235 bank_din0_236 bank_din0_237 bank_din0_238 bank_din0_239
+ bank_din0_240 bank_din0_241 bank_din0_242 bank_din0_243 bank_din0_244
+ bank_din0_245 bank_din0_246 bank_din0_247 bank_din0_248 bank_din0_249
+ bank_din0_250 bank_din0_251 bank_din0_252 bank_din0_253 bank_din0_254
+ bank_din0_255 bank_din0_256 bank_din0_257 bank_din0_258 bank_din0_259
+ bank_din0_260 bank_din0_261 bank_din0_262 bank_din0_263 bank_din0_264
+ bank_din0_265 bank_din0_266 bank_din0_267 bank_din0_268 bank_din0_269
+ bank_din0_270 bank_din0_271 bank_din0_272 bank_din0_273 bank_din0_274
+ bank_din0_275 bank_din0_276 bank_din0_277 bank_din0_278 bank_din0_279
+ bank_din0_280 bank_din0_281 bank_din0_282 bank_din0_283 bank_din0_284
+ bank_din0_285 bank_din0_286 bank_din0_287 bank_din0_288 bank_din0_289
+ bank_din0_290 bank_din0_291 bank_din0_292 bank_din0_293 bank_din0_294
+ bank_din0_295 bank_din0_296 bank_din0_297 bank_din0_298 bank_din0_299
+ bank_din0_300 bank_din0_301 bank_din0_302 bank_din0_303 bank_din0_304
+ bank_din0_305 bank_din0_306 bank_din0_307 bank_din0_308 bank_din0_309
+ bank_din0_310 bank_din0_311 bank_din0_312 bank_din0_313 bank_din0_314
+ bank_din0_315 bank_din0_316 bank_din0_317 bank_din0_318 bank_din0_319
+ bank_din0_320 bank_din0_321 bank_din0_322 bank_din0_323 bank_din0_324
+ bank_din0_325 bank_din0_326 bank_din0_327 bank_din0_328 bank_din0_329
+ bank_din0_330 bank_din0_331 bank_din0_332 bank_din0_333 bank_din0_334
+ bank_din0_335 bank_din0_336 bank_din0_337 bank_din0_338 bank_din0_339
+ bank_din0_340 bank_din0_341 bank_din0_342 bank_din0_343 bank_din0_344
+ bank_din0_345 bank_din0_346 bank_din0_347 bank_din0_348 bank_din0_349
+ bank_din0_350 bank_din0_351 bank_din0_352 bank_din0_353 bank_din0_354
+ bank_din0_355 bank_din0_356 bank_din0_357 bank_din0_358 bank_din0_359
+ bank_din0_360 bank_din0_361 bank_din0_362 bank_din0_363 bank_din0_364
+ bank_din0_365 bank_din0_366 bank_din0_367 bank_din0_368 bank_din0_369
+ bank_din0_370 bank_din0_371 bank_din0_372 bank_din0_373 bank_din0_374
+ bank_din0_375 bank_din0_376 bank_din0_377 bank_din0_378 bank_din0_379
+ bank_din0_380 bank_din0_381 bank_din0_382 bank_din0_383 bank_din0_384
+ bank_din0_385 bank_din0_386 bank_din0_387 bank_din0_388 bank_din0_389
+ bank_din0_390 bank_din0_391 bank_din0_392 bank_din0_393 bank_din0_394
+ bank_din0_395 bank_din0_396 bank_din0_397 bank_din0_398 bank_din0_399
+ bank_din0_400 bank_din0_401 bank_din0_402 bank_din0_403 bank_din0_404
+ bank_din0_405 bank_din0_406 bank_din0_407 bank_din0_408 bank_din0_409
+ bank_din0_410 bank_din0_411 bank_din0_412 bank_din0_413 bank_din0_414
+ bank_din0_415 bank_din0_416 bank_din0_417 bank_din0_418 bank_din0_419
+ bank_din0_420 bank_din0_421 bank_din0_422 bank_din0_423 bank_din0_424
+ bank_din0_425 bank_din0_426 bank_din0_427 bank_din0_428 bank_din0_429
+ bank_din0_430 bank_din0_431 bank_din0_432 bank_din0_433 bank_din0_434
+ bank_din0_435 bank_din0_436 bank_din0_437 bank_din0_438 bank_din0_439
+ bank_din0_440 bank_din0_441 bank_din0_442 bank_din0_443 bank_din0_444
+ bank_din0_445 bank_din0_446 bank_din0_447 bank_din0_448 bank_din0_449
+ bank_din0_450 bank_din0_451 bank_din0_452 bank_din0_453 bank_din0_454
+ bank_din0_455 bank_din0_456 bank_din0_457 bank_din0_458 bank_din0_459
+ bank_din0_460 bank_din0_461 bank_din0_462 bank_din0_463 bank_din0_464
+ bank_din0_465 bank_din0_466 bank_din0_467 bank_din0_468 bank_din0_469
+ bank_din0_470 bank_din0_471 bank_din0_472 bank_din0_473 bank_din0_474
+ bank_din0_475 bank_din0_476 bank_din0_477 bank_din0_478 bank_din0_479
+ bank_din0_480 bank_din0_481 bank_din0_482 bank_din0_483 bank_din0_484
+ bank_din0_485 bank_din0_486 bank_din0_487 bank_din0_488 bank_din0_489
+ bank_din0_490 bank_din0_491 bank_din0_492 bank_din0_493 bank_din0_494
+ bank_din0_495 bank_din0_496 bank_din0_497 bank_din0_498 bank_din0_499
+ bank_din0_500 bank_din0_501 bank_din0_502 bank_din0_503 bank_din0_504
+ bank_din0_505 bank_din0_506 bank_din0_507 bank_din0_508 bank_din0_509
+ bank_din0_510 bank_din0_511 clk_buf0 vdd gnd
+ freepdk45_sram_1rw0r_45x512_data_dff
.ENDS freepdk45_sram_1rw0r_45x512
