../macros/freepdk45_sram_1rw0r_64x40_20/freepdk45_sram_1rw0r_64x40_20.lef