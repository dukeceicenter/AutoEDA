../macros/freepdk45_sram_1w1r_120x16/freepdk45_sram_1w1r_120x16.lef