VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_128x4_1
   CLASS BLOCK ;
   SIZE 91.325 BY 83.985 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.635 1.105 34.77 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 1.105 37.63 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.355 1.105 40.49 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.215 1.105 43.35 1.24 ;
      END
   END din0[3]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14.615 1.105 14.75 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.475 1.105 17.61 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.335 1.105 20.47 1.24 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  8.895 46.71 9.03 46.845 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  8.895 49.44 9.03 49.575 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  8.895 51.65 9.03 51.785 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  8.895 54.38 9.03 54.515 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.575 82.745 73.71 82.88 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.715 82.745 70.85 82.88 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.855 82.745 67.99 82.88 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.155 29.55 82.29 29.685 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.155 26.82 82.29 26.955 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.155 24.61 82.29 24.745 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.155 21.88 82.29 22.015 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 11.09 0.42 11.225 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.905 71.49 91.04 71.625 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 11.175 6.3825 11.31 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.8025 71.405 84.9375 71.54 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.195 1.105 23.33 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.055 1.105 26.19 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.915 1.105 29.05 1.24 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.775 1.105 31.91 1.24 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.6625 68.5175 26.7975 68.6525 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.0625 68.5175 36.1975 68.6525 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.4625 68.5175 45.5975 68.6525 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.8625 68.5175 54.9975 68.6525 ;
      END
   END dout1[3]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  76.4225 35.14 76.5575 35.275 ;
         LAYER metal3 ;
         RECT  76.4225 44.11 76.5575 44.245 ;
         LAYER metal3 ;
         RECT  68.5225 56.07 68.6575 56.205 ;
         LAYER metal3 ;
         RECT  23.3425 16.65 23.4775 16.785 ;
         LAYER metal3 ;
         RECT  14.4325 41.12 14.5675 41.255 ;
         LAYER metal4 ;
         RECT  67.44 27.4825 67.58 57.6325 ;
         LAYER metal3 ;
         RECT  2.425 12.455 2.56 12.59 ;
         LAYER metal4 ;
         RECT  8.61 45.6025 8.75 55.6225 ;
         LAYER metal3 ;
         RECT  14.4325 44.11 14.5675 44.245 ;
         LAYER metal4 ;
         RECT  22.33 30.6525 22.47 54.7125 ;
         LAYER metal3 ;
         RECT  76.4225 32.15 76.5575 32.285 ;
         LAYER metal3 ;
         RECT  64.2275 16.65 64.3625 16.785 ;
         LAYER metal3 ;
         RECT  88.765 70.125 88.9 70.26 ;
         LAYER metal3 ;
         RECT  76.4225 41.12 76.5575 41.255 ;
         LAYER metal4 ;
         RECT  23.41 27.4825 23.55 57.6325 ;
         LAYER metal3 ;
         RECT  14.3325 2.47 14.4675 2.605 ;
         LAYER metal4 ;
         RECT  11.33 12.4525 11.47 27.4125 ;
         LAYER metal4 ;
         RECT  68.52 30.6525 68.66 54.7125 ;
         LAYER metal4 ;
         RECT  79.715 60.2425 79.855 70.2625 ;
         LAYER metal3 ;
         RECT  22.9125 2.47 23.0475 2.605 ;
         LAYER metal4 ;
         RECT  74.39 60.72 74.53 80.62 ;
         LAYER metal3 ;
         RECT  23.4775 65.96 55.6675 66.03 ;
         LAYER metal3 ;
         RECT  23.4775 26.7875 64.3625 26.8575 ;
         LAYER metal3 ;
         RECT  22.3325 29.16 22.4675 29.295 ;
         LAYER metal4 ;
         RECT  82.435 20.7725 82.575 30.7925 ;
         LAYER metal3 ;
         RECT  34.3525 2.47 34.4875 2.605 ;
         LAYER metal4 ;
         RECT  19.08 30.6525 19.22 54.7825 ;
         LAYER metal4 ;
         RECT  16.46 4.565 16.6 24.465 ;
         LAYER metal3 ;
         RECT  71.155 55.2825 71.29 55.4175 ;
         LAYER metal3 ;
         RECT  14.4325 35.14 14.5675 35.275 ;
         LAYER metal3 ;
         RECT  19.7 29.9475 19.835 30.0825 ;
         LAYER metal3 ;
         RECT  14.4325 32.15 14.5675 32.285 ;
         LAYER metal4 ;
         RECT  90.4975 40.4825 90.6375 62.885 ;
         LAYER metal4 ;
         RECT  0.6875 19.83 0.8275 42.2325 ;
         LAYER metal4 ;
         RECT  71.77 30.6525 71.91 54.7825 ;
         LAYER metal3 ;
         RECT  23.4775 17.6175 55.6675 17.6875 ;
         LAYER metal3 ;
         RECT  73.8575 81.38 73.9925 81.515 ;
         LAYER metal3 ;
         RECT  23.4775 58.3275 65.5375 58.3975 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  23.4775 64.0675 55.7025 64.1375 ;
         LAYER metal3 ;
         RECT  12.905 36.635 13.04 36.77 ;
         LAYER metal4 ;
         RECT  76.3325 60.6525 76.4725 80.6875 ;
         LAYER metal3 ;
         RECT  77.95 42.615 78.085 42.75 ;
         LAYER metal4 ;
         RECT  6.105 9.9825 6.245 24.9425 ;
         LAYER metal4 ;
         RECT  11.47 45.5375 11.61 55.6875 ;
         LAYER metal3 ;
         RECT  37.2125 0.0 37.3475 0.135 ;
         LAYER metal3 ;
         RECT  77.95 36.635 78.085 36.77 ;
         LAYER metal4 ;
         RECT  73.36 30.62 73.5 54.7825 ;
         LAYER metal4 ;
         RECT  23.87 27.4825 24.01 57.6325 ;
         LAYER metal4 ;
         RECT  71.21 30.62 71.35 54.745 ;
         LAYER metal3 ;
         RECT  12.905 30.655 13.04 30.79 ;
         LAYER metal3 ;
         RECT  77.95 39.625 78.085 39.76 ;
         LAYER metal3 ;
         RECT  64.2275 14.83 64.3625 14.965 ;
         LAYER metal3 ;
         RECT  12.905 33.645 13.04 33.78 ;
         LAYER metal3 ;
         RECT  77.95 30.655 78.085 30.79 ;
         LAYER metal4 ;
         RECT  2.75 19.8625 2.89 42.265 ;
         LAYER metal3 ;
         RECT  25.7725 0.0 25.9075 0.135 ;
         LAYER metal3 ;
         RECT  23.4775 60.9475 64.395 61.0175 ;
         LAYER metal4 ;
         RECT  66.98 27.4825 67.12 57.6325 ;
         LAYER metal3 ;
         RECT  23.4775 19.6675 55.6675 19.7375 ;
         LAYER metal3 ;
         RECT  88.765 72.595 88.9 72.73 ;
         LAYER metal3 ;
         RECT  77.95 33.645 78.085 33.78 ;
         LAYER metal3 ;
         RECT  23.3425 14.83 23.4775 14.965 ;
         LAYER metal3 ;
         RECT  23.4775 24.1675 64.395 24.2375 ;
         LAYER metal4 ;
         RECT  19.64 30.62 19.78 54.745 ;
         LAYER metal3 ;
         RECT  2.425 9.985 2.56 10.12 ;
         LAYER metal3 ;
         RECT  70.9975 83.85 71.1325 83.985 ;
         LAYER metal4 ;
         RECT  17.49 30.62 17.63 54.7825 ;
         LAYER metal3 ;
         RECT  12.905 39.625 13.04 39.76 ;
         LAYER metal3 ;
         RECT  77.95 45.605 78.085 45.74 ;
         LAYER metal4 ;
         RECT  88.435 40.45 88.575 62.8525 ;
         LAYER metal4 ;
         RECT  84.94 57.7725 85.08 72.7325 ;
         LAYER metal3 ;
         RECT  12.905 42.615 13.04 42.75 ;
         LAYER metal3 ;
         RECT  17.1925 0.0 17.3275 0.135 ;
         LAYER metal3 ;
         RECT  12.905 45.605 13.04 45.74 ;
         LAYER metal4 ;
         RECT  14.5175 4.4975 14.6575 24.5325 ;
         LAYER metal4 ;
         RECT  79.575 20.7075 79.715 30.8575 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 91.185 83.845 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 91.185 83.845 ;
   LAYER  metal3 ;
      RECT  34.495 0.14 34.91 0.965 ;
      RECT  34.91 0.965 37.355 1.38 ;
      RECT  37.77 0.965 40.215 1.38 ;
      RECT  40.63 0.965 43.075 1.38 ;
      RECT  43.49 0.965 91.185 1.38 ;
      RECT  0.14 0.965 14.475 1.38 ;
      RECT  14.89 0.965 17.335 1.38 ;
      RECT  17.75 0.965 20.195 1.38 ;
      RECT  0.14 46.57 8.755 46.985 ;
      RECT  0.14 46.985 8.755 83.845 ;
      RECT  8.755 1.38 9.17 46.57 ;
      RECT  9.17 46.57 34.495 46.985 ;
      RECT  8.755 46.985 9.17 49.3 ;
      RECT  8.755 49.715 9.17 51.51 ;
      RECT  8.755 51.925 9.17 54.24 ;
      RECT  8.755 54.655 9.17 83.845 ;
      RECT  73.435 83.02 73.85 83.845 ;
      RECT  73.85 82.605 91.185 83.02 ;
      RECT  73.85 83.02 91.185 83.845 ;
      RECT  70.99 82.605 73.435 83.02 ;
      RECT  34.91 82.605 67.715 83.02 ;
      RECT  68.13 82.605 70.575 83.02 ;
      RECT  73.85 1.38 82.015 29.41 ;
      RECT  73.85 29.41 82.015 29.825 ;
      RECT  82.015 29.825 82.43 82.605 ;
      RECT  82.43 1.38 91.185 29.41 ;
      RECT  82.43 29.41 91.185 29.825 ;
      RECT  82.015 27.095 82.43 29.41 ;
      RECT  82.015 24.885 82.43 26.68 ;
      RECT  82.015 1.38 82.43 21.74 ;
      RECT  82.015 22.155 82.43 24.47 ;
      RECT  0.14 1.38 0.145 10.95 ;
      RECT  0.14 10.95 0.145 11.365 ;
      RECT  0.14 11.365 0.145 46.57 ;
      RECT  0.145 1.38 0.56 10.95 ;
      RECT  0.145 11.365 0.56 46.57 ;
      RECT  90.765 29.825 91.18 71.35 ;
      RECT  90.765 71.765 91.18 82.605 ;
      RECT  91.18 29.825 91.185 71.35 ;
      RECT  91.18 71.35 91.185 71.765 ;
      RECT  91.18 71.765 91.185 82.605 ;
      RECT  0.56 10.95 6.1075 11.035 ;
      RECT  0.56 11.035 6.1075 11.365 ;
      RECT  6.1075 10.95 6.5225 11.035 ;
      RECT  6.5225 10.95 8.755 11.035 ;
      RECT  6.5225 11.035 8.755 11.365 ;
      RECT  0.56 11.365 6.1075 11.45 ;
      RECT  6.1075 11.45 6.5225 46.57 ;
      RECT  6.5225 11.365 8.755 11.45 ;
      RECT  6.5225 11.45 8.755 46.57 ;
      RECT  82.43 29.825 84.6625 71.265 ;
      RECT  82.43 71.265 84.6625 71.35 ;
      RECT  84.6625 29.825 85.0775 71.265 ;
      RECT  85.0775 71.265 90.765 71.35 ;
      RECT  82.43 71.35 84.6625 71.68 ;
      RECT  82.43 71.68 84.6625 71.765 ;
      RECT  84.6625 71.68 85.0775 71.765 ;
      RECT  85.0775 71.35 90.765 71.68 ;
      RECT  85.0775 71.68 90.765 71.765 ;
      RECT  20.61 0.965 23.055 1.38 ;
      RECT  23.47 0.965 25.915 1.38 ;
      RECT  26.33 0.965 28.775 1.38 ;
      RECT  29.19 0.965 31.635 1.38 ;
      RECT  32.05 0.965 34.495 1.38 ;
      RECT  9.17 68.3775 26.5225 68.7925 ;
      RECT  9.17 68.7925 26.5225 83.845 ;
      RECT  26.5225 68.7925 26.9375 83.845 ;
      RECT  26.9375 68.3775 34.495 68.7925 ;
      RECT  26.9375 68.7925 34.495 83.845 ;
      RECT  34.91 68.3775 35.9225 68.7925 ;
      RECT  34.91 68.7925 35.9225 82.605 ;
      RECT  35.9225 68.7925 36.3375 82.605 ;
      RECT  36.3375 68.7925 73.435 82.605 ;
      RECT  36.3375 68.3775 45.3225 68.7925 ;
      RECT  45.7375 68.3775 54.7225 68.7925 ;
      RECT  55.1375 68.3775 73.435 68.7925 ;
      RECT  73.85 29.825 76.2825 35.0 ;
      RECT  73.85 35.0 76.2825 35.415 ;
      RECT  76.6975 35.0 82.015 35.415 ;
      RECT  76.2825 44.385 76.6975 82.605 ;
      RECT  36.3375 55.93 68.3825 56.345 ;
      RECT  68.3825 1.38 68.7975 55.93 ;
      RECT  68.3825 56.345 68.7975 68.3775 ;
      RECT  68.7975 55.93 73.435 56.345 ;
      RECT  68.7975 56.345 73.435 68.3775 ;
      RECT  9.17 16.51 23.2025 16.925 ;
      RECT  23.6175 16.51 34.495 16.925 ;
      RECT  9.17 40.98 14.2925 41.395 ;
      RECT  14.7075 40.98 23.2025 41.395 ;
      RECT  14.7075 41.395 23.2025 46.57 ;
      RECT  0.56 11.45 2.285 12.315 ;
      RECT  0.56 12.315 2.285 12.73 ;
      RECT  0.56 12.73 2.285 46.57 ;
      RECT  2.285 11.45 2.7 12.315 ;
      RECT  2.285 12.73 2.7 46.57 ;
      RECT  2.7 11.45 6.1075 12.315 ;
      RECT  2.7 12.315 6.1075 12.73 ;
      RECT  2.7 12.73 6.1075 46.57 ;
      RECT  14.2925 41.395 14.7075 43.97 ;
      RECT  14.2925 44.385 14.7075 46.57 ;
      RECT  76.2825 29.825 76.6975 32.01 ;
      RECT  76.2825 32.425 76.6975 35.0 ;
      RECT  36.3375 1.38 64.0875 16.51 ;
      RECT  36.3375 16.51 64.0875 16.925 ;
      RECT  64.5025 1.38 68.3825 16.51 ;
      RECT  64.5025 16.51 68.3825 16.925 ;
      RECT  85.0775 29.825 88.625 69.985 ;
      RECT  85.0775 69.985 88.625 70.4 ;
      RECT  85.0775 70.4 88.625 71.265 ;
      RECT  88.625 29.825 89.04 69.985 ;
      RECT  88.625 70.4 89.04 71.265 ;
      RECT  89.04 29.825 90.765 69.985 ;
      RECT  89.04 69.985 90.765 70.4 ;
      RECT  89.04 70.4 90.765 71.265 ;
      RECT  76.2825 35.415 76.6975 40.98 ;
      RECT  76.2825 41.395 76.6975 43.97 ;
      RECT  9.17 1.38 14.1925 2.33 ;
      RECT  9.17 2.33 14.1925 2.745 ;
      RECT  9.17 2.745 14.1925 16.51 ;
      RECT  14.1925 1.38 14.6075 2.33 ;
      RECT  14.1925 2.745 14.6075 16.51 ;
      RECT  14.6075 1.38 23.2025 2.33 ;
      RECT  14.6075 2.745 23.2025 16.51 ;
      RECT  14.6075 2.33 22.7725 2.745 ;
      RECT  23.1875 2.33 23.2025 2.745 ;
      RECT  34.495 66.17 34.91 83.845 ;
      RECT  9.17 46.985 23.3375 65.82 ;
      RECT  9.17 65.82 23.3375 66.17 ;
      RECT  9.17 66.17 23.3375 68.3775 ;
      RECT  23.3375 66.17 26.5225 68.3775 ;
      RECT  26.5225 66.17 26.9375 68.3775 ;
      RECT  26.9375 66.17 34.495 68.3775 ;
      RECT  34.91 66.17 35.9225 68.3775 ;
      RECT  35.9225 66.17 36.3375 68.3775 ;
      RECT  36.3375 66.17 55.8075 68.3775 ;
      RECT  55.8075 65.82 68.3825 66.17 ;
      RECT  55.8075 66.17 68.3825 68.3775 ;
      RECT  23.2025 16.925 23.3375 26.6475 ;
      RECT  23.2025 26.6475 23.3375 26.9975 ;
      RECT  23.2025 26.9975 23.3375 46.57 ;
      RECT  23.3375 26.9975 23.6175 46.57 ;
      RECT  23.6175 26.9975 34.495 46.57 ;
      RECT  36.3375 26.9975 64.0875 55.93 ;
      RECT  64.0875 26.9975 64.5025 55.93 ;
      RECT  14.7075 16.925 22.1925 29.02 ;
      RECT  14.7075 29.02 22.1925 29.435 ;
      RECT  22.1925 16.925 22.6075 29.02 ;
      RECT  22.1925 29.435 22.6075 40.98 ;
      RECT  22.6075 16.925 23.2025 29.02 ;
      RECT  22.6075 29.02 23.2025 29.435 ;
      RECT  22.6075 29.435 23.2025 40.98 ;
      RECT  23.6175 1.38 34.2125 2.33 ;
      RECT  23.6175 2.33 34.2125 2.745 ;
      RECT  23.6175 2.745 34.2125 16.51 ;
      RECT  34.2125 1.38 34.495 2.33 ;
      RECT  34.2125 2.745 34.495 16.51 ;
      RECT  34.495 1.38 34.6275 2.33 ;
      RECT  34.6275 1.38 34.91 2.33 ;
      RECT  34.6275 2.33 34.91 2.745 ;
      RECT  68.7975 1.38 71.015 55.1425 ;
      RECT  68.7975 55.1425 71.015 55.5575 ;
      RECT  68.7975 55.5575 71.015 55.93 ;
      RECT  71.015 1.38 71.43 55.1425 ;
      RECT  71.015 55.5575 71.43 55.93 ;
      RECT  71.43 1.38 73.435 55.1425 ;
      RECT  71.43 55.1425 73.435 55.5575 ;
      RECT  71.43 55.5575 73.435 55.93 ;
      RECT  14.2925 35.415 14.7075 40.98 ;
      RECT  14.7075 29.435 19.56 29.8075 ;
      RECT  14.7075 29.8075 19.56 30.2225 ;
      RECT  14.7075 30.2225 19.56 40.98 ;
      RECT  19.56 29.435 19.975 29.8075 ;
      RECT  19.56 30.2225 19.975 40.98 ;
      RECT  19.975 29.435 22.1925 29.8075 ;
      RECT  19.975 29.8075 22.1925 30.2225 ;
      RECT  19.975 30.2225 22.1925 40.98 ;
      RECT  14.2925 16.925 14.7075 32.01 ;
      RECT  14.2925 32.425 14.7075 35.0 ;
      RECT  23.3375 16.925 23.6175 17.4775 ;
      RECT  23.6175 16.925 34.495 17.4775 ;
      RECT  36.3375 16.925 55.8075 17.4775 ;
      RECT  55.8075 16.925 64.0875 17.4775 ;
      RECT  55.8075 17.4775 64.0875 17.8275 ;
      RECT  34.91 1.38 35.9225 17.4775 ;
      RECT  35.9225 1.38 36.3375 17.4775 ;
      RECT  34.495 2.745 34.6275 17.4775 ;
      RECT  34.6275 2.745 34.91 17.4775 ;
      RECT  73.435 1.38 73.7175 81.24 ;
      RECT  73.435 81.24 73.7175 81.655 ;
      RECT  73.435 81.655 73.7175 82.605 ;
      RECT  73.7175 1.38 73.85 81.24 ;
      RECT  73.7175 81.655 73.85 82.605 ;
      RECT  73.85 35.415 74.1325 81.24 ;
      RECT  73.85 81.655 74.1325 82.605 ;
      RECT  74.1325 35.415 76.2825 81.24 ;
      RECT  74.1325 81.24 76.2825 81.655 ;
      RECT  74.1325 81.655 76.2825 82.605 ;
      RECT  23.3375 46.985 26.5225 58.1875 ;
      RECT  26.5225 46.985 26.9375 58.1875 ;
      RECT  26.9375 46.985 34.495 58.1875 ;
      RECT  36.3375 56.345 55.8075 58.1875 ;
      RECT  55.8075 56.345 65.6775 58.1875 ;
      RECT  65.6775 56.345 68.3825 58.1875 ;
      RECT  65.6775 58.1875 68.3825 58.5375 ;
      RECT  65.6775 58.5375 68.3825 65.82 ;
      RECT  34.495 26.9975 34.91 58.1875 ;
      RECT  34.91 26.9975 35.9225 58.1875 ;
      RECT  35.9225 26.9975 36.3375 58.1875 ;
      RECT  23.3375 64.2775 26.5225 65.82 ;
      RECT  26.5225 64.2775 26.9375 65.82 ;
      RECT  26.9375 64.2775 34.495 65.82 ;
      RECT  36.3375 64.2775 55.8075 65.82 ;
      RECT  55.8075 64.2775 55.8425 65.82 ;
      RECT  55.8425 63.9275 65.6775 64.2775 ;
      RECT  55.8425 64.2775 65.6775 65.82 ;
      RECT  34.495 64.2775 34.91 65.82 ;
      RECT  34.91 64.2775 35.9225 65.82 ;
      RECT  35.9225 64.2775 36.3375 65.82 ;
      RECT  9.17 16.925 12.765 36.495 ;
      RECT  9.17 36.495 12.765 36.91 ;
      RECT  9.17 36.91 12.765 40.98 ;
      RECT  13.18 16.925 14.2925 36.495 ;
      RECT  13.18 36.495 14.2925 36.91 ;
      RECT  13.18 36.91 14.2925 40.98 ;
      RECT  76.6975 35.415 77.81 42.475 ;
      RECT  76.6975 42.475 77.81 42.89 ;
      RECT  76.6975 42.89 77.81 82.605 ;
      RECT  78.225 35.415 82.015 42.475 ;
      RECT  78.225 42.475 82.015 42.89 ;
      RECT  78.225 42.89 82.015 82.605 ;
      RECT  34.91 0.14 37.0725 0.275 ;
      RECT  34.91 0.275 37.0725 0.965 ;
      RECT  37.0725 0.275 37.4875 0.965 ;
      RECT  37.4875 0.14 91.185 0.275 ;
      RECT  37.4875 0.275 91.185 0.965 ;
      RECT  77.81 35.415 78.225 36.495 ;
      RECT  12.765 16.925 13.18 30.515 ;
      RECT  77.81 36.91 78.225 39.485 ;
      RECT  77.81 39.9 78.225 42.475 ;
      RECT  64.0875 1.38 64.5025 14.69 ;
      RECT  64.0875 15.105 64.5025 16.51 ;
      RECT  12.765 30.93 13.18 33.505 ;
      RECT  12.765 33.92 13.18 36.495 ;
      RECT  76.6975 29.825 77.81 30.515 ;
      RECT  76.6975 30.515 77.81 30.93 ;
      RECT  76.6975 30.93 77.81 35.0 ;
      RECT  77.81 29.825 78.225 30.515 ;
      RECT  78.225 29.825 82.015 30.515 ;
      RECT  78.225 30.515 82.015 30.93 ;
      RECT  78.225 30.93 82.015 35.0 ;
      RECT  0.14 0.275 25.6325 0.965 ;
      RECT  25.6325 0.275 26.0475 0.965 ;
      RECT  26.0475 0.14 34.495 0.275 ;
      RECT  26.0475 0.275 34.495 0.965 ;
      RECT  23.3375 58.5375 26.5225 60.8075 ;
      RECT  23.3375 61.1575 26.5225 63.9275 ;
      RECT  26.5225 58.5375 26.9375 60.8075 ;
      RECT  26.5225 61.1575 26.9375 63.9275 ;
      RECT  26.9375 58.5375 34.495 60.8075 ;
      RECT  26.9375 61.1575 34.495 63.9275 ;
      RECT  36.3375 58.5375 55.8075 60.8075 ;
      RECT  36.3375 61.1575 55.8075 63.9275 ;
      RECT  55.8075 58.5375 55.8425 60.8075 ;
      RECT  55.8075 61.1575 55.8425 63.9275 ;
      RECT  55.8425 58.5375 64.535 60.8075 ;
      RECT  55.8425 61.1575 64.535 63.9275 ;
      RECT  64.535 58.5375 65.6775 60.8075 ;
      RECT  64.535 60.8075 65.6775 61.1575 ;
      RECT  64.535 61.1575 65.6775 63.9275 ;
      RECT  34.495 58.5375 34.91 60.8075 ;
      RECT  34.495 61.1575 34.91 63.9275 ;
      RECT  34.91 58.5375 35.9225 60.8075 ;
      RECT  34.91 61.1575 35.9225 63.9275 ;
      RECT  35.9225 58.5375 36.3375 60.8075 ;
      RECT  35.9225 61.1575 36.3375 63.9275 ;
      RECT  23.3375 17.8275 23.6175 19.5275 ;
      RECT  23.6175 17.8275 34.495 19.5275 ;
      RECT  36.3375 17.8275 55.8075 19.5275 ;
      RECT  34.91 17.8275 35.9225 19.5275 ;
      RECT  35.9225 17.8275 36.3375 19.5275 ;
      RECT  34.495 17.8275 34.6275 19.5275 ;
      RECT  34.6275 17.8275 34.91 19.5275 ;
      RECT  82.43 71.765 88.625 72.455 ;
      RECT  82.43 72.455 88.625 72.87 ;
      RECT  82.43 72.87 88.625 82.605 ;
      RECT  88.625 71.765 89.04 72.455 ;
      RECT  88.625 72.87 89.04 82.605 ;
      RECT  89.04 71.765 90.765 72.455 ;
      RECT  89.04 72.455 90.765 72.87 ;
      RECT  89.04 72.87 90.765 82.605 ;
      RECT  77.81 30.93 78.225 33.505 ;
      RECT  77.81 33.92 78.225 35.0 ;
      RECT  23.2025 1.38 23.6175 14.69 ;
      RECT  23.2025 15.105 23.6175 16.51 ;
      RECT  64.5025 16.925 64.535 24.0275 ;
      RECT  64.5025 24.3775 64.535 55.93 ;
      RECT  64.535 16.925 68.3825 24.0275 ;
      RECT  64.535 24.0275 68.3825 24.3775 ;
      RECT  64.535 24.3775 68.3825 55.93 ;
      RECT  64.0875 16.925 64.5025 24.0275 ;
      RECT  64.0875 24.3775 64.5025 26.6475 ;
      RECT  55.8075 17.8275 64.0875 24.0275 ;
      RECT  55.8075 24.3775 64.0875 26.6475 ;
      RECT  23.3375 19.8775 23.6175 24.0275 ;
      RECT  23.3375 24.3775 23.6175 26.6475 ;
      RECT  23.6175 19.8775 34.495 24.0275 ;
      RECT  23.6175 24.3775 34.495 26.6475 ;
      RECT  36.3375 19.8775 55.8075 24.0275 ;
      RECT  36.3375 24.3775 55.8075 26.6475 ;
      RECT  34.91 19.8775 35.9225 24.0275 ;
      RECT  34.91 24.3775 35.9225 26.6475 ;
      RECT  35.9225 19.8775 36.3375 24.0275 ;
      RECT  35.9225 24.3775 36.3375 26.6475 ;
      RECT  34.495 19.8775 34.6275 24.0275 ;
      RECT  34.495 24.3775 34.6275 26.6475 ;
      RECT  34.6275 19.8775 34.91 24.0275 ;
      RECT  34.6275 24.3775 34.91 26.6475 ;
      RECT  0.56 1.38 2.285 9.845 ;
      RECT  0.56 9.845 2.285 10.26 ;
      RECT  0.56 10.26 2.285 10.95 ;
      RECT  2.285 1.38 2.7 9.845 ;
      RECT  2.285 10.26 2.7 10.95 ;
      RECT  2.7 1.38 8.755 9.845 ;
      RECT  2.7 9.845 8.755 10.26 ;
      RECT  2.7 10.26 8.755 10.95 ;
      RECT  34.91 83.02 70.8575 83.71 ;
      RECT  34.91 83.71 70.8575 83.845 ;
      RECT  70.8575 83.02 71.2725 83.71 ;
      RECT  71.2725 83.02 73.435 83.71 ;
      RECT  71.2725 83.71 73.435 83.845 ;
      RECT  12.765 36.91 13.18 39.485 ;
      RECT  12.765 39.9 13.18 40.98 ;
      RECT  77.81 42.89 78.225 45.465 ;
      RECT  77.81 45.88 78.225 82.605 ;
      RECT  9.17 41.395 12.765 42.475 ;
      RECT  9.17 42.475 12.765 42.89 ;
      RECT  9.17 42.89 12.765 46.57 ;
      RECT  12.765 41.395 13.18 42.475 ;
      RECT  13.18 41.395 14.2925 42.475 ;
      RECT  13.18 42.475 14.2925 42.89 ;
      RECT  13.18 42.89 14.2925 46.57 ;
      RECT  0.14 0.14 17.0525 0.275 ;
      RECT  17.4675 0.14 25.6325 0.275 ;
      RECT  12.765 42.89 13.18 45.465 ;
      RECT  12.765 45.88 13.18 46.57 ;
   LAYER  metal4 ;
      RECT  0.14 57.9125 67.16 83.845 ;
      RECT  67.16 0.14 67.86 27.2025 ;
      RECT  67.16 57.9125 67.86 83.845 ;
      RECT  0.14 45.3225 8.33 55.9025 ;
      RECT  0.14 55.9025 8.33 57.9125 ;
      RECT  8.33 27.2025 9.03 45.3225 ;
      RECT  8.33 55.9025 9.03 57.9125 ;
      RECT  22.05 27.2025 22.75 30.3725 ;
      RECT  22.05 54.9925 22.75 55.9025 ;
      RECT  22.75 27.2025 23.13 30.3725 ;
      RECT  22.75 30.3725 23.13 45.3225 ;
      RECT  22.75 45.3225 23.13 54.9925 ;
      RECT  22.75 54.9925 23.13 55.9025 ;
      RECT  11.05 0.14 11.75 12.1725 ;
      RECT  9.03 27.2025 11.05 27.6925 ;
      RECT  9.03 27.6925 11.05 30.3725 ;
      RECT  11.05 27.6925 11.75 30.3725 ;
      RECT  11.75 27.2025 22.05 27.6925 ;
      RECT  67.86 27.2025 68.24 30.3725 ;
      RECT  67.86 30.3725 68.24 54.9925 ;
      RECT  67.86 54.9925 68.24 57.9125 ;
      RECT  68.24 27.2025 68.94 30.3725 ;
      RECT  68.24 54.9925 68.94 57.9125 ;
      RECT  67.86 57.9125 79.435 59.9625 ;
      RECT  79.435 57.9125 80.135 59.9625 ;
      RECT  79.435 70.5425 80.135 83.845 ;
      RECT  67.86 59.9625 74.11 60.44 ;
      RECT  67.86 60.44 74.11 70.5425 ;
      RECT  74.11 59.9625 74.81 60.44 ;
      RECT  67.86 70.5425 74.11 80.9 ;
      RECT  67.86 80.9 74.11 83.845 ;
      RECT  74.11 80.9 74.81 83.845 ;
      RECT  82.155 0.14 82.855 20.4925 ;
      RECT  82.855 0.14 91.185 20.4925 ;
      RECT  82.855 20.4925 91.185 27.2025 ;
      RECT  82.855 27.2025 91.185 30.3725 ;
      RECT  82.155 31.0725 82.855 54.9925 ;
      RECT  82.855 30.3725 91.185 31.0725 ;
      RECT  18.8 55.0625 19.5 55.9025 ;
      RECT  19.5 55.0625 22.05 55.9025 ;
      RECT  16.18 0.14 16.88 4.285 ;
      RECT  16.88 0.14 67.16 4.285 ;
      RECT  16.88 4.285 67.16 12.1725 ;
      RECT  16.18 24.745 16.88 27.2025 ;
      RECT  16.88 12.1725 67.16 24.745 ;
      RECT  16.88 24.745 67.16 27.2025 ;
      RECT  90.9175 54.9925 91.185 57.9125 ;
      RECT  90.9175 57.9125 91.185 59.9625 ;
      RECT  90.2175 63.165 90.9175 70.5425 ;
      RECT  90.9175 59.9625 91.185 63.165 ;
      RECT  90.9175 63.165 91.185 70.5425 ;
      RECT  90.2175 31.0725 90.9175 40.2025 ;
      RECT  90.9175 31.0725 91.185 40.2025 ;
      RECT  90.9175 40.2025 91.185 54.9925 ;
      RECT  0.14 27.2025 0.4075 42.5125 ;
      RECT  0.14 42.5125 0.4075 45.3225 ;
      RECT  0.4075 42.5125 1.1075 45.3225 ;
      RECT  0.14 12.1725 0.4075 19.55 ;
      RECT  0.14 19.55 0.4075 27.2025 ;
      RECT  0.4075 12.1725 1.1075 19.55 ;
      RECT  68.94 55.0625 71.49 57.9125 ;
      RECT  71.49 55.0625 72.19 57.9125 ;
      RECT  74.81 59.9625 76.0525 60.3725 ;
      RECT  74.81 60.3725 76.0525 60.44 ;
      RECT  76.0525 59.9625 76.7525 60.3725 ;
      RECT  76.7525 59.9625 79.435 60.3725 ;
      RECT  76.7525 60.3725 79.435 60.44 ;
      RECT  74.81 60.44 76.0525 70.5425 ;
      RECT  76.7525 60.44 79.435 70.5425 ;
      RECT  74.81 70.5425 76.0525 80.9 ;
      RECT  76.7525 70.5425 79.435 80.9 ;
      RECT  74.81 80.9 76.0525 80.9675 ;
      RECT  74.81 80.9675 76.0525 83.845 ;
      RECT  76.0525 80.9675 76.7525 83.845 ;
      RECT  76.7525 80.9 79.435 80.9675 ;
      RECT  76.7525 80.9675 79.435 83.845 ;
      RECT  0.14 0.14 5.825 9.7025 ;
      RECT  0.14 9.7025 5.825 12.1725 ;
      RECT  5.825 0.14 6.525 9.7025 ;
      RECT  6.525 0.14 11.05 9.7025 ;
      RECT  6.525 9.7025 11.05 12.1725 ;
      RECT  1.1075 12.1725 5.825 19.55 ;
      RECT  6.525 12.1725 11.05 19.55 ;
      RECT  5.825 25.2225 6.525 27.2025 ;
      RECT  6.525 19.55 11.05 25.2225 ;
      RECT  6.525 25.2225 11.05 27.2025 ;
      RECT  9.03 55.9025 11.19 55.9675 ;
      RECT  9.03 55.9675 11.19 57.9125 ;
      RECT  11.19 55.9675 11.89 57.9125 ;
      RECT  11.89 55.9025 23.13 55.9675 ;
      RECT  11.89 55.9675 23.13 57.9125 ;
      RECT  9.03 30.3725 11.19 45.2575 ;
      RECT  9.03 45.2575 11.19 45.3225 ;
      RECT  11.19 30.3725 11.89 45.2575 ;
      RECT  9.03 45.3225 11.19 54.9925 ;
      RECT  9.03 54.9925 11.19 55.0625 ;
      RECT  9.03 55.0625 11.19 55.9025 ;
      RECT  11.89 55.0625 18.8 55.9025 ;
      RECT  68.94 27.2025 73.08 30.34 ;
      RECT  73.08 27.2025 73.78 30.34 ;
      RECT  72.19 30.3725 73.08 31.0725 ;
      RECT  72.19 31.0725 73.08 54.9925 ;
      RECT  72.19 54.9925 73.08 55.0625 ;
      RECT  68.94 30.3725 70.93 31.0725 ;
      RECT  68.94 31.0725 70.93 54.9925 ;
      RECT  68.94 54.9925 70.93 55.025 ;
      RECT  68.94 55.025 70.93 55.0625 ;
      RECT  70.93 55.025 71.49 55.0625 ;
      RECT  68.94 30.34 70.93 30.3725 ;
      RECT  71.63 30.34 73.08 30.3725 ;
      RECT  1.1075 27.2025 2.47 42.5125 ;
      RECT  3.17 27.2025 8.33 42.5125 ;
      RECT  1.1075 42.5125 2.47 42.545 ;
      RECT  1.1075 42.545 2.47 45.3225 ;
      RECT  2.47 42.545 3.17 45.3225 ;
      RECT  3.17 42.5125 8.33 42.545 ;
      RECT  3.17 42.545 8.33 45.3225 ;
      RECT  1.1075 19.55 2.47 19.5825 ;
      RECT  1.1075 19.5825 2.47 25.2225 ;
      RECT  2.47 19.55 3.17 19.5825 ;
      RECT  3.17 19.55 5.825 19.5825 ;
      RECT  3.17 19.5825 5.825 25.2225 ;
      RECT  1.1075 25.2225 2.47 27.2025 ;
      RECT  3.17 25.2225 5.825 27.2025 ;
      RECT  24.29 55.9025 66.7 57.9125 ;
      RECT  24.29 27.2025 66.7 30.3725 ;
      RECT  24.29 30.3725 66.7 45.3225 ;
      RECT  24.29 45.3225 66.7 54.9925 ;
      RECT  24.29 54.9925 66.7 55.9025 ;
      RECT  11.75 27.6925 19.36 30.34 ;
      RECT  19.36 27.6925 20.06 30.34 ;
      RECT  20.06 27.6925 22.05 30.34 ;
      RECT  20.06 30.34 22.05 30.3725 ;
      RECT  20.06 30.3725 22.05 45.3225 ;
      RECT  20.06 45.3225 22.05 54.9925 ;
      RECT  19.5 55.025 20.06 55.0625 ;
      RECT  20.06 54.9925 22.05 55.025 ;
      RECT  20.06 55.025 22.05 55.0625 ;
      RECT  11.89 30.3725 17.21 45.2575 ;
      RECT  17.91 30.3725 18.8 45.2575 ;
      RECT  11.89 45.2575 17.21 45.3225 ;
      RECT  17.91 45.2575 18.8 45.3225 ;
      RECT  11.89 45.3225 17.21 54.9925 ;
      RECT  17.91 45.3225 18.8 54.9925 ;
      RECT  11.89 54.9925 17.21 55.0625 ;
      RECT  17.91 54.9925 18.8 55.0625 ;
      RECT  11.75 30.34 17.21 30.3725 ;
      RECT  17.91 30.34 19.36 30.3725 ;
      RECT  88.855 57.9125 90.2175 59.9625 ;
      RECT  88.155 63.1325 88.855 63.165 ;
      RECT  88.855 59.9625 90.2175 63.1325 ;
      RECT  88.855 63.1325 90.2175 63.165 ;
      RECT  82.855 31.0725 88.155 40.17 ;
      RECT  82.855 40.17 88.155 40.2025 ;
      RECT  88.155 31.0725 88.855 40.17 ;
      RECT  88.855 31.0725 90.2175 40.17 ;
      RECT  88.855 40.17 90.2175 40.2025 ;
      RECT  82.855 40.2025 88.155 54.9925 ;
      RECT  88.855 40.2025 90.2175 54.9925 ;
      RECT  88.855 55.0625 90.2175 57.9125 ;
      RECT  73.78 54.9925 88.155 55.0625 ;
      RECT  88.855 54.9925 90.2175 55.0625 ;
      RECT  80.135 70.5425 84.66 73.0125 ;
      RECT  80.135 73.0125 84.66 83.845 ;
      RECT  84.66 73.0125 85.36 83.845 ;
      RECT  85.36 70.5425 91.185 73.0125 ;
      RECT  85.36 73.0125 91.185 83.845 ;
      RECT  80.135 63.165 84.66 70.5425 ;
      RECT  85.36 63.165 90.2175 70.5425 ;
      RECT  80.135 57.9125 84.66 59.9625 ;
      RECT  85.36 57.9125 88.155 59.9625 ;
      RECT  80.135 59.9625 84.66 63.1325 ;
      RECT  85.36 59.9625 88.155 63.1325 ;
      RECT  80.135 63.1325 84.66 63.165 ;
      RECT  85.36 63.1325 88.155 63.165 ;
      RECT  72.19 55.0625 84.66 57.4925 ;
      RECT  72.19 57.4925 84.66 57.9125 ;
      RECT  84.66 55.0625 85.36 57.4925 ;
      RECT  85.36 55.0625 88.155 57.4925 ;
      RECT  85.36 57.4925 88.155 57.9125 ;
      RECT  11.75 0.14 14.2375 4.2175 ;
      RECT  11.75 4.2175 14.2375 4.285 ;
      RECT  14.2375 0.14 14.9375 4.2175 ;
      RECT  14.9375 0.14 16.18 4.2175 ;
      RECT  14.9375 4.2175 16.18 4.285 ;
      RECT  11.75 4.285 14.2375 12.1725 ;
      RECT  14.9375 4.285 16.18 12.1725 ;
      RECT  11.75 12.1725 14.2375 24.745 ;
      RECT  14.9375 12.1725 16.18 24.745 ;
      RECT  11.75 24.745 14.2375 24.8125 ;
      RECT  11.75 24.8125 14.2375 27.2025 ;
      RECT  14.2375 24.8125 14.9375 27.2025 ;
      RECT  14.9375 24.745 16.18 24.8125 ;
      RECT  14.9375 24.8125 16.18 27.2025 ;
      RECT  67.86 0.14 79.295 20.4275 ;
      RECT  67.86 20.4275 79.295 20.4925 ;
      RECT  79.295 0.14 79.995 20.4275 ;
      RECT  79.995 0.14 82.155 20.4275 ;
      RECT  79.995 20.4275 82.155 20.4925 ;
      RECT  67.86 20.4925 79.295 27.2025 ;
      RECT  79.995 20.4925 82.155 27.2025 ;
      RECT  73.78 27.2025 79.295 30.34 ;
      RECT  79.995 27.2025 82.155 30.34 ;
      RECT  73.78 30.34 79.295 30.3725 ;
      RECT  79.995 30.34 82.155 30.3725 ;
      RECT  73.78 30.3725 79.295 31.0725 ;
      RECT  79.995 30.3725 82.155 31.0725 ;
      RECT  73.78 31.0725 79.295 31.1375 ;
      RECT  73.78 31.1375 79.295 54.9925 ;
      RECT  79.295 31.1375 79.995 54.9925 ;
      RECT  79.995 31.0725 82.155 31.1375 ;
      RECT  79.995 31.1375 82.155 54.9925 ;
   END
END    freepdk45_sram_1w1r_128x4_1
END    LIBRARY
