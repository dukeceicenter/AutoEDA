../macros/freepdk45_sram_1w1r_28x128_32/freepdk45_sram_1w1r_28x128_32.lef