../macros/freepdk45_sram_1w1r_40x240/freepdk45_sram_1w1r_40x240.lef