/home/yl996/proj/mcp-eda-example/libraries/FreePDK45/OpenRAM/macros/freepdk45_sram_1rw0r_64x40_20/freepdk45_sram_1rw0r_64x40_20.lef