VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1rw0r_64x176_22
   CLASS BLOCK ;
   SIZE 579.145 BY 146.8275 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.0 1.105 76.135 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.86 1.105 78.995 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.72 1.105 81.855 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.58 1.105 84.715 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.44 1.105 87.575 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.3 1.105 90.435 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.16 1.105 93.295 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.02 1.105 96.155 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.88 1.105 99.015 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.74 1.105 101.875 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.6 1.105 104.735 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.46 1.105 107.595 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.32 1.105 110.455 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.18 1.105 113.315 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.04 1.105 116.175 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.9 1.105 119.035 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.76 1.105 121.895 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.62 1.105 124.755 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.48 1.105 127.615 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.34 1.105 130.475 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.2 1.105 133.335 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.06 1.105 136.195 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.92 1.105 139.055 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.78 1.105 141.915 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.64 1.105 144.775 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.5 1.105 147.635 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.36 1.105 150.495 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.22 1.105 153.355 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.08 1.105 156.215 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.94 1.105 159.075 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.8 1.105 161.935 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.66 1.105 164.795 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.52 1.105 167.655 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.38 1.105 170.515 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.24 1.105 173.375 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.1 1.105 176.235 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.96 1.105 179.095 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.82 1.105 181.955 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.68 1.105 184.815 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.54 1.105 187.675 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.4 1.105 190.535 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.26 1.105 193.395 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.12 1.105 196.255 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.98 1.105 199.115 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.84 1.105 201.975 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.7 1.105 204.835 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.56 1.105 207.695 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.42 1.105 210.555 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.28 1.105 213.415 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.14 1.105 216.275 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.0 1.105 219.135 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.86 1.105 221.995 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.72 1.105 224.855 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.58 1.105 227.715 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.44 1.105 230.575 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.3 1.105 233.435 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.16 1.105 236.295 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.02 1.105 239.155 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.88 1.105 242.015 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.74 1.105 244.875 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.6 1.105 247.735 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.46 1.105 250.595 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.32 1.105 253.455 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.18 1.105 256.315 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.04 1.105 259.175 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.9 1.105 262.035 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.76 1.105 264.895 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.62 1.105 267.755 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.48 1.105 270.615 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.34 1.105 273.475 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.2 1.105 276.335 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.06 1.105 279.195 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.92 1.105 282.055 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.78 1.105 284.915 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.64 1.105 287.775 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.5 1.105 290.635 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.36 1.105 293.495 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.22 1.105 296.355 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.08 1.105 299.215 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.94 1.105 302.075 1.24 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.8 1.105 304.935 1.24 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.66 1.105 307.795 1.24 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.52 1.105 310.655 1.24 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.38 1.105 313.515 1.24 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.24 1.105 316.375 1.24 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.1 1.105 319.235 1.24 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.96 1.105 322.095 1.24 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.82 1.105 324.955 1.24 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.68 1.105 327.815 1.24 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.54 1.105 330.675 1.24 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.4 1.105 333.535 1.24 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.26 1.105 336.395 1.24 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.12 1.105 339.255 1.24 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.98 1.105 342.115 1.24 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.84 1.105 344.975 1.24 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.7 1.105 347.835 1.24 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.56 1.105 350.695 1.24 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.42 1.105 353.555 1.24 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.28 1.105 356.415 1.24 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.14 1.105 359.275 1.24 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.0 1.105 362.135 1.24 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.86 1.105 364.995 1.24 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.72 1.105 367.855 1.24 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.58 1.105 370.715 1.24 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.44 1.105 373.575 1.24 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  376.3 1.105 376.435 1.24 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  379.16 1.105 379.295 1.24 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  382.02 1.105 382.155 1.24 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.88 1.105 385.015 1.24 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  387.74 1.105 387.875 1.24 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  390.6 1.105 390.735 1.24 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.46 1.105 393.595 1.24 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.32 1.105 396.455 1.24 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.18 1.105 399.315 1.24 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  402.04 1.105 402.175 1.24 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.9 1.105 405.035 1.24 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.76 1.105 407.895 1.24 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.62 1.105 410.755 1.24 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  413.48 1.105 413.615 1.24 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  416.34 1.105 416.475 1.24 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  419.2 1.105 419.335 1.24 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  422.06 1.105 422.195 1.24 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.92 1.105 425.055 1.24 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.78 1.105 427.915 1.24 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  430.64 1.105 430.775 1.24 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  433.5 1.105 433.635 1.24 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  436.36 1.105 436.495 1.24 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  439.22 1.105 439.355 1.24 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  442.08 1.105 442.215 1.24 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.94 1.105 445.075 1.24 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.8 1.105 447.935 1.24 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  450.66 1.105 450.795 1.24 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.52 1.105 453.655 1.24 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  456.38 1.105 456.515 1.24 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  459.24 1.105 459.375 1.24 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  462.1 1.105 462.235 1.24 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.96 1.105 465.095 1.24 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.82 1.105 467.955 1.24 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.68 1.105 470.815 1.24 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  473.54 1.105 473.675 1.24 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  476.4 1.105 476.535 1.24 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  479.26 1.105 479.395 1.24 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.12 1.105 482.255 1.24 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.98 1.105 485.115 1.24 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.84 1.105 487.975 1.24 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  490.7 1.105 490.835 1.24 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  493.56 1.105 493.695 1.24 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  496.42 1.105 496.555 1.24 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  499.28 1.105 499.415 1.24 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  502.14 1.105 502.275 1.24 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  505.0 1.105 505.135 1.24 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.86 1.105 507.995 1.24 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.72 1.105 510.855 1.24 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  513.58 1.105 513.715 1.24 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  516.44 1.105 516.575 1.24 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  519.3 1.105 519.435 1.24 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  522.16 1.105 522.295 1.24 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  525.02 1.105 525.155 1.24 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.88 1.105 528.015 1.24 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  530.74 1.105 530.875 1.24 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  533.6 1.105 533.735 1.24 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  536.46 1.105 536.595 1.24 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  539.32 1.105 539.455 1.24 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  542.18 1.105 542.315 1.24 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  545.04 1.105 545.175 1.24 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  547.9 1.105 548.035 1.24 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  550.76 1.105 550.895 1.24 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  553.62 1.105 553.755 1.24 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  556.48 1.105 556.615 1.24 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  559.34 1.105 559.475 1.24 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  562.2 1.105 562.335 1.24 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  565.06 1.105 565.195 1.24 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  567.92 1.105 568.055 1.24 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  570.78 1.105 570.915 1.24 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  573.64 1.105 573.775 1.24 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  576.5 1.105 576.635 1.24 ;
      END
   END din0[175]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.4 80.7825 47.535 80.9175 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.4 83.5125 47.535 83.6475 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.4 85.7225 47.535 85.8575 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.4 88.4525 47.535 88.5875 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.4 90.6625 47.535 90.7975 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.4 93.3925 47.535 93.5275 ;
      END
   END addr0[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 36.0625 0.42 36.1975 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 38.7925 0.42 38.9275 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 36.1475 6.6625 36.2825 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.12 1.105 53.255 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.98 1.105 56.115 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.84 1.105 58.975 1.24 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.7 1.105 61.835 1.24 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.56 1.105 64.695 1.24 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.42 1.105 67.555 1.24 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.28 1.105 70.415 1.24 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.14 1.105 73.275 1.24 ;
      END
   END wmask0[7]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.1125 47.7125 73.2475 47.8475 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.8175 47.7125 73.9525 47.8475 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.5225 47.7125 74.6575 47.8475 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.2275 47.7125 75.3625 47.8475 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.9325 47.7125 76.0675 47.8475 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.6375 47.7125 76.7725 47.8475 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.3425 47.7125 77.4775 47.8475 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.0475 47.7125 78.1825 47.8475 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.7525 47.7125 78.8875 47.8475 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.4575 47.7125 79.5925 47.8475 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.1625 47.7125 80.2975 47.8475 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.8675 47.7125 81.0025 47.8475 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.5725 47.7125 81.7075 47.8475 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.2775 47.7125 82.4125 47.8475 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.9825 47.7125 83.1175 47.8475 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.6875 47.7125 83.8225 47.8475 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.3925 47.7125 84.5275 47.8475 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.0975 47.7125 85.2325 47.8475 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.8025 47.7125 85.9375 47.8475 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.5075 47.7125 86.6425 47.8475 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.2125 47.7125 87.3475 47.8475 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.9175 47.7125 88.0525 47.8475 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.6225 47.7125 88.7575 47.8475 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.3275 47.7125 89.4625 47.8475 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.0325 47.7125 90.1675 47.8475 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.7375 47.7125 90.8725 47.8475 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.4425 47.7125 91.5775 47.8475 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.1475 47.7125 92.2825 47.8475 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.8525 47.7125 92.9875 47.8475 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.5575 47.7125 93.6925 47.8475 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.2625 47.7125 94.3975 47.8475 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.9675 47.7125 95.1025 47.8475 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.6725 47.7125 95.8075 47.8475 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.3775 47.7125 96.5125 47.8475 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.0825 47.7125 97.2175 47.8475 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.7875 47.7125 97.9225 47.8475 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.4925 47.7125 98.6275 47.8475 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.1975 47.7125 99.3325 47.8475 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.9025 47.7125 100.0375 47.8475 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.6075 47.7125 100.7425 47.8475 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.3125 47.7125 101.4475 47.8475 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.0175 47.7125 102.1525 47.8475 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.7225 47.7125 102.8575 47.8475 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.4275 47.7125 103.5625 47.8475 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.1325 47.7125 104.2675 47.8475 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.8375 47.7125 104.9725 47.8475 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.5425 47.7125 105.6775 47.8475 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.2475 47.7125 106.3825 47.8475 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.9525 47.7125 107.0875 47.8475 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.6575 47.7125 107.7925 47.8475 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.3625 47.7125 108.4975 47.8475 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.0675 47.7125 109.2025 47.8475 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.7725 47.7125 109.9075 47.8475 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.4775 47.7125 110.6125 47.8475 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.1825 47.7125 111.3175 47.8475 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.8875 47.7125 112.0225 47.8475 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.5925 47.7125 112.7275 47.8475 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.2975 47.7125 113.4325 47.8475 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.0025 47.7125 114.1375 47.8475 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.7075 47.7125 114.8425 47.8475 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.4125 47.7125 115.5475 47.8475 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.1175 47.7125 116.2525 47.8475 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.8225 47.7125 116.9575 47.8475 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.5275 47.7125 117.6625 47.8475 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.2325 47.7125 118.3675 47.8475 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.9375 47.7125 119.0725 47.8475 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.6425 47.7125 119.7775 47.8475 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.3475 47.7125 120.4825 47.8475 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.0525 47.7125 121.1875 47.8475 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.7575 47.7125 121.8925 47.8475 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.4625 47.7125 122.5975 47.8475 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.1675 47.7125 123.3025 47.8475 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.8725 47.7125 124.0075 47.8475 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.5775 47.7125 124.7125 47.8475 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.2825 47.7125 125.4175 47.8475 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.9875 47.7125 126.1225 47.8475 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.6925 47.7125 126.8275 47.8475 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.3975 47.7125 127.5325 47.8475 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.1025 47.7125 128.2375 47.8475 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.8075 47.7125 128.9425 47.8475 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.5125 47.7125 129.6475 47.8475 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.2175 47.7125 130.3525 47.8475 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.9225 47.7125 131.0575 47.8475 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.6275 47.7125 131.7625 47.8475 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.3325 47.7125 132.4675 47.8475 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.0375 47.7125 133.1725 47.8475 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.7425 47.7125 133.8775 47.8475 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.4475 47.7125 134.5825 47.8475 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.1525 47.7125 135.2875 47.8475 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.8575 47.7125 135.9925 47.8475 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.5625 47.7125 136.6975 47.8475 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.2675 47.7125 137.4025 47.8475 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.9725 47.7125 138.1075 47.8475 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.6775 47.7125 138.8125 47.8475 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.3825 47.7125 139.5175 47.8475 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.0875 47.7125 140.2225 47.8475 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.7925 47.7125 140.9275 47.8475 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.4975 47.7125 141.6325 47.8475 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.2025 47.7125 142.3375 47.8475 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.9075 47.7125 143.0425 47.8475 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.6125 47.7125 143.7475 47.8475 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.3175 47.7125 144.4525 47.8475 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.0225 47.7125 145.1575 47.8475 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.7275 47.7125 145.8625 47.8475 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.4325 47.7125 146.5675 47.8475 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.1375 47.7125 147.2725 47.8475 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.8425 47.7125 147.9775 47.8475 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.5475 47.7125 148.6825 47.8475 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.2525 47.7125 149.3875 47.8475 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.9575 47.7125 150.0925 47.8475 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.6625 47.7125 150.7975 47.8475 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.3675 47.7125 151.5025 47.8475 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.0725 47.7125 152.2075 47.8475 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.7775 47.7125 152.9125 47.8475 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.4825 47.7125 153.6175 47.8475 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.1875 47.7125 154.3225 47.8475 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.8925 47.7125 155.0275 47.8475 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.5975 47.7125 155.7325 47.8475 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.3025 47.7125 156.4375 47.8475 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.0075 47.7125 157.1425 47.8475 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.7125 47.7125 157.8475 47.8475 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.4175 47.7125 158.5525 47.8475 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.1225 47.7125 159.2575 47.8475 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.8275 47.7125 159.9625 47.8475 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.5325 47.7125 160.6675 47.8475 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.2375 47.7125 161.3725 47.8475 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.9425 47.7125 162.0775 47.8475 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.6475 47.7125 162.7825 47.8475 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.3525 47.7125 163.4875 47.8475 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.0575 47.7125 164.1925 47.8475 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.7625 47.7125 164.8975 47.8475 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.4675 47.7125 165.6025 47.8475 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.1725 47.7125 166.3075 47.8475 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.8775 47.7125 167.0125 47.8475 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.5825 47.7125 167.7175 47.8475 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.2875 47.7125 168.4225 47.8475 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.9925 47.7125 169.1275 47.8475 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.6975 47.7125 169.8325 47.8475 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.4025 47.7125 170.5375 47.8475 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.1075 47.7125 171.2425 47.8475 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.8125 47.7125 171.9475 47.8475 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.5175 47.7125 172.6525 47.8475 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.2225 47.7125 173.3575 47.8475 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.9275 47.7125 174.0625 47.8475 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.6325 47.7125 174.7675 47.8475 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.3375 47.7125 175.4725 47.8475 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.0425 47.7125 176.1775 47.8475 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.7475 47.7125 176.8825 47.8475 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.4525 47.7125 177.5875 47.8475 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.1575 47.7125 178.2925 47.8475 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.8625 47.7125 178.9975 47.8475 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.5675 47.7125 179.7025 47.8475 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.2725 47.7125 180.4075 47.8475 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.9775 47.7125 181.1125 47.8475 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.6825 47.7125 181.8175 47.8475 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.3875 47.7125 182.5225 47.8475 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.0925 47.7125 183.2275 47.8475 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.7975 47.7125 183.9325 47.8475 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.5025 47.7125 184.6375 47.8475 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.2075 47.7125 185.3425 47.8475 ;
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.9125 47.7125 186.0475 47.8475 ;
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.6175 47.7125 186.7525 47.8475 ;
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.3225 47.7125 187.4575 47.8475 ;
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.0275 47.7125 188.1625 47.8475 ;
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.7325 47.7125 188.8675 47.8475 ;
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.4375 47.7125 189.5725 47.8475 ;
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.1425 47.7125 190.2775 47.8475 ;
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.8475 47.7125 190.9825 47.8475 ;
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.5525 47.7125 191.6875 47.8475 ;
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.2575 47.7125 192.3925 47.8475 ;
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.9625 47.7125 193.0975 47.8475 ;
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.6675 47.7125 193.8025 47.8475 ;
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.3725 47.7125 194.5075 47.8475 ;
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.0775 47.7125 195.2125 47.8475 ;
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.7825 47.7125 195.9175 47.8475 ;
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.4875 47.7125 196.6225 47.8475 ;
      END
   END dout0[175]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  53.2175 67.3925 53.3525 67.5275 ;
         LAYER metal3 ;
         RECT  418.9175 2.47 419.0525 2.605 ;
         LAYER metal3 ;
         RECT  338.8375 2.47 338.9725 2.605 ;
         LAYER metal3 ;
         RECT  110.0375 2.47 110.1725 2.605 ;
         LAYER metal3 ;
         RECT  53.2175 75.5825 53.3525 75.7175 ;
         LAYER metal3 ;
         RECT  75.7175 2.47 75.8525 2.605 ;
         LAYER metal3 ;
         RECT  53.2175 59.2025 53.3525 59.3375 ;
         LAYER metal3 ;
         RECT  247.3175 2.47 247.4525 2.605 ;
         LAYER metal3 ;
         RECT  70.8675 50.3325 197.2925 50.4025 ;
         LAYER metal3 ;
         RECT  53.2175 61.9325 53.3525 62.0675 ;
         LAYER metal3 ;
         RECT  155.7975 2.47 155.9325 2.605 ;
         LAYER metal3 ;
         RECT  212.9975 2.47 213.1325 2.605 ;
         LAYER metal3 ;
         RECT  407.4775 2.47 407.6125 2.605 ;
         LAYER metal3 ;
         RECT  52.8375 2.47 52.9725 2.605 ;
         LAYER metal3 ;
         RECT  315.9575 2.47 316.0925 2.605 ;
         LAYER metal3 ;
         RECT  521.8775 2.47 522.0125 2.605 ;
         LAYER metal3 ;
         RECT  258.7575 2.47 258.8925 2.605 ;
         LAYER metal3 ;
         RECT  69.7225 56.4725 69.8575 56.6075 ;
         LAYER metal4 ;
         RECT  0.0 34.955 0.14 40.035 ;
         LAYER metal3 ;
         RECT  350.2775 2.47 350.4125 2.605 ;
         LAYER metal3 ;
         RECT  453.2375 2.47 453.3725 2.605 ;
         LAYER metal3 ;
         RECT  327.3975 2.47 327.5325 2.605 ;
         LAYER metal3 ;
         RECT  304.5175 2.47 304.6525 2.605 ;
         LAYER metal3 ;
         RECT  293.0775 2.47 293.2125 2.605 ;
         LAYER metal4 ;
         RECT  0.6875 44.8025 0.8275 67.205 ;
         LAYER metal3 ;
         RECT  281.6375 2.47 281.7725 2.605 ;
         LAYER metal3 ;
         RECT  224.4375 2.47 224.5725 2.605 ;
         LAYER metal3 ;
         RECT  87.1575 2.47 87.2925 2.605 ;
         LAYER metal3 ;
         RECT  201.5575 2.47 201.6925 2.605 ;
         LAYER metal3 ;
         RECT  544.7575 2.47 544.8925 2.605 ;
         LAYER metal3 ;
         RECT  441.7975 2.47 441.9325 2.605 ;
         LAYER metal3 ;
         RECT  70.8675 43.405 197.2925 43.475 ;
         LAYER metal3 ;
         RECT  270.1975 2.47 270.3325 2.605 ;
         LAYER metal4 ;
         RECT  58.77 57.835 58.91 145.405 ;
         LAYER metal4 ;
         RECT  70.8 54.925 70.94 146.63 ;
         LAYER metal3 ;
         RECT  98.5975 2.47 98.7325 2.605 ;
         LAYER metal3 ;
         RECT  132.9175 2.47 133.0525 2.605 ;
         LAYER metal3 ;
         RECT  567.6375 2.47 567.7725 2.605 ;
         LAYER metal3 ;
         RECT  487.5575 2.47 487.6925 2.605 ;
         LAYER metal3 ;
         RECT  70.7325 42.4375 70.8675 42.5725 ;
         LAYER metal3 ;
         RECT  235.8775 2.47 236.0125 2.605 ;
         LAYER metal3 ;
         RECT  533.3175 2.47 533.4525 2.605 ;
         LAYER metal3 ;
         RECT  384.5975 2.47 384.7325 2.605 ;
         LAYER metal3 ;
         RECT  556.1975 2.47 556.3325 2.605 ;
         LAYER metal3 ;
         RECT  373.1575 2.47 373.2925 2.605 ;
         LAYER metal3 ;
         RECT  167.2375 2.47 167.3725 2.605 ;
         LAYER metal3 ;
         RECT  396.0375 2.47 396.1725 2.605 ;
         LAYER metal4 ;
         RECT  69.72 57.835 69.86 145.335 ;
         LAYER metal3 ;
         RECT  70.8675 54.23 197.2925 54.3 ;
         LAYER metal3 ;
         RECT  498.9975 2.47 499.1325 2.605 ;
         LAYER metal3 ;
         RECT  510.4375 2.47 510.5725 2.605 ;
         LAYER metal3 ;
         RECT  464.6775 2.47 464.8125 2.605 ;
         LAYER metal3 ;
         RECT  190.1175 2.47 190.2525 2.605 ;
         LAYER metal3 ;
         RECT  144.3575 2.47 144.4925 2.605 ;
         LAYER metal3 ;
         RECT  361.7175 2.47 361.8525 2.605 ;
         LAYER metal4 ;
         RECT  49.835 37.425 49.975 52.385 ;
         LAYER metal3 ;
         RECT  64.2775 2.47 64.4125 2.605 ;
         LAYER metal3 ;
         RECT  121.4775 2.47 121.6125 2.605 ;
         LAYER metal4 ;
         RECT  47.115 79.675 47.255 94.635 ;
         LAYER metal3 ;
         RECT  53.2175 70.1225 53.3525 70.2575 ;
         LAYER metal3 ;
         RECT  430.3575 2.47 430.4925 2.605 ;
         LAYER metal3 ;
         RECT  178.6775 2.47 178.8125 2.605 ;
         LAYER metal3 ;
         RECT  53.2175 78.3125 53.3525 78.4475 ;
         LAYER metal4 ;
         RECT  198.725 54.925 198.865 146.63 ;
         LAYER metal3 ;
         RECT  59.39 57.13 59.525 57.265 ;
         LAYER metal3 ;
         RECT  476.1175 2.47 476.2525 2.605 ;
         LAYER metal3 ;
         RECT  197.1575 42.4375 197.2925 42.5725 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  147.2175 0.0 147.3525 0.135 ;
         LAYER metal3 ;
         RECT  398.8975 0.0 399.0325 0.135 ;
         LAYER metal3 ;
         RECT  158.6575 0.0 158.7925 0.135 ;
         LAYER metal3 ;
         RECT  170.0975 0.0 170.2325 0.135 ;
         LAYER metal3 ;
         RECT  250.1775 0.0 250.3125 0.135 ;
         LAYER metal3 ;
         RECT  387.4575 0.0 387.5925 0.135 ;
         LAYER metal4 ;
         RECT  71.26 54.925 71.4 146.63 ;
         LAYER metal3 ;
         RECT  559.0575 0.0 559.1925 0.135 ;
         LAYER metal3 ;
         RECT  51.69 71.4875 51.825 71.6225 ;
         LAYER metal4 ;
         RECT  4.845 34.89 4.985 40.1 ;
         LAYER metal3 ;
         RECT  101.4575 0.0 101.5925 0.135 ;
         LAYER metal3 ;
         RECT  284.4975 0.0 284.6325 0.135 ;
         LAYER metal3 ;
         RECT  51.69 74.2175 51.825 74.3525 ;
         LAYER metal3 ;
         RECT  51.69 68.7575 51.825 68.8925 ;
         LAYER metal3 ;
         RECT  421.7775 0.0 421.9125 0.135 ;
         LAYER metal3 ;
         RECT  330.2575 0.0 330.3925 0.135 ;
         LAYER metal3 ;
         RECT  238.7375 0.0 238.8725 0.135 ;
         LAYER metal4 ;
         RECT  59.33 57.8025 59.47 145.3675 ;
         LAYER metal3 ;
         RECT  215.8575 0.0 215.9925 0.135 ;
         LAYER metal3 ;
         RECT  90.0175 0.0 90.1525 0.135 ;
         LAYER metal3 ;
         RECT  456.0975 0.0 456.2325 0.135 ;
         LAYER metal3 ;
         RECT  197.1575 40.6175 197.2925 40.7525 ;
         LAYER metal3 ;
         RECT  55.6975 0.0 55.8325 0.135 ;
         LAYER metal3 ;
         RECT  67.1375 0.0 67.2725 0.135 ;
         LAYER metal3 ;
         RECT  536.1775 0.0 536.3125 0.135 ;
         LAYER metal3 ;
         RECT  433.2175 0.0 433.3525 0.135 ;
         LAYER metal3 ;
         RECT  181.5375 0.0 181.6725 0.135 ;
         LAYER metal3 ;
         RECT  51.69 63.2975 51.825 63.4325 ;
         LAYER metal4 ;
         RECT  49.975 79.61 50.115 94.7 ;
         LAYER metal4 ;
         RECT  6.385 34.955 6.525 54.855 ;
         LAYER metal3 ;
         RECT  51.69 79.6775 51.825 79.8125 ;
         LAYER metal3 ;
         RECT  547.6175 0.0 547.7525 0.135 ;
         LAYER metal3 ;
         RECT  112.8975 0.0 113.0325 0.135 ;
         LAYER metal3 ;
         RECT  135.7775 0.0 135.9125 0.135 ;
         LAYER metal3 ;
         RECT  490.4175 0.0 490.5525 0.135 ;
         LAYER metal3 ;
         RECT  376.0175 0.0 376.1525 0.135 ;
         LAYER metal3 ;
         RECT  192.9775 0.0 193.1125 0.135 ;
         LAYER metal3 ;
         RECT  51.69 60.5675 51.825 60.7025 ;
         LAYER metal3 ;
         RECT  70.8675 52.225 197.3275 52.295 ;
         LAYER metal3 ;
         RECT  478.9775 0.0 479.1125 0.135 ;
         LAYER metal3 ;
         RECT  51.69 76.9475 51.825 77.0825 ;
         LAYER metal3 ;
         RECT  70.8675 45.455 197.2925 45.525 ;
         LAYER metal3 ;
         RECT  341.6975 0.0 341.8325 0.135 ;
         LAYER metal3 ;
         RECT  467.5375 0.0 467.6725 0.135 ;
         LAYER metal3 ;
         RECT  273.0575 0.0 273.1925 0.135 ;
         LAYER metal3 ;
         RECT  78.5775 0.0 78.7125 0.135 ;
         LAYER metal3 ;
         RECT  501.8575 0.0 501.9925 0.135 ;
         LAYER metal3 ;
         RECT  353.1375 0.0 353.2725 0.135 ;
         LAYER metal3 ;
         RECT  513.2975 0.0 513.4325 0.135 ;
         LAYER metal3 ;
         RECT  410.3375 0.0 410.4725 0.135 ;
         LAYER metal3 ;
         RECT  364.5775 0.0 364.7125 0.135 ;
         LAYER metal4 ;
         RECT  56.835 57.8025 56.975 145.405 ;
         LAYER metal3 ;
         RECT  204.4175 0.0 204.5525 0.135 ;
         LAYER metal3 ;
         RECT  51.69 66.0275 51.825 66.1625 ;
         LAYER metal4 ;
         RECT  198.265 54.925 198.405 146.63 ;
         LAYER metal3 ;
         RECT  524.7375 0.0 524.8725 0.135 ;
         LAYER metal4 ;
         RECT  2.75 44.835 2.89 67.2375 ;
         LAYER metal3 ;
         RECT  295.9375 0.0 296.0725 0.135 ;
         LAYER metal3 ;
         RECT  444.6575 0.0 444.7925 0.135 ;
         LAYER metal3 ;
         RECT  124.3375 0.0 124.4725 0.135 ;
         LAYER metal3 ;
         RECT  307.3775 0.0 307.5125 0.135 ;
         LAYER metal3 ;
         RECT  70.7325 40.6175 70.8675 40.7525 ;
         LAYER metal3 ;
         RECT  318.8175 0.0 318.9525 0.135 ;
         LAYER metal3 ;
         RECT  51.69 57.8375 51.825 57.9725 ;
         LAYER metal3 ;
         RECT  227.2975 0.0 227.4325 0.135 ;
         LAYER metal3 ;
         RECT  570.4975 0.0 570.6325 0.135 ;
         LAYER metal3 ;
         RECT  261.6175 0.0 261.7525 0.135 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 579.005 146.6875 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 579.005 146.6875 ;
   LAYER  metal3 ;
      RECT  75.86 0.14 76.275 0.965 ;
      RECT  76.275 0.965 78.72 1.38 ;
      RECT  79.135 0.965 81.58 1.38 ;
      RECT  81.995 0.965 84.44 1.38 ;
      RECT  84.855 0.965 87.3 1.38 ;
      RECT  87.715 0.965 90.16 1.38 ;
      RECT  90.575 0.965 93.02 1.38 ;
      RECT  93.435 0.965 95.88 1.38 ;
      RECT  96.295 0.965 98.74 1.38 ;
      RECT  99.155 0.965 101.6 1.38 ;
      RECT  102.015 0.965 104.46 1.38 ;
      RECT  104.875 0.965 107.32 1.38 ;
      RECT  107.735 0.965 110.18 1.38 ;
      RECT  110.595 0.965 113.04 1.38 ;
      RECT  113.455 0.965 115.9 1.38 ;
      RECT  116.315 0.965 118.76 1.38 ;
      RECT  119.175 0.965 121.62 1.38 ;
      RECT  122.035 0.965 124.48 1.38 ;
      RECT  124.895 0.965 127.34 1.38 ;
      RECT  127.755 0.965 130.2 1.38 ;
      RECT  130.615 0.965 133.06 1.38 ;
      RECT  133.475 0.965 135.92 1.38 ;
      RECT  136.335 0.965 138.78 1.38 ;
      RECT  139.195 0.965 141.64 1.38 ;
      RECT  142.055 0.965 144.5 1.38 ;
      RECT  144.915 0.965 147.36 1.38 ;
      RECT  147.775 0.965 150.22 1.38 ;
      RECT  150.635 0.965 153.08 1.38 ;
      RECT  153.495 0.965 155.94 1.38 ;
      RECT  156.355 0.965 158.8 1.38 ;
      RECT  159.215 0.965 161.66 1.38 ;
      RECT  162.075 0.965 164.52 1.38 ;
      RECT  164.935 0.965 167.38 1.38 ;
      RECT  167.795 0.965 170.24 1.38 ;
      RECT  170.655 0.965 173.1 1.38 ;
      RECT  173.515 0.965 175.96 1.38 ;
      RECT  176.375 0.965 178.82 1.38 ;
      RECT  179.235 0.965 181.68 1.38 ;
      RECT  182.095 0.965 184.54 1.38 ;
      RECT  184.955 0.965 187.4 1.38 ;
      RECT  187.815 0.965 190.26 1.38 ;
      RECT  190.675 0.965 193.12 1.38 ;
      RECT  193.535 0.965 195.98 1.38 ;
      RECT  196.395 0.965 198.84 1.38 ;
      RECT  199.255 0.965 201.7 1.38 ;
      RECT  202.115 0.965 204.56 1.38 ;
      RECT  204.975 0.965 207.42 1.38 ;
      RECT  207.835 0.965 210.28 1.38 ;
      RECT  210.695 0.965 213.14 1.38 ;
      RECT  213.555 0.965 216.0 1.38 ;
      RECT  216.415 0.965 218.86 1.38 ;
      RECT  219.275 0.965 221.72 1.38 ;
      RECT  222.135 0.965 224.58 1.38 ;
      RECT  224.995 0.965 227.44 1.38 ;
      RECT  227.855 0.965 230.3 1.38 ;
      RECT  230.715 0.965 233.16 1.38 ;
      RECT  233.575 0.965 236.02 1.38 ;
      RECT  236.435 0.965 238.88 1.38 ;
      RECT  239.295 0.965 241.74 1.38 ;
      RECT  242.155 0.965 244.6 1.38 ;
      RECT  245.015 0.965 247.46 1.38 ;
      RECT  247.875 0.965 250.32 1.38 ;
      RECT  250.735 0.965 253.18 1.38 ;
      RECT  253.595 0.965 256.04 1.38 ;
      RECT  256.455 0.965 258.9 1.38 ;
      RECT  259.315 0.965 261.76 1.38 ;
      RECT  262.175 0.965 264.62 1.38 ;
      RECT  265.035 0.965 267.48 1.38 ;
      RECT  267.895 0.965 270.34 1.38 ;
      RECT  270.755 0.965 273.2 1.38 ;
      RECT  273.615 0.965 276.06 1.38 ;
      RECT  276.475 0.965 278.92 1.38 ;
      RECT  279.335 0.965 281.78 1.38 ;
      RECT  282.195 0.965 284.64 1.38 ;
      RECT  285.055 0.965 287.5 1.38 ;
      RECT  287.915 0.965 290.36 1.38 ;
      RECT  290.775 0.965 293.22 1.38 ;
      RECT  293.635 0.965 296.08 1.38 ;
      RECT  296.495 0.965 298.94 1.38 ;
      RECT  299.355 0.965 301.8 1.38 ;
      RECT  302.215 0.965 304.66 1.38 ;
      RECT  305.075 0.965 307.52 1.38 ;
      RECT  307.935 0.965 310.38 1.38 ;
      RECT  310.795 0.965 313.24 1.38 ;
      RECT  313.655 0.965 316.1 1.38 ;
      RECT  316.515 0.965 318.96 1.38 ;
      RECT  319.375 0.965 321.82 1.38 ;
      RECT  322.235 0.965 324.68 1.38 ;
      RECT  325.095 0.965 327.54 1.38 ;
      RECT  327.955 0.965 330.4 1.38 ;
      RECT  330.815 0.965 333.26 1.38 ;
      RECT  333.675 0.965 336.12 1.38 ;
      RECT  336.535 0.965 338.98 1.38 ;
      RECT  339.395 0.965 341.84 1.38 ;
      RECT  342.255 0.965 344.7 1.38 ;
      RECT  345.115 0.965 347.56 1.38 ;
      RECT  347.975 0.965 350.42 1.38 ;
      RECT  350.835 0.965 353.28 1.38 ;
      RECT  353.695 0.965 356.14 1.38 ;
      RECT  356.555 0.965 359.0 1.38 ;
      RECT  359.415 0.965 361.86 1.38 ;
      RECT  362.275 0.965 364.72 1.38 ;
      RECT  365.135 0.965 367.58 1.38 ;
      RECT  367.995 0.965 370.44 1.38 ;
      RECT  370.855 0.965 373.3 1.38 ;
      RECT  373.715 0.965 376.16 1.38 ;
      RECT  376.575 0.965 379.02 1.38 ;
      RECT  379.435 0.965 381.88 1.38 ;
      RECT  382.295 0.965 384.74 1.38 ;
      RECT  385.155 0.965 387.6 1.38 ;
      RECT  388.015 0.965 390.46 1.38 ;
      RECT  390.875 0.965 393.32 1.38 ;
      RECT  393.735 0.965 396.18 1.38 ;
      RECT  396.595 0.965 399.04 1.38 ;
      RECT  399.455 0.965 401.9 1.38 ;
      RECT  402.315 0.965 404.76 1.38 ;
      RECT  405.175 0.965 407.62 1.38 ;
      RECT  408.035 0.965 410.48 1.38 ;
      RECT  410.895 0.965 413.34 1.38 ;
      RECT  413.755 0.965 416.2 1.38 ;
      RECT  416.615 0.965 419.06 1.38 ;
      RECT  419.475 0.965 421.92 1.38 ;
      RECT  422.335 0.965 424.78 1.38 ;
      RECT  425.195 0.965 427.64 1.38 ;
      RECT  428.055 0.965 430.5 1.38 ;
      RECT  430.915 0.965 433.36 1.38 ;
      RECT  433.775 0.965 436.22 1.38 ;
      RECT  436.635 0.965 439.08 1.38 ;
      RECT  439.495 0.965 441.94 1.38 ;
      RECT  442.355 0.965 444.8 1.38 ;
      RECT  445.215 0.965 447.66 1.38 ;
      RECT  448.075 0.965 450.52 1.38 ;
      RECT  450.935 0.965 453.38 1.38 ;
      RECT  453.795 0.965 456.24 1.38 ;
      RECT  456.655 0.965 459.1 1.38 ;
      RECT  459.515 0.965 461.96 1.38 ;
      RECT  462.375 0.965 464.82 1.38 ;
      RECT  465.235 0.965 467.68 1.38 ;
      RECT  468.095 0.965 470.54 1.38 ;
      RECT  470.955 0.965 473.4 1.38 ;
      RECT  473.815 0.965 476.26 1.38 ;
      RECT  476.675 0.965 479.12 1.38 ;
      RECT  479.535 0.965 481.98 1.38 ;
      RECT  482.395 0.965 484.84 1.38 ;
      RECT  485.255 0.965 487.7 1.38 ;
      RECT  488.115 0.965 490.56 1.38 ;
      RECT  490.975 0.965 493.42 1.38 ;
      RECT  493.835 0.965 496.28 1.38 ;
      RECT  496.695 0.965 499.14 1.38 ;
      RECT  499.555 0.965 502.0 1.38 ;
      RECT  502.415 0.965 504.86 1.38 ;
      RECT  505.275 0.965 507.72 1.38 ;
      RECT  508.135 0.965 510.58 1.38 ;
      RECT  510.995 0.965 513.44 1.38 ;
      RECT  513.855 0.965 516.3 1.38 ;
      RECT  516.715 0.965 519.16 1.38 ;
      RECT  519.575 0.965 522.02 1.38 ;
      RECT  522.435 0.965 524.88 1.38 ;
      RECT  525.295 0.965 527.74 1.38 ;
      RECT  528.155 0.965 530.6 1.38 ;
      RECT  531.015 0.965 533.46 1.38 ;
      RECT  533.875 0.965 536.32 1.38 ;
      RECT  536.735 0.965 539.18 1.38 ;
      RECT  539.595 0.965 542.04 1.38 ;
      RECT  542.455 0.965 544.9 1.38 ;
      RECT  545.315 0.965 547.76 1.38 ;
      RECT  548.175 0.965 550.62 1.38 ;
      RECT  551.035 0.965 553.48 1.38 ;
      RECT  553.895 0.965 556.34 1.38 ;
      RECT  556.755 0.965 559.2 1.38 ;
      RECT  559.615 0.965 562.06 1.38 ;
      RECT  562.475 0.965 564.92 1.38 ;
      RECT  565.335 0.965 567.78 1.38 ;
      RECT  568.195 0.965 570.64 1.38 ;
      RECT  571.055 0.965 573.5 1.38 ;
      RECT  573.915 0.965 576.36 1.38 ;
      RECT  576.775 0.965 579.005 1.38 ;
      RECT  0.14 80.6425 47.26 81.0575 ;
      RECT  0.14 81.0575 47.26 146.6875 ;
      RECT  47.26 1.38 47.675 80.6425 ;
      RECT  47.675 80.6425 75.86 81.0575 ;
      RECT  47.675 81.0575 75.86 146.6875 ;
      RECT  47.26 81.0575 47.675 83.3725 ;
      RECT  47.26 83.7875 47.675 85.5825 ;
      RECT  47.26 85.9975 47.675 88.3125 ;
      RECT  47.26 88.7275 47.675 90.5225 ;
      RECT  47.26 90.9375 47.675 93.2525 ;
      RECT  47.26 93.6675 47.675 146.6875 ;
      RECT  0.14 1.38 0.145 35.9225 ;
      RECT  0.14 35.9225 0.145 36.3375 ;
      RECT  0.14 36.3375 0.145 80.6425 ;
      RECT  0.145 1.38 0.56 35.9225 ;
      RECT  0.56 1.38 47.26 35.9225 ;
      RECT  0.145 36.3375 0.56 38.6525 ;
      RECT  0.145 39.0675 0.56 80.6425 ;
      RECT  0.56 35.9225 6.3875 36.0075 ;
      RECT  0.56 36.0075 6.3875 36.3375 ;
      RECT  6.3875 35.9225 6.8025 36.0075 ;
      RECT  6.8025 35.9225 47.26 36.0075 ;
      RECT  6.8025 36.0075 47.26 36.3375 ;
      RECT  0.56 36.3375 6.3875 36.4225 ;
      RECT  0.56 36.4225 6.3875 80.6425 ;
      RECT  6.3875 36.4225 6.8025 80.6425 ;
      RECT  6.8025 36.3375 47.26 36.4225 ;
      RECT  6.8025 36.4225 47.26 80.6425 ;
      RECT  0.14 0.965 52.98 1.38 ;
      RECT  53.395 0.965 55.84 1.38 ;
      RECT  56.255 0.965 58.7 1.38 ;
      RECT  59.115 0.965 61.56 1.38 ;
      RECT  61.975 0.965 64.42 1.38 ;
      RECT  64.835 0.965 67.28 1.38 ;
      RECT  67.695 0.965 70.14 1.38 ;
      RECT  70.555 0.965 73.0 1.38 ;
      RECT  73.415 0.965 75.86 1.38 ;
      RECT  47.675 47.5725 72.9725 47.9875 ;
      RECT  73.3875 47.5725 73.6775 47.9875 ;
      RECT  74.0925 47.5725 74.3825 47.9875 ;
      RECT  74.7975 47.5725 75.0875 47.9875 ;
      RECT  76.2075 47.5725 76.275 47.9875 ;
      RECT  75.5025 47.5725 75.7925 47.9875 ;
      RECT  76.275 47.5725 76.4975 47.9875 ;
      RECT  76.9125 47.5725 77.2025 47.9875 ;
      RECT  77.6175 47.5725 77.9075 47.9875 ;
      RECT  78.3225 47.5725 78.6125 47.9875 ;
      RECT  79.0275 47.5725 79.3175 47.9875 ;
      RECT  79.7325 47.5725 80.0225 47.9875 ;
      RECT  80.4375 47.5725 80.7275 47.9875 ;
      RECT  81.1425 47.5725 81.4325 47.9875 ;
      RECT  81.8475 47.5725 82.1375 47.9875 ;
      RECT  82.5525 47.5725 82.8425 47.9875 ;
      RECT  83.2575 47.5725 83.5475 47.9875 ;
      RECT  83.9625 47.5725 84.2525 47.9875 ;
      RECT  84.6675 47.5725 84.9575 47.9875 ;
      RECT  85.3725 47.5725 85.6625 47.9875 ;
      RECT  86.0775 47.5725 86.3675 47.9875 ;
      RECT  86.7825 47.5725 87.0725 47.9875 ;
      RECT  87.4875 47.5725 87.7775 47.9875 ;
      RECT  88.1925 47.5725 88.4825 47.9875 ;
      RECT  88.8975 47.5725 89.1875 47.9875 ;
      RECT  89.6025 47.5725 89.8925 47.9875 ;
      RECT  90.3075 47.5725 90.5975 47.9875 ;
      RECT  91.0125 47.5725 91.3025 47.9875 ;
      RECT  91.7175 47.5725 92.0075 47.9875 ;
      RECT  92.4225 47.5725 92.7125 47.9875 ;
      RECT  93.1275 47.5725 93.4175 47.9875 ;
      RECT  93.8325 47.5725 94.1225 47.9875 ;
      RECT  94.5375 47.5725 94.8275 47.9875 ;
      RECT  95.2425 47.5725 95.5325 47.9875 ;
      RECT  95.9475 47.5725 96.2375 47.9875 ;
      RECT  96.6525 47.5725 96.9425 47.9875 ;
      RECT  97.3575 47.5725 97.6475 47.9875 ;
      RECT  98.0625 47.5725 98.3525 47.9875 ;
      RECT  98.7675 47.5725 99.0575 47.9875 ;
      RECT  99.4725 47.5725 99.7625 47.9875 ;
      RECT  100.1775 47.5725 100.4675 47.9875 ;
      RECT  100.8825 47.5725 101.1725 47.9875 ;
      RECT  101.5875 47.5725 101.8775 47.9875 ;
      RECT  102.2925 47.5725 102.5825 47.9875 ;
      RECT  102.9975 47.5725 103.2875 47.9875 ;
      RECT  103.7025 47.5725 103.9925 47.9875 ;
      RECT  104.4075 47.5725 104.6975 47.9875 ;
      RECT  105.1125 47.5725 105.4025 47.9875 ;
      RECT  105.8175 47.5725 106.1075 47.9875 ;
      RECT  106.5225 47.5725 106.8125 47.9875 ;
      RECT  107.2275 47.5725 107.5175 47.9875 ;
      RECT  107.9325 47.5725 108.2225 47.9875 ;
      RECT  108.6375 47.5725 108.9275 47.9875 ;
      RECT  109.3425 47.5725 109.6325 47.9875 ;
      RECT  110.0475 47.5725 110.3375 47.9875 ;
      RECT  110.7525 47.5725 111.0425 47.9875 ;
      RECT  111.4575 47.5725 111.7475 47.9875 ;
      RECT  112.1625 47.5725 112.4525 47.9875 ;
      RECT  112.8675 47.5725 113.1575 47.9875 ;
      RECT  113.5725 47.5725 113.8625 47.9875 ;
      RECT  114.2775 47.5725 114.5675 47.9875 ;
      RECT  114.9825 47.5725 115.2725 47.9875 ;
      RECT  115.6875 47.5725 115.9775 47.9875 ;
      RECT  116.3925 47.5725 116.6825 47.9875 ;
      RECT  117.0975 47.5725 117.3875 47.9875 ;
      RECT  117.8025 47.5725 118.0925 47.9875 ;
      RECT  118.5075 47.5725 118.7975 47.9875 ;
      RECT  119.2125 47.5725 119.5025 47.9875 ;
      RECT  119.9175 47.5725 120.2075 47.9875 ;
      RECT  120.6225 47.5725 120.9125 47.9875 ;
      RECT  121.3275 47.5725 121.6175 47.9875 ;
      RECT  122.0325 47.5725 122.3225 47.9875 ;
      RECT  122.7375 47.5725 123.0275 47.9875 ;
      RECT  123.4425 47.5725 123.7325 47.9875 ;
      RECT  124.1475 47.5725 124.4375 47.9875 ;
      RECT  124.8525 47.5725 125.1425 47.9875 ;
      RECT  125.5575 47.5725 125.8475 47.9875 ;
      RECT  126.2625 47.5725 126.5525 47.9875 ;
      RECT  126.9675 47.5725 127.2575 47.9875 ;
      RECT  127.6725 47.5725 127.9625 47.9875 ;
      RECT  128.3775 47.5725 128.6675 47.9875 ;
      RECT  129.0825 47.5725 129.3725 47.9875 ;
      RECT  129.7875 47.5725 130.0775 47.9875 ;
      RECT  130.4925 47.5725 130.7825 47.9875 ;
      RECT  131.1975 47.5725 131.4875 47.9875 ;
      RECT  131.9025 47.5725 132.1925 47.9875 ;
      RECT  132.6075 47.5725 132.8975 47.9875 ;
      RECT  133.3125 47.5725 133.6025 47.9875 ;
      RECT  134.0175 47.5725 134.3075 47.9875 ;
      RECT  134.7225 47.5725 135.0125 47.9875 ;
      RECT  135.4275 47.5725 135.7175 47.9875 ;
      RECT  136.1325 47.5725 136.4225 47.9875 ;
      RECT  136.8375 47.5725 137.1275 47.9875 ;
      RECT  137.5425 47.5725 137.8325 47.9875 ;
      RECT  138.2475 47.5725 138.5375 47.9875 ;
      RECT  138.9525 47.5725 139.2425 47.9875 ;
      RECT  139.6575 47.5725 139.9475 47.9875 ;
      RECT  140.3625 47.5725 140.6525 47.9875 ;
      RECT  141.0675 47.5725 141.3575 47.9875 ;
      RECT  141.7725 47.5725 142.0625 47.9875 ;
      RECT  142.4775 47.5725 142.7675 47.9875 ;
      RECT  143.1825 47.5725 143.4725 47.9875 ;
      RECT  143.8875 47.5725 144.1775 47.9875 ;
      RECT  144.5925 47.5725 144.8825 47.9875 ;
      RECT  145.2975 47.5725 145.5875 47.9875 ;
      RECT  146.0025 47.5725 146.2925 47.9875 ;
      RECT  146.7075 47.5725 146.9975 47.9875 ;
      RECT  147.4125 47.5725 147.7025 47.9875 ;
      RECT  148.1175 47.5725 148.4075 47.9875 ;
      RECT  148.8225 47.5725 149.1125 47.9875 ;
      RECT  149.5275 47.5725 149.8175 47.9875 ;
      RECT  150.2325 47.5725 150.5225 47.9875 ;
      RECT  150.9375 47.5725 151.2275 47.9875 ;
      RECT  151.6425 47.5725 151.9325 47.9875 ;
      RECT  152.3475 47.5725 152.6375 47.9875 ;
      RECT  153.0525 47.5725 153.3425 47.9875 ;
      RECT  153.7575 47.5725 154.0475 47.9875 ;
      RECT  154.4625 47.5725 154.7525 47.9875 ;
      RECT  155.1675 47.5725 155.4575 47.9875 ;
      RECT  155.8725 47.5725 156.1625 47.9875 ;
      RECT  156.5775 47.5725 156.8675 47.9875 ;
      RECT  157.2825 47.5725 157.5725 47.9875 ;
      RECT  157.9875 47.5725 158.2775 47.9875 ;
      RECT  158.6925 47.5725 158.9825 47.9875 ;
      RECT  159.3975 47.5725 159.6875 47.9875 ;
      RECT  160.1025 47.5725 160.3925 47.9875 ;
      RECT  160.8075 47.5725 161.0975 47.9875 ;
      RECT  161.5125 47.5725 161.8025 47.9875 ;
      RECT  162.2175 47.5725 162.5075 47.9875 ;
      RECT  162.9225 47.5725 163.2125 47.9875 ;
      RECT  163.6275 47.5725 163.9175 47.9875 ;
      RECT  164.3325 47.5725 164.6225 47.9875 ;
      RECT  165.0375 47.5725 165.3275 47.9875 ;
      RECT  165.7425 47.5725 166.0325 47.9875 ;
      RECT  166.4475 47.5725 166.7375 47.9875 ;
      RECT  167.1525 47.5725 167.4425 47.9875 ;
      RECT  167.8575 47.5725 168.1475 47.9875 ;
      RECT  168.5625 47.5725 168.8525 47.9875 ;
      RECT  169.2675 47.5725 169.5575 47.9875 ;
      RECT  169.9725 47.5725 170.2625 47.9875 ;
      RECT  170.6775 47.5725 170.9675 47.9875 ;
      RECT  171.3825 47.5725 171.6725 47.9875 ;
      RECT  172.0875 47.5725 172.3775 47.9875 ;
      RECT  172.7925 47.5725 173.0825 47.9875 ;
      RECT  173.4975 47.5725 173.7875 47.9875 ;
      RECT  174.2025 47.5725 174.4925 47.9875 ;
      RECT  174.9075 47.5725 175.1975 47.9875 ;
      RECT  175.6125 47.5725 175.9025 47.9875 ;
      RECT  176.3175 47.5725 176.6075 47.9875 ;
      RECT  177.0225 47.5725 177.3125 47.9875 ;
      RECT  177.7275 47.5725 178.0175 47.9875 ;
      RECT  178.4325 47.5725 178.7225 47.9875 ;
      RECT  179.1375 47.5725 179.4275 47.9875 ;
      RECT  179.8425 47.5725 180.1325 47.9875 ;
      RECT  180.5475 47.5725 180.8375 47.9875 ;
      RECT  181.2525 47.5725 181.5425 47.9875 ;
      RECT  181.9575 47.5725 182.2475 47.9875 ;
      RECT  182.6625 47.5725 182.9525 47.9875 ;
      RECT  183.3675 47.5725 183.6575 47.9875 ;
      RECT  184.0725 47.5725 184.3625 47.9875 ;
      RECT  184.7775 47.5725 185.0675 47.9875 ;
      RECT  185.4825 47.5725 185.7725 47.9875 ;
      RECT  186.1875 47.5725 186.4775 47.9875 ;
      RECT  186.8925 47.5725 187.1825 47.9875 ;
      RECT  187.5975 47.5725 187.8875 47.9875 ;
      RECT  188.3025 47.5725 188.5925 47.9875 ;
      RECT  189.0075 47.5725 189.2975 47.9875 ;
      RECT  189.7125 47.5725 190.0025 47.9875 ;
      RECT  190.4175 47.5725 190.7075 47.9875 ;
      RECT  191.1225 47.5725 191.4125 47.9875 ;
      RECT  191.8275 47.5725 192.1175 47.9875 ;
      RECT  192.5325 47.5725 192.8225 47.9875 ;
      RECT  193.2375 47.5725 193.5275 47.9875 ;
      RECT  193.9425 47.5725 194.2325 47.9875 ;
      RECT  194.6475 47.5725 194.9375 47.9875 ;
      RECT  195.3525 47.5725 195.6425 47.9875 ;
      RECT  196.0575 47.5725 196.3475 47.9875 ;
      RECT  196.7625 47.5725 579.005 47.9875 ;
      RECT  47.675 67.2525 53.0775 67.6675 ;
      RECT  53.4925 67.2525 72.9725 67.6675 ;
      RECT  53.4925 67.6675 72.9725 80.6425 ;
      RECT  76.9125 1.38 418.7775 2.33 ;
      RECT  418.7775 1.38 419.1925 2.33 ;
      RECT  418.7775 2.745 419.1925 47.5725 ;
      RECT  419.1925 1.38 579.005 2.33 ;
      RECT  419.1925 2.745 579.005 47.5725 ;
      RECT  73.3875 1.38 75.5775 2.33 ;
      RECT  73.3875 2.33 75.5775 2.745 ;
      RECT  75.5775 1.38 75.86 2.33 ;
      RECT  75.86 1.38 75.9925 2.33 ;
      RECT  75.9925 1.38 76.2075 2.33 ;
      RECT  75.9925 2.33 76.2075 2.745 ;
      RECT  53.0775 47.9875 53.4925 59.0625 ;
      RECT  72.9725 47.9875 73.3875 50.1925 ;
      RECT  73.3875 47.9875 75.86 50.1925 ;
      RECT  75.86 47.9875 76.2075 50.1925 ;
      RECT  76.2075 47.9875 76.275 50.1925 ;
      RECT  76.275 47.9875 76.4975 50.1925 ;
      RECT  76.4975 47.9875 76.9125 50.1925 ;
      RECT  76.9125 47.9875 197.4325 50.1925 ;
      RECT  197.4325 47.9875 579.005 50.1925 ;
      RECT  197.4325 50.1925 579.005 50.5425 ;
      RECT  53.4925 47.9875 70.7275 50.1925 ;
      RECT  53.4925 50.1925 70.7275 50.5425 ;
      RECT  70.7275 47.9875 72.9725 50.1925 ;
      RECT  53.0775 59.4775 53.4925 61.7925 ;
      RECT  53.0775 62.2075 53.4925 67.2525 ;
      RECT  407.7525 2.33 418.7775 2.745 ;
      RECT  47.675 1.38 52.6975 2.33 ;
      RECT  47.675 2.33 52.6975 2.745 ;
      RECT  47.675 2.745 52.6975 47.5725 ;
      RECT  52.6975 1.38 53.1125 2.33 ;
      RECT  52.6975 2.745 53.1125 47.5725 ;
      RECT  53.1125 1.38 72.9725 2.33 ;
      RECT  247.5925 2.33 258.6175 2.745 ;
      RECT  53.4925 50.5425 69.5825 56.3325 ;
      RECT  53.4925 56.3325 69.5825 56.7475 ;
      RECT  69.5825 50.5425 69.9975 56.3325 ;
      RECT  69.5825 56.7475 69.9975 67.2525 ;
      RECT  69.9975 50.5425 70.7275 56.3325 ;
      RECT  69.9975 56.3325 70.7275 56.7475 ;
      RECT  69.9975 56.7475 70.7275 67.2525 ;
      RECT  339.1125 2.33 350.1375 2.745 ;
      RECT  316.2325 2.33 327.2575 2.745 ;
      RECT  327.6725 2.33 338.6975 2.745 ;
      RECT  304.7925 2.33 315.8175 2.745 ;
      RECT  293.3525 2.33 304.3775 2.745 ;
      RECT  281.9125 2.33 292.9375 2.745 ;
      RECT  213.2725 2.33 224.2975 2.745 ;
      RECT  76.9125 2.33 87.0175 2.745 ;
      RECT  201.8325 2.33 212.8575 2.745 ;
      RECT  442.0725 2.33 453.0975 2.745 ;
      RECT  72.9725 1.38 73.3875 43.265 ;
      RECT  76.2075 1.38 76.275 43.265 ;
      RECT  76.275 1.38 76.4975 43.265 ;
      RECT  76.4975 1.38 76.9125 43.265 ;
      RECT  197.4325 2.745 418.7775 43.265 ;
      RECT  197.4325 43.265 418.7775 43.615 ;
      RECT  197.4325 43.615 418.7775 47.5725 ;
      RECT  73.3875 2.745 75.5775 43.265 ;
      RECT  75.5775 2.745 75.86 43.265 ;
      RECT  75.86 2.745 75.9925 43.265 ;
      RECT  75.9925 2.745 76.2075 43.265 ;
      RECT  53.1125 43.265 70.7275 43.615 ;
      RECT  53.1125 43.615 70.7275 47.5725 ;
      RECT  259.0325 2.33 270.0575 2.745 ;
      RECT  270.4725 2.33 281.4975 2.745 ;
      RECT  87.4325 2.33 98.4575 2.745 ;
      RECT  98.8725 2.33 109.8975 2.745 ;
      RECT  567.9125 2.33 579.005 2.745 ;
      RECT  53.1125 2.745 70.5925 42.2975 ;
      RECT  53.1125 42.2975 70.5925 42.7125 ;
      RECT  53.1125 42.7125 70.5925 43.265 ;
      RECT  70.5925 42.7125 70.7275 43.265 ;
      RECT  70.7275 42.7125 71.0075 43.265 ;
      RECT  71.0075 2.745 72.9725 42.2975 ;
      RECT  71.0075 42.2975 72.9725 42.7125 ;
      RECT  71.0075 42.7125 72.9725 43.265 ;
      RECT  224.7125 2.33 235.7375 2.745 ;
      RECT  236.1525 2.33 247.1775 2.745 ;
      RECT  522.1525 2.33 533.1775 2.745 ;
      RECT  533.5925 2.33 544.6175 2.745 ;
      RECT  545.0325 2.33 556.0575 2.745 ;
      RECT  556.4725 2.33 567.4975 2.745 ;
      RECT  373.4325 2.33 384.4575 2.745 ;
      RECT  156.0725 2.33 167.0975 2.745 ;
      RECT  384.8725 2.33 395.8975 2.745 ;
      RECT  396.3125 2.33 407.3375 2.745 ;
      RECT  72.9725 54.44 73.3875 80.6425 ;
      RECT  73.3875 54.44 75.86 80.6425 ;
      RECT  75.86 54.44 76.2075 146.6875 ;
      RECT  76.2075 54.44 76.275 146.6875 ;
      RECT  76.275 54.44 76.4975 146.6875 ;
      RECT  76.4975 54.44 76.9125 146.6875 ;
      RECT  76.9125 54.44 197.4325 146.6875 ;
      RECT  70.7275 54.44 72.9725 67.2525 ;
      RECT  487.8325 2.33 498.8575 2.745 ;
      RECT  499.2725 2.33 510.2975 2.745 ;
      RECT  510.7125 2.33 521.7375 2.745 ;
      RECT  453.5125 2.33 464.5375 2.745 ;
      RECT  190.3925 2.33 201.4175 2.745 ;
      RECT  133.1925 2.33 144.2175 2.745 ;
      RECT  144.6325 2.33 155.6575 2.745 ;
      RECT  350.5525 2.33 361.5775 2.745 ;
      RECT  361.9925 2.33 373.0175 2.745 ;
      RECT  53.1125 2.33 64.1375 2.745 ;
      RECT  64.5525 2.33 72.9725 2.745 ;
      RECT  110.3125 2.33 121.3375 2.745 ;
      RECT  121.7525 2.33 132.7775 2.745 ;
      RECT  53.0775 67.6675 53.4925 69.9825 ;
      RECT  53.0775 70.3975 53.4925 75.4425 ;
      RECT  419.1925 2.33 430.2175 2.745 ;
      RECT  430.6325 2.33 441.6575 2.745 ;
      RECT  167.5125 2.33 178.5375 2.745 ;
      RECT  178.9525 2.33 189.9775 2.745 ;
      RECT  53.0775 75.8575 53.4925 78.1725 ;
      RECT  53.0775 78.5875 53.4925 80.6425 ;
      RECT  53.4925 56.7475 59.25 56.99 ;
      RECT  53.4925 56.99 59.25 57.405 ;
      RECT  53.4925 57.405 59.25 67.2525 ;
      RECT  59.25 56.7475 59.665 56.99 ;
      RECT  59.25 57.405 59.665 67.2525 ;
      RECT  59.665 56.7475 69.5825 56.99 ;
      RECT  59.665 56.99 69.5825 57.405 ;
      RECT  59.665 57.405 69.5825 67.2525 ;
      RECT  464.9525 2.33 475.9775 2.745 ;
      RECT  476.3925 2.33 487.4175 2.745 ;
      RECT  76.9125 2.745 197.0175 42.2975 ;
      RECT  76.9125 42.2975 197.0175 42.7125 ;
      RECT  76.9125 42.7125 197.0175 43.265 ;
      RECT  197.0175 42.7125 197.4325 43.265 ;
      RECT  76.275 0.275 147.0775 0.965 ;
      RECT  147.0775 0.275 147.4925 0.965 ;
      RECT  147.4925 0.275 579.005 0.965 ;
      RECT  147.4925 0.14 158.5175 0.275 ;
      RECT  158.9325 0.14 169.9575 0.275 ;
      RECT  387.7325 0.14 398.7575 0.275 ;
      RECT  47.675 67.6675 51.55 71.3475 ;
      RECT  47.675 71.3475 51.55 71.7625 ;
      RECT  47.675 71.7625 51.55 80.6425 ;
      RECT  51.965 67.6675 53.0775 71.3475 ;
      RECT  51.965 71.3475 53.0775 71.7625 ;
      RECT  51.965 71.7625 53.0775 80.6425 ;
      RECT  51.55 71.7625 51.965 74.0775 ;
      RECT  51.55 67.6675 51.965 68.6175 ;
      RECT  51.55 69.0325 51.965 71.3475 ;
      RECT  239.0125 0.14 250.0375 0.275 ;
      RECT  90.2925 0.14 101.3175 0.275 ;
      RECT  197.0175 2.745 197.4325 40.4775 ;
      RECT  197.0175 40.8925 197.4325 42.2975 ;
      RECT  0.14 0.14 55.5575 0.275 ;
      RECT  0.14 0.275 55.5575 0.965 ;
      RECT  55.5575 0.275 55.9725 0.965 ;
      RECT  55.9725 0.275 75.86 0.965 ;
      RECT  55.9725 0.14 66.9975 0.275 ;
      RECT  67.4125 0.14 75.86 0.275 ;
      RECT  422.0525 0.14 433.0775 0.275 ;
      RECT  170.3725 0.14 181.3975 0.275 ;
      RECT  47.675 47.9875 51.55 63.1575 ;
      RECT  47.675 63.1575 51.55 63.5725 ;
      RECT  47.675 63.5725 51.55 67.2525 ;
      RECT  51.965 47.9875 53.0775 63.1575 ;
      RECT  51.965 63.1575 53.0775 63.5725 ;
      RECT  51.965 63.5725 53.0775 67.2525 ;
      RECT  51.55 79.9525 51.965 80.6425 ;
      RECT  536.4525 0.14 547.4775 0.275 ;
      RECT  547.8925 0.14 558.9175 0.275 ;
      RECT  101.7325 0.14 112.7575 0.275 ;
      RECT  136.0525 0.14 147.0775 0.275 ;
      RECT  376.2925 0.14 387.3175 0.275 ;
      RECT  181.8125 0.14 192.8375 0.275 ;
      RECT  51.55 60.8425 51.965 63.1575 ;
      RECT  197.4325 50.5425 197.4675 52.085 ;
      RECT  197.4325 52.435 197.4675 146.6875 ;
      RECT  197.4675 50.5425 579.005 52.085 ;
      RECT  197.4675 52.085 579.005 52.435 ;
      RECT  197.4675 52.435 579.005 146.6875 ;
      RECT  72.9725 50.5425 73.3875 52.085 ;
      RECT  72.9725 52.435 73.3875 54.09 ;
      RECT  73.3875 50.5425 75.86 52.085 ;
      RECT  73.3875 52.435 75.86 54.09 ;
      RECT  75.86 50.5425 76.2075 52.085 ;
      RECT  75.86 52.435 76.2075 54.09 ;
      RECT  76.2075 50.5425 76.275 52.085 ;
      RECT  76.2075 52.435 76.275 54.09 ;
      RECT  76.275 50.5425 76.4975 52.085 ;
      RECT  76.275 52.435 76.4975 54.09 ;
      RECT  76.4975 50.5425 76.9125 52.085 ;
      RECT  76.4975 52.435 76.9125 54.09 ;
      RECT  76.9125 50.5425 197.4325 52.085 ;
      RECT  76.9125 52.435 197.4325 54.09 ;
      RECT  70.7275 50.5425 72.9725 52.085 ;
      RECT  70.7275 52.435 72.9725 54.09 ;
      RECT  479.2525 0.14 490.2775 0.275 ;
      RECT  51.55 74.4925 51.965 76.8075 ;
      RECT  51.55 77.2225 51.965 79.5375 ;
      RECT  72.9725 43.615 73.3875 45.315 ;
      RECT  72.9725 45.665 73.3875 47.5725 ;
      RECT  76.2075 43.615 76.275 45.315 ;
      RECT  76.2075 45.665 76.275 47.5725 ;
      RECT  76.275 43.615 76.4975 45.315 ;
      RECT  76.275 45.665 76.4975 47.5725 ;
      RECT  76.4975 43.615 76.9125 45.315 ;
      RECT  76.4975 45.665 76.9125 47.5725 ;
      RECT  76.9125 43.615 197.4325 45.315 ;
      RECT  76.9125 45.665 197.4325 47.5725 ;
      RECT  73.3875 43.615 75.5775 45.315 ;
      RECT  73.3875 45.665 75.5775 47.5725 ;
      RECT  75.5775 43.615 75.86 45.315 ;
      RECT  75.5775 45.665 75.86 47.5725 ;
      RECT  75.86 43.615 75.9925 45.315 ;
      RECT  75.86 45.665 75.9925 47.5725 ;
      RECT  75.9925 43.615 76.2075 45.315 ;
      RECT  75.9925 45.665 76.2075 47.5725 ;
      RECT  70.7275 43.615 72.9725 45.315 ;
      RECT  70.7275 45.665 72.9725 47.5725 ;
      RECT  330.5325 0.14 341.5575 0.275 ;
      RECT  456.3725 0.14 467.3975 0.275 ;
      RECT  467.8125 0.14 478.8375 0.275 ;
      RECT  273.3325 0.14 284.3575 0.275 ;
      RECT  76.275 0.14 78.4375 0.275 ;
      RECT  78.8525 0.14 89.8775 0.275 ;
      RECT  490.6925 0.14 501.7175 0.275 ;
      RECT  341.9725 0.14 352.9975 0.275 ;
      RECT  502.1325 0.14 513.1575 0.275 ;
      RECT  399.1725 0.14 410.1975 0.275 ;
      RECT  410.6125 0.14 421.6375 0.275 ;
      RECT  353.4125 0.14 364.4375 0.275 ;
      RECT  364.8525 0.14 375.8775 0.275 ;
      RECT  193.2525 0.14 204.2775 0.275 ;
      RECT  204.6925 0.14 215.7175 0.275 ;
      RECT  51.55 63.5725 51.965 65.8875 ;
      RECT  51.55 66.3025 51.965 67.2525 ;
      RECT  513.5725 0.14 524.5975 0.275 ;
      RECT  525.0125 0.14 536.0375 0.275 ;
      RECT  284.7725 0.14 295.7975 0.275 ;
      RECT  433.4925 0.14 444.5175 0.275 ;
      RECT  444.9325 0.14 455.9575 0.275 ;
      RECT  113.1725 0.14 124.1975 0.275 ;
      RECT  124.6125 0.14 135.6375 0.275 ;
      RECT  296.2125 0.14 307.2375 0.275 ;
      RECT  70.5925 2.745 70.7275 40.4775 ;
      RECT  70.5925 40.8925 70.7275 42.2975 ;
      RECT  70.7275 2.745 71.0075 40.4775 ;
      RECT  70.7275 40.8925 71.0075 42.2975 ;
      RECT  307.6525 0.14 318.6775 0.275 ;
      RECT  319.0925 0.14 330.1175 0.275 ;
      RECT  51.55 47.9875 51.965 57.6975 ;
      RECT  51.55 58.1125 51.965 60.4275 ;
      RECT  216.1325 0.14 227.1575 0.275 ;
      RECT  227.5725 0.14 238.5975 0.275 ;
      RECT  559.3325 0.14 570.3575 0.275 ;
      RECT  570.7725 0.14 579.005 0.275 ;
      RECT  250.4525 0.14 261.4775 0.275 ;
      RECT  261.8925 0.14 272.9175 0.275 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 0.42 34.675 ;
      RECT  0.14 40.315 0.4075 44.5225 ;
      RECT  0.14 44.5225 0.4075 67.485 ;
      RECT  0.14 67.485 0.4075 146.6875 ;
      RECT  0.4075 40.315 0.42 44.5225 ;
      RECT  0.4075 67.485 0.42 146.6875 ;
      RECT  0.42 40.315 1.1075 44.5225 ;
      RECT  0.42 67.485 1.1075 146.6875 ;
      RECT  1.1075 145.685 58.49 146.6875 ;
      RECT  58.49 145.685 59.19 146.6875 ;
      RECT  59.19 44.5225 70.52 54.645 ;
      RECT  70.52 44.5225 71.22 54.645 ;
      RECT  71.22 44.5225 579.005 54.645 ;
      RECT  59.19 145.685 70.52 146.6875 ;
      RECT  70.14 57.555 70.52 67.485 ;
      RECT  69.44 145.615 70.14 145.685 ;
      RECT  70.14 67.485 70.52 145.615 ;
      RECT  70.14 145.615 70.52 145.685 ;
      RECT  49.555 34.675 50.255 37.145 ;
      RECT  50.255 34.675 579.005 37.145 ;
      RECT  50.255 37.145 579.005 40.315 ;
      RECT  50.255 40.315 579.005 44.5225 ;
      RECT  49.555 52.665 50.255 57.555 ;
      RECT  50.255 44.5225 58.49 52.665 ;
      RECT  1.1075 79.395 46.835 94.915 ;
      RECT  1.1075 94.915 46.835 145.685 ;
      RECT  46.835 67.485 47.535 79.395 ;
      RECT  46.835 94.915 47.535 145.685 ;
      RECT  199.145 54.645 579.005 57.555 ;
      RECT  199.145 57.555 579.005 67.485 ;
      RECT  199.145 67.485 579.005 145.685 ;
      RECT  199.145 145.685 579.005 146.6875 ;
      RECT  0.42 0.14 4.565 34.61 ;
      RECT  0.42 34.61 4.565 34.675 ;
      RECT  4.565 0.14 5.265 34.61 ;
      RECT  5.265 0.14 579.005 34.61 ;
      RECT  5.265 34.61 579.005 34.675 ;
      RECT  0.42 34.675 4.565 37.145 ;
      RECT  0.42 37.145 4.565 40.315 ;
      RECT  1.1075 40.315 4.565 40.38 ;
      RECT  1.1075 40.38 4.565 44.5225 ;
      RECT  4.565 40.38 5.265 44.5225 ;
      RECT  58.49 44.5225 59.05 57.5225 ;
      RECT  58.49 57.5225 59.05 57.555 ;
      RECT  59.05 44.5225 59.19 57.5225 ;
      RECT  59.19 54.645 59.75 57.5225 ;
      RECT  59.75 54.645 70.52 57.5225 ;
      RECT  59.75 57.5225 70.52 57.555 ;
      RECT  59.75 57.555 69.44 67.485 ;
      RECT  59.75 67.485 69.44 145.615 ;
      RECT  59.19 145.6475 59.75 145.685 ;
      RECT  59.75 145.615 69.44 145.6475 ;
      RECT  59.75 145.6475 69.44 145.685 ;
      RECT  47.535 67.485 49.695 79.33 ;
      RECT  47.535 79.33 49.695 79.395 ;
      RECT  49.695 67.485 50.395 79.33 ;
      RECT  47.535 79.395 49.695 94.915 ;
      RECT  47.535 94.915 49.695 94.98 ;
      RECT  47.535 94.98 49.695 145.685 ;
      RECT  49.695 94.98 50.395 145.685 ;
      RECT  6.805 44.5225 49.555 52.665 ;
      RECT  6.105 55.135 6.805 57.555 ;
      RECT  6.805 52.665 49.555 55.135 ;
      RECT  6.805 55.135 49.555 57.555 ;
      RECT  5.265 34.675 6.105 37.145 ;
      RECT  6.805 34.675 49.555 37.145 ;
      RECT  5.265 37.145 6.105 40.315 ;
      RECT  6.805 37.145 49.555 40.315 ;
      RECT  5.265 40.315 6.105 40.38 ;
      RECT  6.805 40.315 49.555 40.38 ;
      RECT  5.265 40.38 6.105 44.5225 ;
      RECT  6.805 40.38 49.555 44.5225 ;
      RECT  57.255 57.555 58.49 67.485 ;
      RECT  50.255 52.665 56.555 57.5225 ;
      RECT  50.255 57.5225 56.555 57.555 ;
      RECT  56.555 52.665 57.255 57.5225 ;
      RECT  57.255 52.665 58.49 57.5225 ;
      RECT  57.255 57.5225 58.49 57.555 ;
      RECT  50.395 67.485 56.555 79.33 ;
      RECT  57.255 67.485 58.49 79.33 ;
      RECT  50.395 79.33 56.555 79.395 ;
      RECT  57.255 79.33 58.49 79.395 ;
      RECT  50.395 79.395 56.555 94.915 ;
      RECT  57.255 79.395 58.49 94.915 ;
      RECT  50.395 94.915 56.555 94.98 ;
      RECT  57.255 94.915 58.49 94.98 ;
      RECT  50.395 94.98 56.555 145.685 ;
      RECT  57.255 94.98 58.49 145.685 ;
      RECT  71.68 54.645 197.985 57.555 ;
      RECT  71.68 57.555 197.985 67.485 ;
      RECT  71.68 67.485 197.985 145.685 ;
      RECT  71.68 145.685 197.985 146.6875 ;
      RECT  1.1075 67.485 2.47 67.5175 ;
      RECT  1.1075 67.5175 2.47 79.395 ;
      RECT  2.47 67.5175 3.17 79.395 ;
      RECT  3.17 67.485 46.835 67.5175 ;
      RECT  3.17 67.5175 46.835 79.395 ;
      RECT  1.1075 44.5225 2.47 44.555 ;
      RECT  1.1075 44.555 2.47 52.665 ;
      RECT  2.47 44.5225 3.17 44.555 ;
      RECT  3.17 44.5225 6.105 44.555 ;
      RECT  3.17 44.555 6.105 52.665 ;
      RECT  1.1075 52.665 2.47 55.135 ;
      RECT  3.17 52.665 6.105 55.135 ;
      RECT  1.1075 55.135 2.47 57.555 ;
      RECT  3.17 55.135 6.105 57.555 ;
      RECT  1.1075 57.555 2.47 67.485 ;
      RECT  3.17 57.555 56.555 67.485 ;
   END
END    freepdk45_sram_1rw0r_64x176_22
END    LIBRARY
