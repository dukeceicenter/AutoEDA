../macros/freepdk45_sram_1w1r_48x32_32/freepdk45_sram_1w1r_48x32_32.lef