../macros/freepdk45_sram_1w1r_128x4_1/freepdk45_sram_1w1r_128x4_1.lef