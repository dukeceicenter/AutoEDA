VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_128x124_31
   CLASS BLOCK ;
   SIZE 407.98 BY 244.585 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.555 1.105 53.69 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.415 1.105 56.55 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.275 1.105 59.41 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.135 1.105 62.27 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.995 1.105 65.13 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.855 1.105 67.99 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.715 1.105 70.85 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.575 1.105 73.71 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.435 1.105 76.57 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.295 1.105 79.43 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.155 1.105 82.29 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.015 1.105 85.15 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.875 1.105 88.01 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.735 1.105 90.87 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.595 1.105 93.73 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.455 1.105 96.59 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.315 1.105 99.45 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.175 1.105 102.31 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.035 1.105 105.17 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.895 1.105 108.03 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.755 1.105 110.89 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.615 1.105 113.75 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.475 1.105 116.61 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.335 1.105 119.47 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.195 1.105 122.33 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.055 1.105 125.19 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.915 1.105 128.05 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.775 1.105 130.91 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.635 1.105 133.77 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.495 1.105 136.63 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.355 1.105 139.49 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.215 1.105 142.35 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.075 1.105 145.21 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.935 1.105 148.07 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.795 1.105 150.93 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.655 1.105 153.79 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.515 1.105 156.65 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.375 1.105 159.51 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.235 1.105 162.37 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.095 1.105 165.23 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.955 1.105 168.09 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.815 1.105 170.95 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.675 1.105 173.81 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.535 1.105 176.67 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.395 1.105 179.53 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.255 1.105 182.39 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.115 1.105 185.25 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.975 1.105 188.11 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.835 1.105 190.97 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.695 1.105 193.83 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.555 1.105 196.69 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.415 1.105 199.55 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.275 1.105 202.41 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.135 1.105 205.27 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.995 1.105 208.13 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.855 1.105 210.99 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.715 1.105 213.85 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.575 1.105 216.71 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.435 1.105 219.57 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.295 1.105 222.43 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.155 1.105 225.29 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.015 1.105 228.15 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.875 1.105 231.01 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.735 1.105 233.87 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.595 1.105 236.73 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.455 1.105 239.59 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.315 1.105 242.45 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.175 1.105 245.31 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.035 1.105 248.17 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.895 1.105 251.03 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.755 1.105 253.89 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.615 1.105 256.75 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.475 1.105 259.61 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.335 1.105 262.47 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.195 1.105 265.33 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.055 1.105 268.19 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.915 1.105 271.05 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.775 1.105 273.91 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.635 1.105 276.77 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.495 1.105 279.63 1.24 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  282.355 1.105 282.49 1.24 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.215 1.105 285.35 1.24 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.075 1.105 288.21 1.24 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.935 1.105 291.07 1.24 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.795 1.105 293.93 1.24 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.655 1.105 296.79 1.24 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.515 1.105 299.65 1.24 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  302.375 1.105 302.51 1.24 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.235 1.105 305.37 1.24 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.095 1.105 308.23 1.24 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.955 1.105 311.09 1.24 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.815 1.105 313.95 1.24 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.675 1.105 316.81 1.24 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.535 1.105 319.67 1.24 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  322.395 1.105 322.53 1.24 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.255 1.105 325.39 1.24 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.115 1.105 328.25 1.24 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.975 1.105 331.11 1.24 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.835 1.105 333.97 1.24 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.695 1.105 336.83 1.24 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.555 1.105 339.69 1.24 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.415 1.105 342.55 1.24 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.275 1.105 345.41 1.24 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.135 1.105 348.27 1.24 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.995 1.105 351.13 1.24 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.855 1.105 353.99 1.24 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.715 1.105 356.85 1.24 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.575 1.105 359.71 1.24 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.435 1.105 362.57 1.24 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.295 1.105 365.43 1.24 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.155 1.105 368.29 1.24 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  371.015 1.105 371.15 1.24 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.875 1.105 374.01 1.24 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  376.735 1.105 376.87 1.24 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  379.595 1.105 379.73 1.24 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  382.455 1.105 382.59 1.24 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  385.315 1.105 385.45 1.24 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  388.175 1.105 388.31 1.24 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  391.035 1.105 391.17 1.24 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.895 1.105 394.03 1.24 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.755 1.105 396.89 1.24 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.615 1.105 399.75 1.24 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  402.475 1.105 402.61 1.24 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  405.335 1.105 405.47 1.24 ;
      END
   END din0[123]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.395 66.0725 36.53 66.2075 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.395 68.8025 36.53 68.9375 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.395 71.0125 36.53 71.1475 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.395 73.7425 36.53 73.8775 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.395 75.9525 36.53 76.0875 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.395 78.6825 36.53 78.8175 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.395 80.8925 36.53 81.0275 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.305 33.9625 231.44 34.0975 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.305 31.2325 231.44 31.3675 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.305 29.0225 231.44 29.1575 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.305 26.2925 231.44 26.4275 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.305 24.0825 231.44 24.2175 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.305 21.3525 231.44 21.4875 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.305 19.1425 231.44 19.2775 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 15.5025 0.42 15.6375 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.555 243.3425 267.69 243.4775 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 15.5875 6.3825 15.7225 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.4525 243.2575 261.5875 243.3925 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.115 1.105 42.25 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.975 1.105 45.11 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.835 1.105 47.97 1.24 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.695 1.105 50.83 1.24 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.9375 236.6325 61.0725 236.7675 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.1125 236.6325 62.2475 236.7675 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.2875 236.6325 63.4225 236.7675 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.4625 236.6325 64.5975 236.7675 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.6375 236.6325 65.7725 236.7675 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.8125 236.6325 66.9475 236.7675 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.9875 236.6325 68.1225 236.7675 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.1625 236.6325 69.2975 236.7675 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.3375 236.6325 70.4725 236.7675 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.5125 236.6325 71.6475 236.7675 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.6875 236.6325 72.8225 236.7675 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.8625 236.6325 73.9975 236.7675 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.0375 236.6325 75.1725 236.7675 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.2125 236.6325 76.3475 236.7675 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.3875 236.6325 77.5225 236.7675 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.5625 236.6325 78.6975 236.7675 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.7375 236.6325 79.8725 236.7675 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.9125 236.6325 81.0475 236.7675 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.0875 236.6325 82.2225 236.7675 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.2625 236.6325 83.3975 236.7675 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.4375 236.6325 84.5725 236.7675 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.6125 236.6325 85.7475 236.7675 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.7875 236.6325 86.9225 236.7675 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.9625 236.6325 88.0975 236.7675 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.1375 236.6325 89.2725 236.7675 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.3125 236.6325 90.4475 236.7675 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.4875 236.6325 91.6225 236.7675 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.6625 236.6325 92.7975 236.7675 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.8375 236.6325 93.9725 236.7675 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.0125 236.6325 95.1475 236.7675 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.1875 236.6325 96.3225 236.7675 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.3625 236.6325 97.4975 236.7675 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.5375 236.6325 98.6725 236.7675 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.7125 236.6325 99.8475 236.7675 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.8875 236.6325 101.0225 236.7675 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.0625 236.6325 102.1975 236.7675 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.2375 236.6325 103.3725 236.7675 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.4125 236.6325 104.5475 236.7675 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.5875 236.6325 105.7225 236.7675 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.7625 236.6325 106.8975 236.7675 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.9375 236.6325 108.0725 236.7675 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.1125 236.6325 109.2475 236.7675 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.2875 236.6325 110.4225 236.7675 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.4625 236.6325 111.5975 236.7675 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.6375 236.6325 112.7725 236.7675 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.8125 236.6325 113.9475 236.7675 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.9875 236.6325 115.1225 236.7675 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.1625 236.6325 116.2975 236.7675 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.3375 236.6325 117.4725 236.7675 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.5125 236.6325 118.6475 236.7675 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.6875 236.6325 119.8225 236.7675 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.8625 236.6325 120.9975 236.7675 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.0375 236.6325 122.1725 236.7675 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.2125 236.6325 123.3475 236.7675 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.3875 236.6325 124.5225 236.7675 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.5625 236.6325 125.6975 236.7675 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.7375 236.6325 126.8725 236.7675 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.9125 236.6325 128.0475 236.7675 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.0875 236.6325 129.2225 236.7675 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.2625 236.6325 130.3975 236.7675 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.4375 236.6325 131.5725 236.7675 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.6125 236.6325 132.7475 236.7675 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.7875 236.6325 133.9225 236.7675 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.9625 236.6325 135.0975 236.7675 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.1375 236.6325 136.2725 236.7675 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.3125 236.6325 137.4475 236.7675 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.4875 236.6325 138.6225 236.7675 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.6625 236.6325 139.7975 236.7675 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.8375 236.6325 140.9725 236.7675 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.0125 236.6325 142.1475 236.7675 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.1875 236.6325 143.3225 236.7675 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.3625 236.6325 144.4975 236.7675 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.5375 236.6325 145.6725 236.7675 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.7125 236.6325 146.8475 236.7675 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.8875 236.6325 148.0225 236.7675 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.0625 236.6325 149.1975 236.7675 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.2375 236.6325 150.3725 236.7675 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.4125 236.6325 151.5475 236.7675 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.5875 236.6325 152.7225 236.7675 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.7625 236.6325 153.8975 236.7675 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.9375 236.6325 155.0725 236.7675 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.1125 236.6325 156.2475 236.7675 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.2875 236.6325 157.4225 236.7675 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.4625 236.6325 158.5975 236.7675 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.6375 236.6325 159.7725 236.7675 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.8125 236.6325 160.9475 236.7675 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.9875 236.6325 162.1225 236.7675 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.1625 236.6325 163.2975 236.7675 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.3375 236.6325 164.4725 236.7675 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.5125 236.6325 165.6475 236.7675 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.6875 236.6325 166.8225 236.7675 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.8625 236.6325 167.9975 236.7675 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.0375 236.6325 169.1725 236.7675 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.2125 236.6325 170.3475 236.7675 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.3875 236.6325 171.5225 236.7675 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.5625 236.6325 172.6975 236.7675 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.7375 236.6325 173.8725 236.7675 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.9125 236.6325 175.0475 236.7675 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.0875 236.6325 176.2225 236.7675 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.2625 236.6325 177.3975 236.7675 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.4375 236.6325 178.5725 236.7675 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.6125 236.6325 179.7475 236.7675 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.7875 236.6325 180.9225 236.7675 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.9625 236.6325 182.0975 236.7675 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.1375 236.6325 183.2725 236.7675 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.3125 236.6325 184.4475 236.7675 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.4875 236.6325 185.6225 236.7675 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.6625 236.6325 186.7975 236.7675 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.8375 236.6325 187.9725 236.7675 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.0125 236.6325 189.1475 236.7675 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.1875 236.6325 190.3225 236.7675 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.3625 236.6325 191.4975 236.7675 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.5375 236.6325 192.6725 236.7675 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.7125 236.6325 193.8475 236.7675 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.8875 236.6325 195.0225 236.7675 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.0625 236.6325 196.1975 236.7675 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.2375 236.6325 197.3725 236.7675 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.4125 236.6325 198.5475 236.7675 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.5875 236.6325 199.7225 236.7675 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.7625 236.6325 200.8975 236.7675 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.9375 236.6325 202.0725 236.7675 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.1125 236.6325 203.2475 236.7675 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.2875 236.6325 204.4225 236.7675 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.4625 236.6325 205.5975 236.7675 ;
      END
   END dout1[123]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  373.5925 2.47 373.7275 2.605 ;
         LAYER metal3 ;
         RECT  327.8325 2.47 327.9675 2.605 ;
         LAYER metal3 ;
         RECT  57.7525 25.765 206.2675 25.835 ;
         LAYER metal4 ;
         RECT  56.605 35.065 56.745 226.565 ;
         LAYER metal3 ;
         RECT  57.7525 234.0775 206.2675 234.1475 ;
         LAYER metal3 ;
         RECT  224.7325 57.4925 224.8675 57.6275 ;
         LAYER metal3 ;
         RECT  201.9925 2.47 202.1275 2.605 ;
         LAYER metal3 ;
         RECT  236.3125 2.47 236.4475 2.605 ;
         LAYER metal3 ;
         RECT  2.425 16.8675 2.56 17.0025 ;
         LAYER metal3 ;
         RECT  179.1125 2.47 179.2475 2.605 ;
         LAYER metal3 ;
         RECT  87.5925 2.47 87.7275 2.605 ;
         LAYER metal3 ;
         RECT  293.5125 2.47 293.6475 2.605 ;
         LAYER metal3 ;
         RECT  224.3875 45.5325 224.5225 45.6675 ;
         LAYER metal3 ;
         RECT  282.0725 2.47 282.2075 2.605 ;
         LAYER metal3 ;
         RECT  156.2325 2.47 156.3675 2.605 ;
         LAYER metal3 ;
         RECT  53.2725 2.47 53.4075 2.605 ;
         LAYER metal3 ;
         RECT  42.7725 60.4825 42.9075 60.6175 ;
         LAYER metal3 ;
         RECT  396.4725 2.47 396.6075 2.605 ;
         LAYER metal3 ;
         RECT  42.7725 63.4725 42.9075 63.6075 ;
         LAYER metal3 ;
         RECT  57.7525 31.2 206.7375 31.27 ;
         LAYER metal3 ;
         RECT  43.1175 48.5225 43.2525 48.6575 ;
         LAYER metal4 ;
         RECT  267.1475 212.335 267.2875 234.7375 ;
         LAYER metal4 ;
         RECT  231.585 17.71 231.725 35.205 ;
         LAYER metal3 ;
         RECT  121.9125 2.47 122.0475 2.605 ;
         LAYER metal3 ;
         RECT  49.85 34.36 49.985 34.495 ;
         LAYER metal3 ;
         RECT  385.0325 2.47 385.1675 2.605 ;
         LAYER metal3 ;
         RECT  224.8725 2.47 225.0075 2.605 ;
         LAYER metal4 ;
         RECT  210.895 35.065 211.035 226.565 ;
         LAYER metal3 ;
         RECT  41.8325 2.47 41.9675 2.605 ;
         LAYER metal3 ;
         RECT  247.7525 2.47 247.8875 2.605 ;
         LAYER metal4 ;
         RECT  209.815 31.895 209.955 229.485 ;
         LAYER metal4 ;
         RECT  218.27 35.065 218.41 226.635 ;
         LAYER metal3 ;
         RECT  224.7325 63.4725 224.8675 63.6075 ;
         LAYER metal3 ;
         RECT  316.3925 2.47 316.5275 2.605 ;
         LAYER metal3 ;
         RECT  190.5525 2.47 190.6875 2.605 ;
         LAYER metal3 ;
         RECT  224.3875 39.5525 224.5225 39.6875 ;
         LAYER metal3 ;
         RECT  57.6175 24.7975 57.7525 24.9325 ;
         LAYER metal4 ;
         RECT  0.6875 24.2425 0.8275 46.645 ;
         LAYER metal3 ;
         RECT  224.3875 48.5225 224.5225 48.6575 ;
         LAYER metal3 ;
         RECT  210.8975 227.9225 211.0325 228.0575 ;
         LAYER metal3 ;
         RECT  167.6725 2.47 167.8075 2.605 ;
         LAYER metal3 ;
         RECT  43.1175 36.5625 43.2525 36.6975 ;
         LAYER metal3 ;
         RECT  217.655 227.135 217.79 227.27 ;
         LAYER metal3 ;
         RECT  270.6325 2.47 270.7675 2.605 ;
         LAYER metal3 ;
         RECT  43.1175 45.5325 43.2525 45.6675 ;
         LAYER metal3 ;
         RECT  64.7125 2.47 64.8475 2.605 ;
         LAYER metal3 ;
         RECT  42.7725 57.4925 42.9075 57.6275 ;
         LAYER metal3 ;
         RECT  110.4725 2.47 110.6075 2.605 ;
         LAYER metal3 ;
         RECT  56.6075 33.5725 56.7425 33.7075 ;
         LAYER metal3 ;
         RECT  206.6025 24.7975 206.7375 24.9325 ;
         LAYER metal3 ;
         RECT  76.1525 2.47 76.2875 2.605 ;
         LAYER metal3 ;
         RECT  224.3875 36.5625 224.5225 36.6975 ;
         LAYER metal3 ;
         RECT  339.2725 2.47 339.4075 2.605 ;
         LAYER metal3 ;
         RECT  350.7125 2.47 350.8475 2.605 ;
         LAYER metal3 ;
         RECT  144.7925 2.47 144.9275 2.605 ;
         LAYER metal3 ;
         RECT  304.9525 2.47 305.0875 2.605 ;
         LAYER metal4 ;
         RECT  38.83 16.865 38.97 31.825 ;
         LAYER metal3 ;
         RECT  213.4325 2.47 213.5675 2.605 ;
         LAYER metal4 ;
         RECT  228.865 232.095 229.005 242.115 ;
         LAYER metal4 ;
         RECT  57.685 31.895 57.825 229.485 ;
         LAYER metal3 ;
         RECT  57.7525 230.18 207.9125 230.25 ;
         LAYER metal3 ;
         RECT  42.7725 54.5025 42.9075 54.6375 ;
         LAYER metal3 ;
         RECT  43.1175 39.5525 43.2525 39.6875 ;
         LAYER metal3 ;
         RECT  224.7325 54.5025 224.8675 54.6375 ;
         LAYER metal4 ;
         RECT  49.23 35.065 49.37 226.635 ;
         LAYER metal3 ;
         RECT  224.7325 60.4825 224.8675 60.6175 ;
         LAYER metal3 ;
         RECT  259.1925 2.47 259.3275 2.605 ;
         LAYER metal3 ;
         RECT  265.415 241.9775 265.55 242.1125 ;
         LAYER metal4 ;
         RECT  36.11 64.965 36.25 82.46 ;
         LAYER metal3 ;
         RECT  99.0325 2.47 99.1675 2.605 ;
         LAYER metal3 ;
         RECT  133.3525 2.47 133.4875 2.605 ;
         LAYER metal3 ;
         RECT  362.1525 2.47 362.2875 2.605 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  239.1725 0.0 239.3075 0.135 ;
         LAYER metal3 ;
         RECT  170.5325 0.0 170.6675 0.135 ;
         LAYER metal3 ;
         RECT  136.2125 0.0 136.3475 0.135 ;
         LAYER metal3 ;
         RECT  225.915 44.0375 226.05 44.1725 ;
         LAYER metal3 ;
         RECT  41.59 44.0375 41.725 44.1725 ;
         LAYER metal3 ;
         RECT  57.7525 27.815 206.2675 27.885 ;
         LAYER metal4 ;
         RECT  209.355 31.895 209.495 229.485 ;
         LAYER metal3 ;
         RECT  181.9725 0.0 182.1075 0.135 ;
         LAYER metal3 ;
         RECT  387.8925 0.0 388.0275 0.135 ;
         LAYER metal4 ;
         RECT  265.085 212.3025 265.225 234.705 ;
         LAYER metal3 ;
         RECT  225.915 35.0675 226.05 35.2025 ;
         LAYER metal3 ;
         RECT  273.4925 0.0 273.6275 0.135 ;
         LAYER metal3 ;
         RECT  226.54 64.9675 226.675 65.1025 ;
         LAYER metal3 ;
         RECT  399.3325 0.0 399.4675 0.135 ;
         LAYER metal3 ;
         RECT  159.0925 0.0 159.2275 0.135 ;
         LAYER metal4 ;
         RECT  6.105 14.395 6.245 29.355 ;
         LAYER metal3 ;
         RECT  226.54 53.0075 226.675 53.1425 ;
         LAYER metal4 ;
         RECT  49.79 35.0325 49.93 226.5975 ;
         LAYER metal3 ;
         RECT  342.1325 0.0 342.2675 0.135 ;
         LAYER metal3 ;
         RECT  41.59 50.0175 41.725 50.1525 ;
         LAYER metal3 ;
         RECT  225.915 47.0275 226.05 47.1625 ;
         LAYER metal3 ;
         RECT  2.425 14.3975 2.56 14.5325 ;
         LAYER metal3 ;
         RECT  284.9325 0.0 285.0675 0.135 ;
         LAYER metal3 ;
         RECT  67.5725 0.0 67.7075 0.135 ;
         LAYER metal3 ;
         RECT  250.6125 0.0 250.7475 0.135 ;
         LAYER metal3 ;
         RECT  307.8125 0.0 307.9475 0.135 ;
         LAYER metal3 ;
         RECT  227.7325 0.0 227.8675 0.135 ;
         LAYER metal3 ;
         RECT  41.59 47.0275 41.725 47.1625 ;
         LAYER metal3 ;
         RECT  353.5725 0.0 353.7075 0.135 ;
         LAYER metal3 ;
         RECT  296.3725 0.0 296.5075 0.135 ;
         LAYER metal4 ;
         RECT  217.71 35.0325 217.85 226.5975 ;
         LAYER metal3 ;
         RECT  57.7525 232.185 206.3025 232.255 ;
         LAYER metal3 ;
         RECT  40.965 55.9975 41.1 56.1325 ;
         LAYER metal3 ;
         RECT  226.54 55.9975 226.675 56.1325 ;
         LAYER metal3 ;
         RECT  113.3325 0.0 113.4675 0.135 ;
         LAYER metal3 ;
         RECT  206.6025 22.9775 206.7375 23.1125 ;
         LAYER metal4 ;
         RECT  58.145 31.895 58.285 229.485 ;
         LAYER metal3 ;
         RECT  41.59 38.0575 41.725 38.1925 ;
         LAYER metal3 ;
         RECT  226.54 61.9775 226.675 62.1125 ;
         LAYER metal3 ;
         RECT  330.6925 0.0 330.8275 0.135 ;
         LAYER metal4 ;
         RECT  261.59 229.625 261.73 244.585 ;
         LAYER metal3 ;
         RECT  90.4525 0.0 90.5875 0.135 ;
         LAYER metal3 ;
         RECT  262.0525 0.0 262.1875 0.135 ;
         LAYER metal3 ;
         RECT  376.4525 0.0 376.5875 0.135 ;
         LAYER metal3 ;
         RECT  124.7725 0.0 124.9075 0.135 ;
         LAYER metal3 ;
         RECT  147.6525 0.0 147.7875 0.135 ;
         LAYER metal3 ;
         RECT  204.8525 0.0 204.9875 0.135 ;
         LAYER metal3 ;
         RECT  44.6925 0.0 44.8275 0.135 ;
         LAYER metal3 ;
         RECT  193.4125 0.0 193.5475 0.135 ;
         LAYER metal4 ;
         RECT  220.205 35.0325 220.345 226.635 ;
         LAYER metal3 ;
         RECT  216.2925 0.0 216.4275 0.135 ;
         LAYER metal4 ;
         RECT  228.725 17.775 228.865 35.27 ;
         LAYER metal3 ;
         RECT  225.915 38.0575 226.05 38.1925 ;
         LAYER metal3 ;
         RECT  226.54 58.9875 226.675 59.1225 ;
         LAYER metal3 ;
         RECT  41.59 35.0675 41.725 35.2025 ;
         LAYER metal3 ;
         RECT  56.1325 0.0 56.2675 0.135 ;
         LAYER metal3 ;
         RECT  79.0125 0.0 79.1475 0.135 ;
         LAYER metal3 ;
         RECT  365.0125 0.0 365.1475 0.135 ;
         LAYER metal3 ;
         RECT  57.6175 22.9775 57.7525 23.1125 ;
         LAYER metal3 ;
         RECT  225.915 41.0475 226.05 41.1825 ;
         LAYER metal3 ;
         RECT  40.965 64.9675 41.1 65.1025 ;
         LAYER metal3 ;
         RECT  225.915 50.0175 226.05 50.1525 ;
         LAYER metal4 ;
         RECT  38.97 64.9 39.11 82.395 ;
         LAYER metal3 ;
         RECT  40.965 58.9875 41.1 59.1225 ;
         LAYER metal3 ;
         RECT  319.2525 0.0 319.3875 0.135 ;
         LAYER metal3 ;
         RECT  41.59 41.0475 41.725 41.1825 ;
         LAYER metal4 ;
         RECT  47.295 35.0325 47.435 226.635 ;
         LAYER metal3 ;
         RECT  40.965 53.0075 41.1 53.1425 ;
         LAYER metal3 ;
         RECT  101.8925 0.0 102.0275 0.135 ;
         LAYER metal4 ;
         RECT  2.75 24.275 2.89 46.6775 ;
         LAYER metal3 ;
         RECT  265.415 244.4475 265.55 244.5825 ;
         LAYER metal3 ;
         RECT  40.965 61.9775 41.1 62.1125 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 407.84 244.445 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 407.84 244.445 ;
   LAYER  metal3 ;
      RECT  53.415 0.14 53.83 0.965 ;
      RECT  53.83 0.965 56.275 1.38 ;
      RECT  56.69 0.965 59.135 1.38 ;
      RECT  59.55 0.965 61.995 1.38 ;
      RECT  62.41 0.965 64.855 1.38 ;
      RECT  65.27 0.965 67.715 1.38 ;
      RECT  68.13 0.965 70.575 1.38 ;
      RECT  70.99 0.965 73.435 1.38 ;
      RECT  73.85 0.965 76.295 1.38 ;
      RECT  76.71 0.965 79.155 1.38 ;
      RECT  79.57 0.965 82.015 1.38 ;
      RECT  82.43 0.965 84.875 1.38 ;
      RECT  85.29 0.965 87.735 1.38 ;
      RECT  88.15 0.965 90.595 1.38 ;
      RECT  91.01 0.965 93.455 1.38 ;
      RECT  93.87 0.965 96.315 1.38 ;
      RECT  96.73 0.965 99.175 1.38 ;
      RECT  99.59 0.965 102.035 1.38 ;
      RECT  102.45 0.965 104.895 1.38 ;
      RECT  105.31 0.965 107.755 1.38 ;
      RECT  108.17 0.965 110.615 1.38 ;
      RECT  111.03 0.965 113.475 1.38 ;
      RECT  113.89 0.965 116.335 1.38 ;
      RECT  116.75 0.965 119.195 1.38 ;
      RECT  119.61 0.965 122.055 1.38 ;
      RECT  122.47 0.965 124.915 1.38 ;
      RECT  125.33 0.965 127.775 1.38 ;
      RECT  128.19 0.965 130.635 1.38 ;
      RECT  131.05 0.965 133.495 1.38 ;
      RECT  133.91 0.965 136.355 1.38 ;
      RECT  136.77 0.965 139.215 1.38 ;
      RECT  139.63 0.965 142.075 1.38 ;
      RECT  142.49 0.965 144.935 1.38 ;
      RECT  145.35 0.965 147.795 1.38 ;
      RECT  148.21 0.965 150.655 1.38 ;
      RECT  151.07 0.965 153.515 1.38 ;
      RECT  153.93 0.965 156.375 1.38 ;
      RECT  156.79 0.965 159.235 1.38 ;
      RECT  159.65 0.965 162.095 1.38 ;
      RECT  162.51 0.965 164.955 1.38 ;
      RECT  165.37 0.965 167.815 1.38 ;
      RECT  168.23 0.965 170.675 1.38 ;
      RECT  171.09 0.965 173.535 1.38 ;
      RECT  173.95 0.965 176.395 1.38 ;
      RECT  176.81 0.965 179.255 1.38 ;
      RECT  179.67 0.965 182.115 1.38 ;
      RECT  182.53 0.965 184.975 1.38 ;
      RECT  185.39 0.965 187.835 1.38 ;
      RECT  188.25 0.965 190.695 1.38 ;
      RECT  191.11 0.965 193.555 1.38 ;
      RECT  193.97 0.965 196.415 1.38 ;
      RECT  196.83 0.965 199.275 1.38 ;
      RECT  199.69 0.965 202.135 1.38 ;
      RECT  202.55 0.965 204.995 1.38 ;
      RECT  205.41 0.965 207.855 1.38 ;
      RECT  208.27 0.965 210.715 1.38 ;
      RECT  211.13 0.965 213.575 1.38 ;
      RECT  213.99 0.965 216.435 1.38 ;
      RECT  216.85 0.965 219.295 1.38 ;
      RECT  219.71 0.965 222.155 1.38 ;
      RECT  222.57 0.965 225.015 1.38 ;
      RECT  225.43 0.965 227.875 1.38 ;
      RECT  228.29 0.965 230.735 1.38 ;
      RECT  231.15 0.965 233.595 1.38 ;
      RECT  234.01 0.965 236.455 1.38 ;
      RECT  236.87 0.965 239.315 1.38 ;
      RECT  239.73 0.965 242.175 1.38 ;
      RECT  242.59 0.965 245.035 1.38 ;
      RECT  245.45 0.965 247.895 1.38 ;
      RECT  248.31 0.965 250.755 1.38 ;
      RECT  251.17 0.965 253.615 1.38 ;
      RECT  254.03 0.965 256.475 1.38 ;
      RECT  256.89 0.965 259.335 1.38 ;
      RECT  259.75 0.965 262.195 1.38 ;
      RECT  262.61 0.965 265.055 1.38 ;
      RECT  265.47 0.965 267.915 1.38 ;
      RECT  268.33 0.965 270.775 1.38 ;
      RECT  271.19 0.965 273.635 1.38 ;
      RECT  274.05 0.965 276.495 1.38 ;
      RECT  276.91 0.965 279.355 1.38 ;
      RECT  279.77 0.965 282.215 1.38 ;
      RECT  282.63 0.965 285.075 1.38 ;
      RECT  285.49 0.965 287.935 1.38 ;
      RECT  288.35 0.965 290.795 1.38 ;
      RECT  291.21 0.965 293.655 1.38 ;
      RECT  294.07 0.965 296.515 1.38 ;
      RECT  296.93 0.965 299.375 1.38 ;
      RECT  299.79 0.965 302.235 1.38 ;
      RECT  302.65 0.965 305.095 1.38 ;
      RECT  305.51 0.965 307.955 1.38 ;
      RECT  308.37 0.965 310.815 1.38 ;
      RECT  311.23 0.965 313.675 1.38 ;
      RECT  314.09 0.965 316.535 1.38 ;
      RECT  316.95 0.965 319.395 1.38 ;
      RECT  319.81 0.965 322.255 1.38 ;
      RECT  322.67 0.965 325.115 1.38 ;
      RECT  325.53 0.965 327.975 1.38 ;
      RECT  328.39 0.965 330.835 1.38 ;
      RECT  331.25 0.965 333.695 1.38 ;
      RECT  334.11 0.965 336.555 1.38 ;
      RECT  336.97 0.965 339.415 1.38 ;
      RECT  339.83 0.965 342.275 1.38 ;
      RECT  342.69 0.965 345.135 1.38 ;
      RECT  345.55 0.965 347.995 1.38 ;
      RECT  348.41 0.965 350.855 1.38 ;
      RECT  351.27 0.965 353.715 1.38 ;
      RECT  354.13 0.965 356.575 1.38 ;
      RECT  356.99 0.965 359.435 1.38 ;
      RECT  359.85 0.965 362.295 1.38 ;
      RECT  362.71 0.965 365.155 1.38 ;
      RECT  365.57 0.965 368.015 1.38 ;
      RECT  368.43 0.965 370.875 1.38 ;
      RECT  371.29 0.965 373.735 1.38 ;
      RECT  374.15 0.965 376.595 1.38 ;
      RECT  377.01 0.965 379.455 1.38 ;
      RECT  379.87 0.965 382.315 1.38 ;
      RECT  382.73 0.965 385.175 1.38 ;
      RECT  385.59 0.965 388.035 1.38 ;
      RECT  388.45 0.965 390.895 1.38 ;
      RECT  391.31 0.965 393.755 1.38 ;
      RECT  394.17 0.965 396.615 1.38 ;
      RECT  397.03 0.965 399.475 1.38 ;
      RECT  399.89 0.965 402.335 1.38 ;
      RECT  402.75 0.965 405.195 1.38 ;
      RECT  405.61 0.965 407.84 1.38 ;
      RECT  0.14 65.9325 36.255 66.3475 ;
      RECT  0.14 66.3475 36.255 244.445 ;
      RECT  36.255 1.38 36.67 65.9325 ;
      RECT  36.67 65.9325 53.415 66.3475 ;
      RECT  36.67 66.3475 53.415 244.445 ;
      RECT  36.255 66.3475 36.67 68.6625 ;
      RECT  36.255 69.0775 36.67 70.8725 ;
      RECT  36.255 71.2875 36.67 73.6025 ;
      RECT  36.255 74.0175 36.67 75.8125 ;
      RECT  36.255 76.2275 36.67 78.5425 ;
      RECT  36.255 78.9575 36.67 80.7525 ;
      RECT  36.255 81.1675 36.67 244.445 ;
      RECT  231.165 34.2375 231.58 244.445 ;
      RECT  231.58 33.8225 407.84 34.2375 ;
      RECT  231.165 31.5075 231.58 33.8225 ;
      RECT  231.165 29.2975 231.58 31.0925 ;
      RECT  231.165 26.5675 231.58 28.8825 ;
      RECT  231.165 24.3575 231.58 26.1525 ;
      RECT  231.165 21.6275 231.58 23.9425 ;
      RECT  231.165 1.38 231.58 19.0025 ;
      RECT  231.165 19.4175 231.58 21.2125 ;
      RECT  0.14 1.38 0.145 15.3625 ;
      RECT  0.14 15.3625 0.145 15.7775 ;
      RECT  0.14 15.7775 0.145 65.9325 ;
      RECT  0.145 1.38 0.56 15.3625 ;
      RECT  0.145 15.7775 0.56 65.9325 ;
      RECT  267.415 34.2375 267.83 243.2025 ;
      RECT  267.415 243.6175 267.83 244.445 ;
      RECT  267.83 34.2375 407.84 243.2025 ;
      RECT  267.83 243.2025 407.84 243.6175 ;
      RECT  267.83 243.6175 407.84 244.445 ;
      RECT  0.56 15.3625 6.1075 15.4475 ;
      RECT  0.56 15.4475 6.1075 15.7775 ;
      RECT  6.1075 15.3625 6.5225 15.4475 ;
      RECT  6.5225 15.3625 36.255 15.4475 ;
      RECT  6.5225 15.4475 36.255 15.7775 ;
      RECT  0.56 15.7775 6.1075 15.8625 ;
      RECT  6.1075 15.8625 6.5225 65.9325 ;
      RECT  6.5225 15.7775 36.255 15.8625 ;
      RECT  6.5225 15.8625 36.255 65.9325 ;
      RECT  231.58 34.2375 261.3125 243.1175 ;
      RECT  231.58 243.1175 261.3125 243.2025 ;
      RECT  261.3125 34.2375 261.7275 243.1175 ;
      RECT  261.7275 243.1175 267.415 243.2025 ;
      RECT  231.58 243.2025 261.3125 243.5325 ;
      RECT  231.58 243.5325 261.3125 243.6175 ;
      RECT  261.3125 243.5325 261.7275 243.6175 ;
      RECT  261.7275 243.2025 267.415 243.5325 ;
      RECT  261.7275 243.5325 267.415 243.6175 ;
      RECT  0.14 0.965 41.975 1.38 ;
      RECT  42.39 0.965 44.835 1.38 ;
      RECT  45.25 0.965 47.695 1.38 ;
      RECT  48.11 0.965 50.555 1.38 ;
      RECT  50.97 0.965 53.415 1.38 ;
      RECT  53.83 236.4925 60.7975 236.9075 ;
      RECT  53.83 236.9075 60.7975 244.445 ;
      RECT  60.7975 236.9075 61.2125 244.445 ;
      RECT  61.2125 236.9075 231.165 244.445 ;
      RECT  61.2125 236.4925 61.9725 236.9075 ;
      RECT  62.3875 236.4925 63.1475 236.9075 ;
      RECT  63.5625 236.4925 64.3225 236.9075 ;
      RECT  64.7375 236.4925 65.4975 236.9075 ;
      RECT  65.9125 236.4925 66.6725 236.9075 ;
      RECT  67.0875 236.4925 67.8475 236.9075 ;
      RECT  68.2625 236.4925 69.0225 236.9075 ;
      RECT  69.4375 236.4925 70.1975 236.9075 ;
      RECT  70.6125 236.4925 71.3725 236.9075 ;
      RECT  71.7875 236.4925 72.5475 236.9075 ;
      RECT  72.9625 236.4925 73.7225 236.9075 ;
      RECT  74.1375 236.4925 74.8975 236.9075 ;
      RECT  75.3125 236.4925 76.0725 236.9075 ;
      RECT  76.4875 236.4925 77.2475 236.9075 ;
      RECT  77.6625 236.4925 78.4225 236.9075 ;
      RECT  78.8375 236.4925 79.5975 236.9075 ;
      RECT  80.0125 236.4925 80.7725 236.9075 ;
      RECT  81.1875 236.4925 81.9475 236.9075 ;
      RECT  82.3625 236.4925 83.1225 236.9075 ;
      RECT  83.5375 236.4925 84.2975 236.9075 ;
      RECT  84.7125 236.4925 85.4725 236.9075 ;
      RECT  85.8875 236.4925 86.6475 236.9075 ;
      RECT  87.0625 236.4925 87.8225 236.9075 ;
      RECT  88.2375 236.4925 88.9975 236.9075 ;
      RECT  89.4125 236.4925 90.1725 236.9075 ;
      RECT  90.5875 236.4925 91.3475 236.9075 ;
      RECT  91.7625 236.4925 92.5225 236.9075 ;
      RECT  92.9375 236.4925 93.6975 236.9075 ;
      RECT  94.1125 236.4925 94.8725 236.9075 ;
      RECT  95.2875 236.4925 96.0475 236.9075 ;
      RECT  96.4625 236.4925 97.2225 236.9075 ;
      RECT  97.6375 236.4925 98.3975 236.9075 ;
      RECT  98.8125 236.4925 99.5725 236.9075 ;
      RECT  99.9875 236.4925 100.7475 236.9075 ;
      RECT  101.1625 236.4925 101.9225 236.9075 ;
      RECT  102.3375 236.4925 103.0975 236.9075 ;
      RECT  103.5125 236.4925 104.2725 236.9075 ;
      RECT  104.6875 236.4925 105.4475 236.9075 ;
      RECT  105.8625 236.4925 106.6225 236.9075 ;
      RECT  107.0375 236.4925 107.7975 236.9075 ;
      RECT  108.2125 236.4925 108.9725 236.9075 ;
      RECT  109.3875 236.4925 110.1475 236.9075 ;
      RECT  110.5625 236.4925 111.3225 236.9075 ;
      RECT  111.7375 236.4925 112.4975 236.9075 ;
      RECT  112.9125 236.4925 113.6725 236.9075 ;
      RECT  114.0875 236.4925 114.8475 236.9075 ;
      RECT  115.2625 236.4925 116.0225 236.9075 ;
      RECT  116.4375 236.4925 117.1975 236.9075 ;
      RECT  117.6125 236.4925 118.3725 236.9075 ;
      RECT  118.7875 236.4925 119.5475 236.9075 ;
      RECT  119.9625 236.4925 120.7225 236.9075 ;
      RECT  121.1375 236.4925 121.8975 236.9075 ;
      RECT  122.3125 236.4925 123.0725 236.9075 ;
      RECT  123.4875 236.4925 124.2475 236.9075 ;
      RECT  124.6625 236.4925 125.4225 236.9075 ;
      RECT  125.8375 236.4925 126.5975 236.9075 ;
      RECT  127.0125 236.4925 127.7725 236.9075 ;
      RECT  128.1875 236.4925 128.9475 236.9075 ;
      RECT  129.3625 236.4925 130.1225 236.9075 ;
      RECT  130.5375 236.4925 131.2975 236.9075 ;
      RECT  131.7125 236.4925 132.4725 236.9075 ;
      RECT  132.8875 236.4925 133.6475 236.9075 ;
      RECT  134.0625 236.4925 134.8225 236.9075 ;
      RECT  135.2375 236.4925 135.9975 236.9075 ;
      RECT  136.4125 236.4925 137.1725 236.9075 ;
      RECT  137.5875 236.4925 138.3475 236.9075 ;
      RECT  138.7625 236.4925 139.5225 236.9075 ;
      RECT  139.9375 236.4925 140.6975 236.9075 ;
      RECT  141.1125 236.4925 141.8725 236.9075 ;
      RECT  142.2875 236.4925 143.0475 236.9075 ;
      RECT  143.4625 236.4925 144.2225 236.9075 ;
      RECT  144.6375 236.4925 145.3975 236.9075 ;
      RECT  145.8125 236.4925 146.5725 236.9075 ;
      RECT  146.9875 236.4925 147.7475 236.9075 ;
      RECT  148.1625 236.4925 148.9225 236.9075 ;
      RECT  149.3375 236.4925 150.0975 236.9075 ;
      RECT  150.5125 236.4925 151.2725 236.9075 ;
      RECT  151.6875 236.4925 152.4475 236.9075 ;
      RECT  152.8625 236.4925 153.6225 236.9075 ;
      RECT  154.0375 236.4925 154.7975 236.9075 ;
      RECT  155.2125 236.4925 155.9725 236.9075 ;
      RECT  156.3875 236.4925 157.1475 236.9075 ;
      RECT  157.5625 236.4925 158.3225 236.9075 ;
      RECT  158.7375 236.4925 159.4975 236.9075 ;
      RECT  159.9125 236.4925 160.6725 236.9075 ;
      RECT  161.0875 236.4925 161.8475 236.9075 ;
      RECT  162.2625 236.4925 163.0225 236.9075 ;
      RECT  163.4375 236.4925 164.1975 236.9075 ;
      RECT  164.6125 236.4925 165.3725 236.9075 ;
      RECT  165.7875 236.4925 166.5475 236.9075 ;
      RECT  166.9625 236.4925 167.7225 236.9075 ;
      RECT  168.1375 236.4925 168.8975 236.9075 ;
      RECT  169.3125 236.4925 170.0725 236.9075 ;
      RECT  170.4875 236.4925 171.2475 236.9075 ;
      RECT  171.6625 236.4925 172.4225 236.9075 ;
      RECT  172.8375 236.4925 173.5975 236.9075 ;
      RECT  174.0125 236.4925 174.7725 236.9075 ;
      RECT  175.1875 236.4925 175.9475 236.9075 ;
      RECT  176.3625 236.4925 177.1225 236.9075 ;
      RECT  177.5375 236.4925 178.2975 236.9075 ;
      RECT  178.7125 236.4925 179.4725 236.9075 ;
      RECT  179.8875 236.4925 180.6475 236.9075 ;
      RECT  181.0625 236.4925 181.8225 236.9075 ;
      RECT  182.2375 236.4925 182.9975 236.9075 ;
      RECT  183.4125 236.4925 184.1725 236.9075 ;
      RECT  184.5875 236.4925 185.3475 236.9075 ;
      RECT  185.7625 236.4925 186.5225 236.9075 ;
      RECT  186.9375 236.4925 187.6975 236.9075 ;
      RECT  188.1125 236.4925 188.8725 236.9075 ;
      RECT  189.2875 236.4925 190.0475 236.9075 ;
      RECT  190.4625 236.4925 191.2225 236.9075 ;
      RECT  191.6375 236.4925 192.3975 236.9075 ;
      RECT  192.8125 236.4925 193.5725 236.9075 ;
      RECT  193.9875 236.4925 194.7475 236.9075 ;
      RECT  195.1625 236.4925 195.9225 236.9075 ;
      RECT  196.3375 236.4925 197.0975 236.9075 ;
      RECT  197.5125 236.4925 198.2725 236.9075 ;
      RECT  198.6875 236.4925 199.4475 236.9075 ;
      RECT  199.8625 236.4925 200.6225 236.9075 ;
      RECT  201.0375 236.4925 201.7975 236.9075 ;
      RECT  202.2125 236.4925 202.9725 236.9075 ;
      RECT  203.3875 236.4925 204.1475 236.9075 ;
      RECT  204.5625 236.4925 205.3225 236.9075 ;
      RECT  205.7375 236.4925 231.165 236.9075 ;
      RECT  231.58 1.38 373.4525 2.33 ;
      RECT  231.58 2.745 373.4525 33.8225 ;
      RECT  373.4525 1.38 373.8675 2.33 ;
      RECT  373.4525 2.745 373.8675 33.8225 ;
      RECT  373.8675 1.38 407.84 2.33 ;
      RECT  373.8675 2.745 407.84 33.8225 ;
      RECT  53.83 25.625 57.6125 25.975 ;
      RECT  206.4075 25.625 231.165 25.975 ;
      RECT  53.83 34.2375 57.6125 233.9375 ;
      RECT  53.83 233.9375 57.6125 234.2875 ;
      RECT  53.83 234.2875 57.6125 236.4925 ;
      RECT  57.6125 234.2875 60.7975 236.4925 ;
      RECT  60.7975 234.2875 61.2125 236.4925 ;
      RECT  61.2125 234.2875 206.4075 236.4925 ;
      RECT  206.4075 233.9375 231.165 234.2875 ;
      RECT  206.4075 234.2875 231.165 236.4925 ;
      RECT  206.4075 57.3525 224.5925 57.7675 ;
      RECT  225.0075 57.3525 231.165 57.7675 ;
      RECT  57.6125 1.38 201.8525 2.33 ;
      RECT  201.8525 1.38 202.2675 2.33 ;
      RECT  201.8525 2.745 202.2675 25.625 ;
      RECT  202.2675 1.38 206.4075 2.33 ;
      RECT  202.2675 2.33 206.4075 2.745 ;
      RECT  202.2675 2.745 206.4075 25.625 ;
      RECT  231.58 2.33 236.1725 2.745 ;
      RECT  0.56 15.8625 2.285 16.7275 ;
      RECT  0.56 16.7275 2.285 17.1425 ;
      RECT  0.56 17.1425 2.285 65.9325 ;
      RECT  2.285 15.8625 2.7 16.7275 ;
      RECT  2.285 17.1425 2.7 65.9325 ;
      RECT  2.7 15.8625 6.1075 16.7275 ;
      RECT  2.7 16.7275 6.1075 17.1425 ;
      RECT  2.7 17.1425 6.1075 65.9325 ;
      RECT  206.4075 34.2375 224.2475 45.3925 ;
      RECT  206.4075 45.3925 224.2475 45.8075 ;
      RECT  206.4075 45.8075 224.2475 57.3525 ;
      RECT  224.6625 34.2375 225.0075 45.3925 ;
      RECT  224.6625 45.3925 225.0075 45.8075 ;
      RECT  282.3475 2.33 293.3725 2.745 ;
      RECT  53.415 1.38 53.5475 2.33 ;
      RECT  53.415 2.745 53.5475 244.445 ;
      RECT  53.5475 1.38 53.83 2.33 ;
      RECT  53.5475 2.33 53.83 2.745 ;
      RECT  53.5475 2.745 53.83 244.445 ;
      RECT  36.67 1.38 53.1325 2.33 ;
      RECT  53.1325 1.38 53.415 2.33 ;
      RECT  53.1325 2.745 53.415 65.9325 ;
      RECT  36.67 60.3425 42.6325 60.7575 ;
      RECT  43.0475 60.3425 53.1325 60.7575 ;
      RECT  43.0475 60.7575 53.1325 65.9325 ;
      RECT  396.7475 2.33 407.84 2.745 ;
      RECT  42.6325 60.7575 43.0475 63.3325 ;
      RECT  42.6325 63.7475 43.0475 65.9325 ;
      RECT  57.6125 31.41 206.4075 33.8225 ;
      RECT  206.4075 25.975 206.8775 31.06 ;
      RECT  206.4075 31.41 206.8775 33.8225 ;
      RECT  206.8775 25.975 231.165 31.06 ;
      RECT  206.8775 31.06 231.165 31.41 ;
      RECT  206.8775 31.41 231.165 33.8225 ;
      RECT  42.6325 2.745 42.9775 48.3825 ;
      RECT  42.6325 48.3825 42.9775 48.7975 ;
      RECT  43.0475 48.7975 43.3925 60.3425 ;
      RECT  43.3925 48.3825 53.1325 48.7975 ;
      RECT  43.3925 48.7975 53.1325 60.3425 ;
      RECT  43.3925 2.745 49.71 34.22 ;
      RECT  43.3925 34.22 49.71 34.635 ;
      RECT  43.3925 34.635 49.71 48.3825 ;
      RECT  49.71 2.745 50.125 34.22 ;
      RECT  49.71 34.635 50.125 48.3825 ;
      RECT  50.125 2.745 53.1325 34.22 ;
      RECT  50.125 34.22 53.1325 34.635 ;
      RECT  50.125 34.635 53.1325 48.3825 ;
      RECT  373.8675 2.33 384.8925 2.745 ;
      RECT  385.3075 2.33 396.3325 2.745 ;
      RECT  206.4075 1.38 224.7325 2.33 ;
      RECT  224.7325 1.38 225.1475 2.33 ;
      RECT  224.7325 2.745 225.1475 25.625 ;
      RECT  225.1475 1.38 231.165 2.33 ;
      RECT  225.1475 2.33 231.165 2.745 ;
      RECT  225.1475 2.745 231.165 25.625 ;
      RECT  36.67 2.33 41.6925 2.745 ;
      RECT  42.1075 2.33 53.1325 2.745 ;
      RECT  236.5875 2.33 247.6125 2.745 ;
      RECT  224.5925 63.7475 225.0075 233.9375 ;
      RECT  316.6675 2.33 327.6925 2.745 ;
      RECT  179.3875 2.33 190.4125 2.745 ;
      RECT  190.8275 2.33 201.8525 2.745 ;
      RECT  224.2475 39.8275 224.5925 45.3925 ;
      RECT  224.5925 39.8275 224.6625 45.3925 ;
      RECT  53.83 1.38 57.4775 24.6575 ;
      RECT  53.83 24.6575 57.4775 25.0725 ;
      RECT  53.83 25.0725 57.4775 25.625 ;
      RECT  57.4775 25.0725 57.6125 25.625 ;
      RECT  57.6125 25.0725 57.8925 25.625 ;
      RECT  57.8925 2.745 201.8525 24.6575 ;
      RECT  57.8925 24.6575 201.8525 25.0725 ;
      RECT  57.8925 25.0725 201.8525 25.625 ;
      RECT  224.2475 45.8075 224.5925 48.3825 ;
      RECT  224.2475 48.7975 224.5925 57.3525 ;
      RECT  224.5925 45.8075 224.6625 48.3825 ;
      RECT  206.4075 57.7675 210.7575 227.7825 ;
      RECT  206.4075 227.7825 210.7575 228.1975 ;
      RECT  210.7575 57.7675 211.1725 227.7825 ;
      RECT  210.7575 228.1975 211.1725 233.9375 ;
      RECT  211.1725 227.7825 224.5925 228.1975 ;
      RECT  211.1725 228.1975 224.5925 233.9375 ;
      RECT  156.5075 2.33 167.5325 2.745 ;
      RECT  167.9475 2.33 178.9725 2.745 ;
      RECT  42.9775 2.745 43.0475 36.4225 ;
      RECT  43.0475 2.745 43.3925 36.4225 ;
      RECT  211.1725 57.7675 217.515 226.995 ;
      RECT  211.1725 226.995 217.515 227.41 ;
      RECT  211.1725 227.41 217.515 227.7825 ;
      RECT  217.515 57.7675 217.93 226.995 ;
      RECT  217.515 227.41 217.93 227.7825 ;
      RECT  217.93 57.7675 224.5925 226.995 ;
      RECT  217.93 226.995 224.5925 227.41 ;
      RECT  217.93 227.41 224.5925 227.7825 ;
      RECT  270.9075 2.33 281.9325 2.745 ;
      RECT  42.9775 45.8075 43.0475 48.3825 ;
      RECT  43.0475 45.8075 43.3925 48.3825 ;
      RECT  57.6125 2.33 64.5725 2.745 ;
      RECT  42.6325 57.7675 42.9775 60.3425 ;
      RECT  42.9775 57.7675 43.0475 60.3425 ;
      RECT  110.7475 2.33 121.7725 2.745 ;
      RECT  53.83 33.8225 56.4675 33.8475 ;
      RECT  53.83 33.8475 56.4675 34.2375 ;
      RECT  56.4675 33.8475 56.8825 34.2375 ;
      RECT  56.8825 33.8225 231.165 33.8475 ;
      RECT  56.8825 33.8475 231.165 34.2375 ;
      RECT  53.83 25.975 56.4675 33.4325 ;
      RECT  53.83 33.4325 56.4675 33.8225 ;
      RECT  56.4675 25.975 56.8825 33.4325 ;
      RECT  56.8825 25.975 57.6125 33.4325 ;
      RECT  56.8825 33.4325 57.6125 33.8225 ;
      RECT  206.4075 2.745 206.4625 24.6575 ;
      RECT  206.4075 24.6575 206.4625 25.0725 ;
      RECT  206.4075 25.0725 206.4625 25.625 ;
      RECT  206.4625 25.0725 206.8775 25.625 ;
      RECT  206.8775 2.745 224.7325 24.6575 ;
      RECT  206.8775 24.6575 224.7325 25.0725 ;
      RECT  206.8775 25.0725 224.7325 25.625 ;
      RECT  64.9875 2.33 76.0125 2.745 ;
      RECT  76.4275 2.33 87.4525 2.745 ;
      RECT  224.2475 34.2375 224.5925 36.4225 ;
      RECT  224.2475 36.8375 224.5925 39.4125 ;
      RECT  224.5925 34.2375 224.6625 36.4225 ;
      RECT  224.5925 36.8375 224.6625 39.4125 ;
      RECT  328.1075 2.33 339.1325 2.745 ;
      RECT  339.5475 2.33 350.5725 2.745 ;
      RECT  145.0675 2.33 156.0925 2.745 ;
      RECT  293.7875 2.33 304.8125 2.745 ;
      RECT  305.2275 2.33 316.2525 2.745 ;
      RECT  206.4075 2.33 213.2925 2.745 ;
      RECT  213.7075 2.33 224.7325 2.745 ;
      RECT  57.6125 34.2375 60.7975 230.04 ;
      RECT  60.7975 34.2375 61.2125 230.04 ;
      RECT  61.2125 34.2375 206.4075 230.04 ;
      RECT  206.4075 228.1975 208.0525 230.04 ;
      RECT  208.0525 228.1975 210.7575 230.04 ;
      RECT  208.0525 230.04 210.7575 230.39 ;
      RECT  208.0525 230.39 210.7575 233.9375 ;
      RECT  42.6325 48.7975 42.9775 54.3625 ;
      RECT  42.6325 54.7775 42.9775 57.3525 ;
      RECT  42.9775 48.7975 43.0475 54.3625 ;
      RECT  42.9775 54.7775 43.0475 57.3525 ;
      RECT  42.9775 36.8375 43.0475 39.4125 ;
      RECT  42.9775 39.8275 43.0475 45.3925 ;
      RECT  43.0475 36.8375 43.3925 39.4125 ;
      RECT  43.0475 39.8275 43.3925 45.3925 ;
      RECT  224.6625 45.8075 225.0075 54.3625 ;
      RECT  224.6625 54.7775 225.0075 57.3525 ;
      RECT  224.5925 48.7975 224.6625 54.3625 ;
      RECT  224.5925 54.7775 224.6625 57.3525 ;
      RECT  224.5925 57.7675 225.0075 60.3425 ;
      RECT  224.5925 60.7575 225.0075 63.3325 ;
      RECT  248.0275 2.33 259.0525 2.745 ;
      RECT  259.4675 2.33 270.4925 2.745 ;
      RECT  261.7275 34.2375 265.275 241.8375 ;
      RECT  261.7275 241.8375 265.275 242.2525 ;
      RECT  261.7275 242.2525 265.275 243.1175 ;
      RECT  265.275 34.2375 265.69 241.8375 ;
      RECT  265.275 242.2525 265.69 243.1175 ;
      RECT  265.69 34.2375 267.415 241.8375 ;
      RECT  265.69 241.8375 267.415 242.2525 ;
      RECT  265.69 242.2525 267.415 243.1175 ;
      RECT  87.8675 2.33 98.8925 2.745 ;
      RECT  99.3075 2.33 110.3325 2.745 ;
      RECT  122.1875 2.33 133.2125 2.745 ;
      RECT  133.6275 2.33 144.6525 2.745 ;
      RECT  350.9875 2.33 362.0125 2.745 ;
      RECT  362.4275 2.33 373.4525 2.745 ;
      RECT  53.83 0.275 239.0325 0.965 ;
      RECT  239.0325 0.275 239.4475 0.965 ;
      RECT  239.4475 0.275 407.84 0.965 ;
      RECT  225.0075 34.2375 225.775 43.8975 ;
      RECT  225.0075 43.8975 225.775 44.3125 ;
      RECT  225.0075 44.3125 225.775 57.3525 ;
      RECT  226.19 34.2375 231.165 43.8975 ;
      RECT  226.19 43.8975 231.165 44.3125 ;
      RECT  36.67 2.745 41.45 43.8975 ;
      RECT  36.67 43.8975 41.45 44.3125 ;
      RECT  41.865 2.745 42.6325 43.8975 ;
      RECT  41.865 43.8975 42.6325 44.3125 ;
      RECT  41.865 44.3125 42.6325 60.3425 ;
      RECT  57.6125 25.975 206.4075 27.675 ;
      RECT  57.6125 28.025 206.4075 31.06 ;
      RECT  170.8075 0.14 181.8325 0.275 ;
      RECT  225.775 34.2375 226.19 34.9275 ;
      RECT  225.0075 57.7675 226.4 64.8275 ;
      RECT  225.0075 64.8275 226.4 65.2425 ;
      RECT  225.0075 65.2425 226.4 233.9375 ;
      RECT  226.4 65.2425 226.815 233.9375 ;
      RECT  226.815 57.7675 231.165 64.8275 ;
      RECT  226.815 64.8275 231.165 65.2425 ;
      RECT  226.815 65.2425 231.165 233.9375 ;
      RECT  388.1675 0.14 399.1925 0.275 ;
      RECT  399.6075 0.14 407.84 0.275 ;
      RECT  159.3675 0.14 170.3925 0.275 ;
      RECT  226.19 44.3125 226.4 52.8675 ;
      RECT  226.19 52.8675 226.4 53.2825 ;
      RECT  226.19 53.2825 226.4 57.3525 ;
      RECT  226.4 44.3125 226.815 52.8675 ;
      RECT  226.815 44.3125 231.165 52.8675 ;
      RECT  226.815 52.8675 231.165 53.2825 ;
      RECT  226.815 53.2825 231.165 57.3525 ;
      RECT  41.45 50.2925 41.865 60.3425 ;
      RECT  225.775 44.3125 226.19 46.8875 ;
      RECT  0.56 1.38 2.285 14.2575 ;
      RECT  0.56 14.2575 2.285 14.6725 ;
      RECT  0.56 14.6725 2.285 15.3625 ;
      RECT  2.285 1.38 2.7 14.2575 ;
      RECT  2.285 14.6725 2.7 15.3625 ;
      RECT  2.7 1.38 36.255 14.2575 ;
      RECT  2.7 14.2575 36.255 14.6725 ;
      RECT  2.7 14.6725 36.255 15.3625 ;
      RECT  273.7675 0.14 284.7925 0.275 ;
      RECT  239.4475 0.14 250.4725 0.275 ;
      RECT  228.0075 0.14 239.0325 0.275 ;
      RECT  41.45 44.3125 41.865 46.8875 ;
      RECT  41.45 47.3025 41.865 49.8775 ;
      RECT  342.4075 0.14 353.4325 0.275 ;
      RECT  285.2075 0.14 296.2325 0.275 ;
      RECT  296.6475 0.14 307.6725 0.275 ;
      RECT  57.6125 230.39 60.7975 232.045 ;
      RECT  57.6125 232.395 60.7975 233.9375 ;
      RECT  60.7975 230.39 61.2125 232.045 ;
      RECT  60.7975 232.395 61.2125 233.9375 ;
      RECT  61.2125 230.39 206.4075 232.045 ;
      RECT  61.2125 232.395 206.4075 233.9375 ;
      RECT  206.4075 230.39 206.4425 232.045 ;
      RECT  206.4075 232.395 206.4425 233.9375 ;
      RECT  206.4425 230.39 208.0525 232.045 ;
      RECT  206.4425 232.045 208.0525 232.395 ;
      RECT  206.4425 232.395 208.0525 233.9375 ;
      RECT  36.67 44.3125 40.825 55.8575 ;
      RECT  36.67 55.8575 40.825 56.2725 ;
      RECT  36.67 56.2725 40.825 60.3425 ;
      RECT  41.24 44.3125 41.45 55.8575 ;
      RECT  41.24 55.8575 41.45 56.2725 ;
      RECT  41.24 56.2725 41.45 60.3425 ;
      RECT  226.4 53.2825 226.815 55.8575 ;
      RECT  226.4 56.2725 226.815 57.3525 ;
      RECT  206.4625 2.745 206.8775 22.8375 ;
      RECT  206.4625 23.2525 206.8775 24.6575 ;
      RECT  226.4 62.2525 226.815 64.8275 ;
      RECT  330.9675 0.14 341.9925 0.275 ;
      RECT  250.8875 0.14 261.9125 0.275 ;
      RECT  262.3275 0.14 273.3525 0.275 ;
      RECT  376.7275 0.14 387.7525 0.275 ;
      RECT  113.6075 0.14 124.6325 0.275 ;
      RECT  125.0475 0.14 136.0725 0.275 ;
      RECT  136.4875 0.14 147.5125 0.275 ;
      RECT  147.9275 0.14 158.9525 0.275 ;
      RECT  0.14 0.14 44.5525 0.275 ;
      RECT  0.14 0.275 44.5525 0.965 ;
      RECT  44.5525 0.275 44.9675 0.965 ;
      RECT  44.9675 0.14 53.415 0.275 ;
      RECT  44.9675 0.275 53.415 0.965 ;
      RECT  182.2475 0.14 193.2725 0.275 ;
      RECT  193.6875 0.14 204.7125 0.275 ;
      RECT  205.1275 0.14 216.1525 0.275 ;
      RECT  216.5675 0.14 227.5925 0.275 ;
      RECT  225.775 35.3425 226.19 37.9175 ;
      RECT  226.4 57.7675 226.815 58.8475 ;
      RECT  226.4 59.2625 226.815 61.8375 ;
      RECT  41.45 2.745 41.865 34.9275 ;
      RECT  41.45 35.3425 41.865 37.9175 ;
      RECT  53.83 0.14 55.9925 0.275 ;
      RECT  56.4075 0.14 67.4325 0.275 ;
      RECT  67.8475 0.14 78.8725 0.275 ;
      RECT  79.2875 0.14 90.3125 0.275 ;
      RECT  353.8475 0.14 364.8725 0.275 ;
      RECT  365.2875 0.14 376.3125 0.275 ;
      RECT  57.4775 1.38 57.6125 22.8375 ;
      RECT  57.4775 23.2525 57.6125 24.6575 ;
      RECT  57.6125 2.745 57.8925 22.8375 ;
      RECT  57.6125 23.2525 57.8925 24.6575 ;
      RECT  225.775 38.3325 226.19 40.9075 ;
      RECT  225.775 41.3225 226.19 43.8975 ;
      RECT  36.67 60.7575 40.825 64.8275 ;
      RECT  36.67 64.8275 40.825 65.2425 ;
      RECT  36.67 65.2425 40.825 65.9325 ;
      RECT  40.825 65.2425 41.24 65.9325 ;
      RECT  41.24 60.7575 42.6325 64.8275 ;
      RECT  41.24 64.8275 42.6325 65.2425 ;
      RECT  41.24 65.2425 42.6325 65.9325 ;
      RECT  225.775 47.3025 226.19 49.8775 ;
      RECT  225.775 50.2925 226.19 57.3525 ;
      RECT  40.825 56.2725 41.24 58.8475 ;
      RECT  40.825 59.2625 41.24 60.3425 ;
      RECT  308.0875 0.14 319.1125 0.275 ;
      RECT  319.5275 0.14 330.5525 0.275 ;
      RECT  41.45 38.3325 41.865 40.9075 ;
      RECT  41.45 41.3225 41.865 43.8975 ;
      RECT  40.825 44.3125 41.24 52.8675 ;
      RECT  40.825 53.2825 41.24 55.8575 ;
      RECT  90.7275 0.14 101.7525 0.275 ;
      RECT  102.1675 0.14 113.1925 0.275 ;
      RECT  231.58 243.6175 265.275 244.3075 ;
      RECT  231.58 244.3075 265.275 244.445 ;
      RECT  265.275 243.6175 265.69 244.3075 ;
      RECT  265.69 243.6175 267.415 244.3075 ;
      RECT  265.69 244.3075 267.415 244.445 ;
      RECT  40.825 60.7575 41.24 61.8375 ;
      RECT  40.825 62.2525 41.24 64.8275 ;
   LAYER  metal4 ;
      RECT  56.325 0.14 57.025 34.785 ;
      RECT  56.325 226.845 57.025 244.445 ;
      RECT  266.8675 34.785 267.5675 212.055 ;
      RECT  267.5675 34.785 407.84 212.055 ;
      RECT  267.5675 212.055 407.84 226.845 ;
      RECT  266.8675 235.0175 267.5675 244.445 ;
      RECT  267.5675 226.845 407.84 235.0175 ;
      RECT  267.5675 235.0175 407.84 244.445 ;
      RECT  57.025 0.14 231.305 17.43 ;
      RECT  231.305 0.14 232.005 17.43 ;
      RECT  232.005 0.14 407.84 17.43 ;
      RECT  232.005 17.43 407.84 34.785 ;
      RECT  231.305 35.485 232.005 212.055 ;
      RECT  232.005 34.785 266.8675 35.485 ;
      RECT  57.025 229.765 209.535 235.0175 ;
      RECT  209.535 229.765 210.235 235.0175 ;
      RECT  57.025 17.43 209.535 31.615 ;
      RECT  209.535 17.43 210.235 31.615 ;
      RECT  210.235 212.055 210.615 226.845 ;
      RECT  210.235 34.785 210.615 35.485 ;
      RECT  210.235 35.485 210.615 212.055 ;
      RECT  210.235 226.915 217.99 229.765 ;
      RECT  217.99 226.915 218.69 229.765 ;
      RECT  0.14 0.14 0.4075 23.9625 ;
      RECT  0.14 23.9625 0.4075 34.785 ;
      RECT  0.4075 0.14 1.1075 23.9625 ;
      RECT  0.14 34.785 0.4075 46.925 ;
      RECT  0.14 46.925 0.4075 226.845 ;
      RECT  0.4075 46.925 1.1075 226.845 ;
      RECT  38.55 0.14 39.25 16.585 ;
      RECT  39.25 0.14 56.325 16.585 ;
      RECT  39.25 16.585 56.325 23.9625 ;
      RECT  38.55 32.105 39.25 34.785 ;
      RECT  39.25 23.9625 56.325 32.105 ;
      RECT  57.025 235.0175 228.585 242.395 ;
      RECT  57.025 242.395 228.585 244.445 ;
      RECT  228.585 242.395 229.285 244.445 ;
      RECT  210.235 229.765 228.585 231.815 ;
      RECT  210.235 231.815 228.585 235.0175 ;
      RECT  228.585 229.765 229.285 231.815 ;
      RECT  57.025 226.845 57.405 229.765 ;
      RECT  57.025 31.615 57.405 34.785 ;
      RECT  57.025 212.055 57.405 226.845 ;
      RECT  57.025 34.785 57.405 35.485 ;
      RECT  57.025 35.485 57.405 212.055 ;
      RECT  0.14 226.915 48.95 244.445 ;
      RECT  48.95 226.915 49.65 244.445 ;
      RECT  49.65 226.915 56.325 244.445 ;
      RECT  1.1075 64.685 35.83 82.74 ;
      RECT  1.1075 82.74 35.83 226.845 ;
      RECT  35.83 46.925 36.53 64.685 ;
      RECT  35.83 82.74 36.53 226.845 ;
      RECT  232.005 35.485 264.805 212.0225 ;
      RECT  232.005 212.0225 264.805 212.055 ;
      RECT  264.805 35.485 265.505 212.0225 ;
      RECT  265.505 35.485 266.8675 212.0225 ;
      RECT  265.505 212.0225 266.8675 212.055 ;
      RECT  265.505 212.055 266.8675 226.845 ;
      RECT  265.505 226.845 266.8675 226.915 ;
      RECT  265.505 226.915 266.8675 229.765 ;
      RECT  265.505 229.765 266.8675 231.815 ;
      RECT  264.805 234.985 265.505 235.0175 ;
      RECT  265.505 231.815 266.8675 234.985 ;
      RECT  265.505 234.985 266.8675 235.0175 ;
      RECT  1.1075 0.14 5.825 14.115 ;
      RECT  1.1075 14.115 5.825 16.585 ;
      RECT  5.825 0.14 6.525 14.115 ;
      RECT  6.525 0.14 38.55 14.115 ;
      RECT  6.525 14.115 38.55 16.585 ;
      RECT  1.1075 16.585 5.825 23.9625 ;
      RECT  6.525 16.585 38.55 23.9625 ;
      RECT  5.825 29.635 6.525 32.105 ;
      RECT  6.525 23.9625 38.55 29.635 ;
      RECT  6.525 29.635 38.55 32.105 ;
      RECT  39.25 32.105 49.51 34.7525 ;
      RECT  49.51 32.105 50.21 34.7525 ;
      RECT  50.21 32.105 56.325 34.7525 ;
      RECT  50.21 34.7525 56.325 34.785 ;
      RECT  49.65 226.8775 50.21 226.915 ;
      RECT  50.21 226.845 56.325 226.8775 ;
      RECT  50.21 226.8775 56.325 226.915 ;
      RECT  50.21 34.785 56.325 46.925 ;
      RECT  50.21 46.925 56.325 226.845 ;
      RECT  210.235 31.615 217.43 34.7525 ;
      RECT  210.235 34.7525 217.43 34.785 ;
      RECT  217.43 31.615 218.13 34.7525 ;
      RECT  211.315 212.055 217.43 226.845 ;
      RECT  211.315 34.785 217.43 35.485 ;
      RECT  211.315 35.485 217.43 212.055 ;
      RECT  210.235 226.845 217.43 226.8775 ;
      RECT  210.235 226.8775 217.43 226.915 ;
      RECT  217.43 226.8775 217.99 226.915 ;
      RECT  58.565 226.845 209.075 229.765 ;
      RECT  58.565 31.615 209.075 34.785 ;
      RECT  58.565 212.055 209.075 226.845 ;
      RECT  58.565 34.785 209.075 35.485 ;
      RECT  58.565 35.485 209.075 212.055 ;
      RECT  229.285 235.0175 261.31 242.395 ;
      RECT  262.01 235.0175 266.8675 242.395 ;
      RECT  229.285 242.395 261.31 244.445 ;
      RECT  262.01 242.395 266.8675 244.445 ;
      RECT  218.69 226.915 261.31 229.345 ;
      RECT  218.69 229.345 261.31 229.765 ;
      RECT  261.31 226.915 262.01 229.345 ;
      RECT  262.01 226.915 264.805 229.345 ;
      RECT  262.01 229.345 264.805 229.765 ;
      RECT  229.285 229.765 261.31 231.815 ;
      RECT  262.01 229.765 264.805 231.815 ;
      RECT  229.285 231.815 261.31 234.985 ;
      RECT  262.01 231.815 264.805 234.985 ;
      RECT  229.285 234.985 261.31 235.0175 ;
      RECT  262.01 234.985 264.805 235.0175 ;
      RECT  218.69 34.785 219.925 35.485 ;
      RECT  218.69 35.485 219.925 212.055 ;
      RECT  218.69 212.055 219.925 226.845 ;
      RECT  220.625 212.055 264.805 226.845 ;
      RECT  218.69 226.845 219.925 226.915 ;
      RECT  220.625 226.845 264.805 226.915 ;
      RECT  218.13 34.7525 219.925 34.785 ;
      RECT  210.235 17.43 228.445 17.495 ;
      RECT  210.235 17.495 228.445 31.615 ;
      RECT  228.445 17.43 229.145 17.495 ;
      RECT  229.145 17.43 231.305 17.495 ;
      RECT  229.145 17.495 231.305 31.615 ;
      RECT  218.13 31.615 228.445 34.7525 ;
      RECT  229.145 31.615 231.305 34.7525 ;
      RECT  220.625 34.785 228.445 35.485 ;
      RECT  229.145 34.785 231.305 35.485 ;
      RECT  220.625 35.485 228.445 35.55 ;
      RECT  220.625 35.55 228.445 212.055 ;
      RECT  228.445 35.55 229.145 212.055 ;
      RECT  229.145 35.485 231.305 35.55 ;
      RECT  229.145 35.55 231.305 212.055 ;
      RECT  220.625 34.7525 228.445 34.785 ;
      RECT  229.145 34.7525 231.305 34.785 ;
      RECT  36.53 46.925 38.69 64.62 ;
      RECT  36.53 64.62 38.69 64.685 ;
      RECT  38.69 46.925 39.39 64.62 ;
      RECT  36.53 64.685 38.69 82.675 ;
      RECT  36.53 82.675 38.69 82.74 ;
      RECT  38.69 82.675 39.39 82.74 ;
      RECT  0.14 226.845 47.015 226.915 ;
      RECT  47.715 226.845 48.95 226.915 ;
      RECT  47.715 34.785 48.95 46.925 ;
      RECT  36.53 82.74 47.015 226.845 ;
      RECT  47.715 82.74 48.95 226.845 ;
      RECT  39.25 34.7525 47.015 34.785 ;
      RECT  47.715 34.7525 49.51 34.785 ;
      RECT  39.39 46.925 47.015 64.62 ;
      RECT  47.715 46.925 48.95 64.62 ;
      RECT  39.39 64.62 47.015 64.685 ;
      RECT  47.715 64.62 48.95 64.685 ;
      RECT  39.39 64.685 47.015 82.675 ;
      RECT  47.715 64.685 48.95 82.675 ;
      RECT  39.39 82.675 47.015 82.74 ;
      RECT  47.715 82.675 48.95 82.74 ;
      RECT  1.1075 32.105 2.47 34.785 ;
      RECT  3.17 32.105 38.55 34.785 ;
      RECT  1.1075 46.925 2.47 46.9575 ;
      RECT  1.1075 46.9575 2.47 64.685 ;
      RECT  2.47 46.9575 3.17 64.685 ;
      RECT  3.17 46.925 35.83 46.9575 ;
      RECT  3.17 46.9575 35.83 64.685 ;
      RECT  1.1075 23.9625 2.47 23.995 ;
      RECT  1.1075 23.995 2.47 29.635 ;
      RECT  2.47 23.9625 3.17 23.995 ;
      RECT  3.17 23.9625 5.825 23.995 ;
      RECT  3.17 23.995 5.825 29.635 ;
      RECT  1.1075 29.635 2.47 32.105 ;
      RECT  3.17 29.635 5.825 32.105 ;
      RECT  1.1075 34.785 2.47 46.925 ;
      RECT  3.17 34.785 47.015 46.925 ;
   END
END    freepdk45_sram_1w1r_128x124_31
END    LIBRARY
