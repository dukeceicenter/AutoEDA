../macros/freepdk45_sram_1rw0r_512x45/freepdk45_sram_1rw0r_512x45.lef