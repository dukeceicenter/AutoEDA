VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_256x48_12
   CLASS BLOCK ;
   SIZE 200.425 BY 230.19 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.465 1.1075 40.6 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.325 1.1075 43.46 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.185 1.1075 46.32 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.045 1.1075 49.18 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.905 1.1075 52.04 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.765 1.1075 54.9 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.625 1.1075 57.76 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.485 1.1075 60.62 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.345 1.1075 63.48 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.205 1.1075 66.34 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.065 1.1075 69.2 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.925 1.1075 72.06 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.785 1.1075 74.92 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.645 1.1075 77.78 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.505 1.1075 80.64 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.365 1.1075 83.5 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.225 1.1075 86.36 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.085 1.1075 89.22 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.945 1.1075 92.08 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.805 1.1075 94.94 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.665 1.1075 97.8 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.525 1.1075 100.66 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.385 1.1075 103.52 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.245 1.1075 106.38 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.105 1.1075 109.24 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.965 1.1075 112.1 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.825 1.1075 114.96 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.685 1.1075 117.82 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.545 1.1075 120.68 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.405 1.1075 123.54 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.265 1.1075 126.4 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.125 1.1075 129.26 1.2425 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.985 1.1075 132.12 1.2425 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.845 1.1075 134.98 1.2425 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.705 1.1075 137.84 1.2425 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.565 1.1075 140.7 1.2425 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.425 1.1075 143.56 1.2425 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.285 1.1075 146.42 1.2425 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.145 1.1075 149.28 1.2425 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.005 1.1075 152.14 1.2425 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.865 1.1075 155.0 1.2425 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.725 1.1075 157.86 1.2425 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.585 1.1075 160.72 1.2425 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.445 1.1075 163.58 1.2425 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.305 1.1075 166.44 1.2425 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.165 1.1075 169.3 1.2425 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.025 1.1075 172.16 1.2425 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.885 1.1075 175.02 1.2425 ;
      END
   END din0[47]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.165 1.1075 26.3 1.2425 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.445 51.6775 20.58 51.8125 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.445 54.4075 20.58 54.5425 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.445 56.6175 20.58 56.7525 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.445 59.3475 20.58 59.4825 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.445 61.5575 20.58 61.6925 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.445 64.2875 20.58 64.4225 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.445 66.4975 20.58 66.6325 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.125 227.615 171.26 227.75 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.705 19.5675 179.84 19.7025 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.705 16.8375 179.84 16.9725 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.705 14.6275 179.84 14.7625 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.705 11.8975 179.84 12.0325 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.705 9.6875 179.84 9.8225 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.705 6.9575 179.84 7.0925 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.705 4.7475 179.84 4.8825 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.005 228.9475 200.14 229.0825 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.9025 228.8625 194.0375 228.9975 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.025 1.1075 29.16 1.2425 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.885 1.1075 32.02 1.2425 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.745 1.1075 34.88 1.2425 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.605 1.1075 37.74 1.2425 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.6125 225.1925 43.7475 225.3275 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.9625 225.1925 46.0975 225.3275 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.3125 225.1925 48.4475 225.3275 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.6625 225.1925 50.7975 225.3275 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.0125 225.1925 53.1475 225.3275 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.3625 225.1925 55.4975 225.3275 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.7125 225.1925 57.8475 225.3275 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.0625 225.1925 60.1975 225.3275 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.4125 225.1925 62.5475 225.3275 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.7625 225.1925 64.8975 225.3275 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.1125 225.1925 67.2475 225.3275 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.4625 225.1925 69.5975 225.3275 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.8125 225.1925 71.9475 225.3275 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.1625 225.1925 74.2975 225.3275 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.5125 225.1925 76.6475 225.3275 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.8625 225.1925 78.9975 225.3275 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.2125 225.1925 81.3475 225.3275 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.5625 225.1925 83.6975 225.3275 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.9125 225.1925 86.0475 225.3275 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.2625 225.1925 88.3975 225.3275 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.6125 225.1925 90.7475 225.3275 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.9625 225.1925 93.0975 225.3275 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.3125 225.1925 95.4475 225.3275 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.6625 225.1925 97.7975 225.3275 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.0125 225.1925 100.1475 225.3275 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.3625 225.1925 102.4975 225.3275 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.7125 225.1925 104.8475 225.3275 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.0625 225.1925 107.1975 225.3275 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.4125 225.1925 109.5475 225.3275 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.7625 225.1925 111.8975 225.3275 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.1125 225.1925 114.2475 225.3275 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.4625 225.1925 116.5975 225.3275 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.8125 225.1925 118.9475 225.3275 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.1625 225.1925 121.2975 225.3275 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.5125 225.1925 123.6475 225.3275 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.8625 225.1925 125.9975 225.3275 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.2125 225.1925 128.3475 225.3275 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.5625 225.1925 130.6975 225.3275 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.9125 225.1925 133.0475 225.3275 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.2625 225.1925 135.3975 225.3275 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.6125 225.1925 137.7475 225.3275 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.9625 225.1925 140.0975 225.3275 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.3125 225.1925 142.4475 225.3275 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.6625 225.1925 144.7975 225.3275 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.0125 225.1925 147.1475 225.3275 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.3625 225.1925 149.4975 225.3275 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.7125 225.1925 151.8475 225.3275 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.0625 225.1925 154.1975 225.3275 ;
      END
   END dout1[47]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  28.7425 2.4725 28.8775 2.6075 ;
         LAYER metal3 ;
         RECT  156.3775 7.4475 156.5125 7.5825 ;
         LAYER metal3 ;
         RECT  173.1325 43.0975 173.2675 43.2325 ;
         LAYER metal4 ;
         RECT  33.28 20.67 33.42 212.24 ;
         LAYER metal3 ;
         RECT  85.9425 2.4725 86.0775 2.6075 ;
         LAYER metal3 ;
         RECT  166.0225 2.4725 166.1575 2.6075 ;
         LAYER metal4 ;
         RECT  179.985 3.315 180.125 20.81 ;
         LAYER metal4 ;
         RECT  20.16 50.57 20.3 68.065 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal3 ;
         RECT  166.055 212.74 166.19 212.875 ;
         LAYER metal3 ;
         RECT  39.2825 19.1775 39.4175 19.3125 ;
         LAYER metal4 ;
         RECT  39.28 20.67 39.42 212.17 ;
         LAYER metal3 ;
         RECT  31.99 11.9075 32.125 12.0425 ;
         LAYER metal3 ;
         RECT  172.7875 31.1375 172.9225 31.2725 ;
         LAYER metal4 ;
         RECT  177.265 217.7 177.405 227.72 ;
         LAYER metal3 ;
         RECT  51.6225 2.4725 51.7575 2.6075 ;
         LAYER metal3 ;
         RECT  131.7025 2.4725 131.8375 2.6075 ;
         LAYER metal3 ;
         RECT  26.8225 46.0875 26.9575 46.2225 ;
         LAYER metal3 ;
         RECT  74.5025 2.4725 74.6375 2.6075 ;
         LAYER metal3 ;
         RECT  40.4275 8.415 154.8675 8.485 ;
         LAYER metal4 ;
         RECT  40.36 17.5 40.5 215.09 ;
         LAYER metal3 ;
         RECT  171.4075 226.25 171.5425 226.385 ;
         LAYER metal3 ;
         RECT  154.5825 2.4725 154.7175 2.6075 ;
         LAYER metal3 ;
         RECT  40.4275 215.785 157.6875 215.855 ;
         LAYER metal3 ;
         RECT  40.1825 2.4725 40.3175 2.6075 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
         LAYER metal4 ;
         RECT  160.67 20.67 160.81 212.17 ;
         LAYER metal3 ;
         RECT  27.1675 22.1675 27.3025 22.3025 ;
         LAYER metal3 ;
         RECT  26.8225 43.0975 26.9575 43.2325 ;
         LAYER metal4 ;
         RECT  159.59 17.5 159.73 215.09 ;
         LAYER metal3 ;
         RECT  40.4275 16.805 156.5125 16.875 ;
         LAYER metal3 ;
         RECT  160.6725 213.5275 160.8075 213.6625 ;
         LAYER metal4 ;
         RECT  199.5975 197.94 199.7375 220.3425 ;
         LAYER metal4 ;
         RECT  166.67 20.67 166.81 212.24 ;
         LAYER metal3 ;
         RECT  172.7875 25.1575 172.9225 25.2925 ;
         LAYER metal3 ;
         RECT  27.1675 34.1275 27.3025 34.2625 ;
         LAYER metal4 ;
         RECT  22.88 2.47 23.02 17.43 ;
         LAYER metal3 ;
         RECT  25.8825 2.4725 26.0175 2.6075 ;
         LAYER metal3 ;
         RECT  120.2625 2.4725 120.3975 2.6075 ;
         LAYER metal3 ;
         RECT  173.1325 46.0875 173.2675 46.2225 ;
         LAYER metal3 ;
         RECT  172.7875 22.1675 172.9225 22.3025 ;
         LAYER metal3 ;
         RECT  27.1675 31.1375 27.3025 31.2725 ;
         LAYER metal3 ;
         RECT  27.1675 25.1575 27.3025 25.2925 ;
         LAYER metal3 ;
         RECT  172.7875 34.1275 172.9225 34.2625 ;
         LAYER metal3 ;
         RECT  173.1325 40.1075 173.2675 40.2425 ;
         LAYER metal3 ;
         RECT  197.865 227.5825 198.0 227.7175 ;
         LAYER metal3 ;
         RECT  40.4275 222.6375 154.8675 222.7075 ;
         LAYER metal3 ;
         RECT  40.2925 7.4475 40.4275 7.5825 ;
         LAYER metal3 ;
         RECT  26.8225 49.0775 26.9575 49.2125 ;
         LAYER metal3 ;
         RECT  97.3825 2.4725 97.5175 2.6075 ;
         LAYER metal3 ;
         RECT  143.1425 2.4725 143.2775 2.6075 ;
         LAYER metal3 ;
         RECT  173.1325 49.0775 173.2675 49.2125 ;
         LAYER metal3 ;
         RECT  167.965 220.6175 168.1 220.7525 ;
         LAYER metal3 ;
         RECT  26.8225 40.1075 26.9575 40.2425 ;
         LAYER metal3 ;
         RECT  33.9 19.965 34.035 20.1 ;
         LAYER metal3 ;
         RECT  63.0625 2.4725 63.1975 2.6075 ;
         LAYER metal3 ;
         RECT  108.8225 2.4725 108.9575 2.6075 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  25.015 44.5925 25.15 44.7275 ;
         LAYER metal4 ;
         RECT  23.02 50.505 23.16 68.0 ;
         LAYER metal3 ;
         RECT  111.6825 0.0025 111.8175 0.1375 ;
         LAYER metal3 ;
         RECT  174.94 47.5825 175.075 47.7175 ;
         LAYER metal3 ;
         RECT  100.2425 0.0025 100.3775 0.1375 ;
         LAYER metal3 ;
         RECT  31.99 9.4375 32.125 9.5725 ;
         LAYER metal3 ;
         RECT  40.2925 5.6275 40.4275 5.7625 ;
         LAYER metal3 ;
         RECT  54.4825 0.0025 54.6175 0.1375 ;
         LAYER metal3 ;
         RECT  40.4275 218.405 156.545 218.475 ;
         LAYER metal3 ;
         RECT  25.015 38.6125 25.15 38.7475 ;
         LAYER metal3 ;
         RECT  40.4275 220.745 154.9025 220.815 ;
         LAYER metal3 ;
         RECT  25.64 20.6725 25.775 20.8075 ;
         LAYER metal3 ;
         RECT  167.965 218.1475 168.1 218.2825 ;
         LAYER metal3 ;
         RECT  25.015 47.5825 25.15 47.7175 ;
         LAYER metal3 ;
         RECT  174.315 26.6525 174.45 26.7875 ;
         LAYER metal4 ;
         RECT  177.125 3.38 177.265 20.875 ;
         LAYER metal3 ;
         RECT  25.64 26.6525 25.775 26.7875 ;
         LAYER metal4 ;
         RECT  166.11 20.6375 166.25 212.2025 ;
         LAYER metal3 ;
         RECT  168.8825 0.0025 169.0175 0.1375 ;
         LAYER metal4 ;
         RECT  194.04 215.23 194.18 230.19 ;
         LAYER metal3 ;
         RECT  174.94 38.6125 175.075 38.7475 ;
         LAYER metal3 ;
         RECT  40.4275 14.185 156.545 14.255 ;
         LAYER metal3 ;
         RECT  77.3625 0.0025 77.4975 0.1375 ;
         LAYER metal3 ;
         RECT  174.315 32.6325 174.45 32.7675 ;
         LAYER metal4 ;
         RECT  31.345 20.6375 31.485 212.24 ;
         LAYER metal3 ;
         RECT  156.3775 5.6275 156.5125 5.7625 ;
         LAYER metal3 ;
         RECT  25.64 32.6325 25.775 32.7675 ;
         LAYER metal4 ;
         RECT  40.82 17.5 40.96 215.09 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal3 ;
         RECT  25.64 23.6625 25.775 23.7975 ;
         LAYER metal3 ;
         RECT  123.1225 0.0025 123.2575 0.1375 ;
         LAYER metal3 ;
         RECT  31.99 14.3775 32.125 14.5125 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal3 ;
         RECT  25.64 35.6225 25.775 35.7575 ;
         LAYER metal3 ;
         RECT  174.94 44.5925 175.075 44.7275 ;
         LAYER metal3 ;
         RECT  25.015 41.6025 25.15 41.7375 ;
         LAYER metal3 ;
         RECT  174.315 29.6425 174.45 29.7775 ;
         LAYER metal3 ;
         RECT  197.865 230.0525 198.0 230.1875 ;
         LAYER metal3 ;
         RECT  28.7425 0.0025 28.8775 0.1375 ;
         LAYER metal3 ;
         RECT  40.4275 10.465 154.8675 10.535 ;
         LAYER metal3 ;
         RECT  168.5475 228.72 168.6825 228.855 ;
         LAYER metal4 ;
         RECT  197.535 197.9075 197.675 220.31 ;
         LAYER metal3 ;
         RECT  31.6025 0.0025 31.7375 0.1375 ;
         LAYER metal3 ;
         RECT  146.0025 0.0025 146.1375 0.1375 ;
         LAYER metal3 ;
         RECT  65.9225 0.0025 66.0575 0.1375 ;
         LAYER metal3 ;
         RECT  157.4425 0.0025 157.5775 0.1375 ;
         LAYER metal3 ;
         RECT  134.5625 0.0025 134.6975 0.1375 ;
         LAYER metal3 ;
         RECT  174.315 35.6225 174.45 35.7575 ;
         LAYER metal3 ;
         RECT  174.94 41.6025 175.075 41.7375 ;
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal3 ;
         RECT  167.965 223.0875 168.1 223.2225 ;
         LAYER metal3 ;
         RECT  174.315 20.6725 174.45 20.8075 ;
         LAYER metal4 ;
         RECT  168.605 20.6375 168.745 212.24 ;
         LAYER metal3 ;
         RECT  174.94 50.5725 175.075 50.7075 ;
         LAYER metal3 ;
         RECT  25.64 29.6425 25.775 29.7775 ;
         LAYER metal3 ;
         RECT  43.0425 0.0025 43.1775 0.1375 ;
         LAYER metal4 ;
         RECT  159.13 17.5 159.27 215.09 ;
         LAYER metal3 ;
         RECT  88.8025 0.0025 88.9375 0.1375 ;
         LAYER metal3 ;
         RECT  25.015 50.5725 25.15 50.7075 ;
         LAYER metal3 ;
         RECT  174.315 23.6625 174.45 23.7975 ;
         LAYER metal4 ;
         RECT  33.84 20.6375 33.98 212.2025 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 200.285 230.05 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 200.285 230.05 ;
   LAYER  metal3 ;
      RECT  40.325 0.14 40.74 0.9675 ;
      RECT  40.74 0.9675 43.185 1.3825 ;
      RECT  43.6 0.9675 46.045 1.3825 ;
      RECT  46.46 0.9675 48.905 1.3825 ;
      RECT  49.32 0.9675 51.765 1.3825 ;
      RECT  52.18 0.9675 54.625 1.3825 ;
      RECT  55.04 0.9675 57.485 1.3825 ;
      RECT  57.9 0.9675 60.345 1.3825 ;
      RECT  60.76 0.9675 63.205 1.3825 ;
      RECT  63.62 0.9675 66.065 1.3825 ;
      RECT  66.48 0.9675 68.925 1.3825 ;
      RECT  69.34 0.9675 71.785 1.3825 ;
      RECT  72.2 0.9675 74.645 1.3825 ;
      RECT  75.06 0.9675 77.505 1.3825 ;
      RECT  77.92 0.9675 80.365 1.3825 ;
      RECT  80.78 0.9675 83.225 1.3825 ;
      RECT  83.64 0.9675 86.085 1.3825 ;
      RECT  86.5 0.9675 88.945 1.3825 ;
      RECT  89.36 0.9675 91.805 1.3825 ;
      RECT  92.22 0.9675 94.665 1.3825 ;
      RECT  95.08 0.9675 97.525 1.3825 ;
      RECT  97.94 0.9675 100.385 1.3825 ;
      RECT  100.8 0.9675 103.245 1.3825 ;
      RECT  103.66 0.9675 106.105 1.3825 ;
      RECT  106.52 0.9675 108.965 1.3825 ;
      RECT  109.38 0.9675 111.825 1.3825 ;
      RECT  112.24 0.9675 114.685 1.3825 ;
      RECT  115.1 0.9675 117.545 1.3825 ;
      RECT  117.96 0.9675 120.405 1.3825 ;
      RECT  120.82 0.9675 123.265 1.3825 ;
      RECT  123.68 0.9675 126.125 1.3825 ;
      RECT  126.54 0.9675 128.985 1.3825 ;
      RECT  129.4 0.9675 131.845 1.3825 ;
      RECT  132.26 0.9675 134.705 1.3825 ;
      RECT  135.12 0.9675 137.565 1.3825 ;
      RECT  137.98 0.9675 140.425 1.3825 ;
      RECT  140.84 0.9675 143.285 1.3825 ;
      RECT  143.7 0.9675 146.145 1.3825 ;
      RECT  146.56 0.9675 149.005 1.3825 ;
      RECT  149.42 0.9675 151.865 1.3825 ;
      RECT  152.28 0.9675 154.725 1.3825 ;
      RECT  155.14 0.9675 157.585 1.3825 ;
      RECT  158.0 0.9675 160.445 1.3825 ;
      RECT  160.86 0.9675 163.305 1.3825 ;
      RECT  163.72 0.9675 166.165 1.3825 ;
      RECT  166.58 0.9675 169.025 1.3825 ;
      RECT  169.44 0.9675 171.885 1.3825 ;
      RECT  172.3 0.9675 174.745 1.3825 ;
      RECT  175.16 0.9675 200.285 1.3825 ;
      RECT  0.14 51.5375 20.305 51.9525 ;
      RECT  0.14 51.9525 20.305 230.05 ;
      RECT  20.305 1.3825 20.72 51.5375 ;
      RECT  20.72 51.5375 40.325 51.9525 ;
      RECT  20.305 51.9525 20.72 54.2675 ;
      RECT  20.305 54.6825 20.72 56.4775 ;
      RECT  20.305 56.8925 20.72 59.2075 ;
      RECT  20.305 59.6225 20.72 61.4175 ;
      RECT  20.305 61.8325 20.72 64.1475 ;
      RECT  20.305 64.5625 20.72 66.3575 ;
      RECT  20.305 66.7725 20.72 230.05 ;
      RECT  40.74 227.475 170.985 227.89 ;
      RECT  170.985 227.89 171.4 230.05 ;
      RECT  171.4 1.3825 179.565 19.4275 ;
      RECT  171.4 19.4275 179.565 19.8425 ;
      RECT  179.565 19.8425 179.98 227.475 ;
      RECT  179.98 1.3825 200.285 19.4275 ;
      RECT  179.98 19.4275 200.285 19.8425 ;
      RECT  179.565 17.1125 179.98 19.4275 ;
      RECT  179.565 14.9025 179.98 16.6975 ;
      RECT  179.565 12.1725 179.98 14.4875 ;
      RECT  179.565 9.9625 179.98 11.7575 ;
      RECT  179.565 7.2325 179.98 9.5475 ;
      RECT  179.565 1.3825 179.98 4.6075 ;
      RECT  179.565 5.0225 179.98 6.8175 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  199.865 227.89 200.28 228.8075 ;
      RECT  199.865 229.2225 200.28 230.05 ;
      RECT  200.28 227.89 200.285 228.8075 ;
      RECT  200.28 228.8075 200.285 229.2225 ;
      RECT  200.28 229.2225 200.285 230.05 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 51.5375 ;
      RECT  6.5225 1.3825 20.305 1.4675 ;
      RECT  6.5225 1.4675 20.305 51.5375 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 26.025 1.0525 ;
      RECT  6.5225 1.0525 26.025 1.3825 ;
      RECT  171.4 227.89 193.7625 228.7225 ;
      RECT  171.4 228.7225 193.7625 228.8075 ;
      RECT  193.7625 227.89 194.1775 228.7225 ;
      RECT  194.1775 227.89 199.865 228.7225 ;
      RECT  194.1775 228.7225 199.865 228.8075 ;
      RECT  171.4 228.8075 193.7625 229.1375 ;
      RECT  171.4 229.1375 193.7625 229.2225 ;
      RECT  193.7625 229.1375 194.1775 229.2225 ;
      RECT  194.1775 228.8075 199.865 229.1375 ;
      RECT  194.1775 229.1375 199.865 229.2225 ;
      RECT  26.44 0.9675 28.885 1.3825 ;
      RECT  29.3 0.9675 31.745 1.3825 ;
      RECT  32.16 0.9675 34.605 1.3825 ;
      RECT  35.02 0.9675 37.465 1.3825 ;
      RECT  37.88 0.9675 40.325 1.3825 ;
      RECT  40.74 225.0525 43.4725 225.4675 ;
      RECT  40.74 225.4675 43.4725 227.475 ;
      RECT  43.4725 225.4675 43.8875 227.475 ;
      RECT  43.8875 225.4675 170.985 227.475 ;
      RECT  43.8875 225.0525 45.8225 225.4675 ;
      RECT  46.2375 225.0525 48.1725 225.4675 ;
      RECT  48.5875 225.0525 50.5225 225.4675 ;
      RECT  50.9375 225.0525 52.8725 225.4675 ;
      RECT  53.2875 225.0525 55.2225 225.4675 ;
      RECT  55.6375 225.0525 57.5725 225.4675 ;
      RECT  57.9875 225.0525 59.9225 225.4675 ;
      RECT  60.3375 225.0525 62.2725 225.4675 ;
      RECT  62.6875 225.0525 64.6225 225.4675 ;
      RECT  65.0375 225.0525 66.9725 225.4675 ;
      RECT  67.3875 225.0525 69.3225 225.4675 ;
      RECT  69.7375 225.0525 71.6725 225.4675 ;
      RECT  72.0875 225.0525 74.0225 225.4675 ;
      RECT  74.4375 225.0525 76.3725 225.4675 ;
      RECT  76.7875 225.0525 78.7225 225.4675 ;
      RECT  79.1375 225.0525 81.0725 225.4675 ;
      RECT  81.4875 225.0525 83.4225 225.4675 ;
      RECT  83.8375 225.0525 85.7725 225.4675 ;
      RECT  86.1875 225.0525 88.1225 225.4675 ;
      RECT  88.5375 225.0525 90.4725 225.4675 ;
      RECT  90.8875 225.0525 92.8225 225.4675 ;
      RECT  93.2375 225.0525 95.1725 225.4675 ;
      RECT  95.5875 225.0525 97.5225 225.4675 ;
      RECT  97.9375 225.0525 99.8725 225.4675 ;
      RECT  100.2875 225.0525 102.2225 225.4675 ;
      RECT  102.6375 225.0525 104.5725 225.4675 ;
      RECT  104.9875 225.0525 106.9225 225.4675 ;
      RECT  107.3375 225.0525 109.2725 225.4675 ;
      RECT  109.6875 225.0525 111.6225 225.4675 ;
      RECT  112.0375 225.0525 113.9725 225.4675 ;
      RECT  114.3875 225.0525 116.3225 225.4675 ;
      RECT  116.7375 225.0525 118.6725 225.4675 ;
      RECT  119.0875 225.0525 121.0225 225.4675 ;
      RECT  121.4375 225.0525 123.3725 225.4675 ;
      RECT  123.7875 225.0525 125.7225 225.4675 ;
      RECT  126.1375 225.0525 128.0725 225.4675 ;
      RECT  128.4875 225.0525 130.4225 225.4675 ;
      RECT  130.8375 225.0525 132.7725 225.4675 ;
      RECT  133.1875 225.0525 135.1225 225.4675 ;
      RECT  135.5375 225.0525 137.4725 225.4675 ;
      RECT  137.8875 225.0525 139.8225 225.4675 ;
      RECT  140.2375 225.0525 142.1725 225.4675 ;
      RECT  142.5875 225.0525 144.5225 225.4675 ;
      RECT  144.9375 225.0525 146.8725 225.4675 ;
      RECT  147.2875 225.0525 149.2225 225.4675 ;
      RECT  149.6375 225.0525 151.5725 225.4675 ;
      RECT  151.9875 225.0525 153.9225 225.4675 ;
      RECT  154.3375 225.0525 170.985 225.4675 ;
      RECT  20.72 1.3825 28.6025 2.3325 ;
      RECT  28.6025 1.3825 29.0175 2.3325 ;
      RECT  28.6025 2.7475 29.0175 51.5375 ;
      RECT  29.0175 1.3825 40.325 2.3325 ;
      RECT  43.8875 7.3075 156.2375 7.7225 ;
      RECT  156.6525 7.3075 170.985 7.7225 ;
      RECT  171.4 42.9575 172.9925 43.3725 ;
      RECT  173.4075 42.9575 179.565 43.3725 ;
      RECT  43.8875 1.3825 85.8025 2.3325 ;
      RECT  43.8875 2.7475 85.8025 7.3075 ;
      RECT  85.8025 1.3825 86.2175 2.3325 ;
      RECT  85.8025 2.7475 86.2175 7.3075 ;
      RECT  86.2175 1.3825 156.2375 2.3325 ;
      RECT  86.2175 2.7475 156.2375 7.3075 ;
      RECT  156.6525 1.3825 165.8825 2.3325 ;
      RECT  156.6525 2.3325 165.8825 2.7475 ;
      RECT  156.6525 2.7475 165.8825 7.3075 ;
      RECT  165.8825 1.3825 166.2975 2.3325 ;
      RECT  165.8825 2.7475 166.2975 7.3075 ;
      RECT  166.2975 1.3825 170.985 2.3325 ;
      RECT  166.2975 2.3325 170.985 2.7475 ;
      RECT  166.2975 2.7475 170.985 7.3075 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 51.5375 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 51.5375 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 51.5375 ;
      RECT  156.6525 212.6 165.915 213.015 ;
      RECT  165.915 7.7225 166.33 212.6 ;
      RECT  165.915 213.015 166.33 225.0525 ;
      RECT  166.33 7.7225 170.985 212.6 ;
      RECT  166.33 212.6 170.985 213.015 ;
      RECT  29.0175 19.0375 39.1425 19.4525 ;
      RECT  39.1425 2.7475 39.5575 19.0375 ;
      RECT  39.1425 19.4525 39.5575 51.5375 ;
      RECT  39.5575 19.0375 40.325 19.4525 ;
      RECT  39.5575 19.4525 40.325 51.5375 ;
      RECT  29.0175 2.7475 31.85 11.7675 ;
      RECT  29.0175 11.7675 31.85 12.1825 ;
      RECT  29.0175 12.1825 31.85 19.0375 ;
      RECT  32.265 2.7475 39.1425 11.7675 ;
      RECT  32.265 11.7675 39.1425 12.1825 ;
      RECT  32.265 12.1825 39.1425 19.0375 ;
      RECT  171.4 19.8425 172.6475 30.9975 ;
      RECT  171.4 30.9975 172.6475 31.4125 ;
      RECT  171.4 31.4125 172.6475 42.9575 ;
      RECT  173.0625 19.8425 173.4075 30.9975 ;
      RECT  173.0625 30.9975 173.4075 31.4125 ;
      RECT  43.8875 2.3325 51.4825 2.7475 ;
      RECT  20.72 45.9475 26.6825 46.3625 ;
      RECT  27.0975 45.9475 28.6025 46.3625 ;
      RECT  27.0975 46.3625 28.6025 51.5375 ;
      RECT  74.7775 2.3325 85.8025 2.7475 ;
      RECT  40.74 1.3825 43.4725 8.275 ;
      RECT  43.4725 1.3825 43.8875 8.275 ;
      RECT  43.8875 7.7225 155.0075 8.275 ;
      RECT  155.0075 7.7225 156.2375 8.275 ;
      RECT  155.0075 8.275 156.2375 8.625 ;
      RECT  39.5575 8.275 40.2875 8.625 ;
      RECT  39.5575 8.625 40.2875 19.0375 ;
      RECT  170.985 1.3825 171.2675 226.11 ;
      RECT  170.985 226.11 171.2675 226.525 ;
      RECT  170.985 226.525 171.2675 227.475 ;
      RECT  171.2675 1.3825 171.4 226.11 ;
      RECT  171.2675 226.525 171.4 227.475 ;
      RECT  171.4 43.3725 171.6825 226.11 ;
      RECT  171.4 226.525 171.6825 227.475 ;
      RECT  171.6825 43.3725 172.9925 226.11 ;
      RECT  171.6825 226.11 172.9925 226.525 ;
      RECT  171.6825 226.525 172.9925 227.475 ;
      RECT  154.8575 2.3325 156.2375 2.7475 ;
      RECT  20.72 51.9525 40.2875 215.645 ;
      RECT  20.72 215.645 40.2875 215.995 ;
      RECT  20.72 215.995 40.2875 230.05 ;
      RECT  40.2875 51.9525 40.325 215.645 ;
      RECT  156.6525 213.015 157.8275 215.645 ;
      RECT  157.8275 215.645 165.915 215.995 ;
      RECT  157.8275 215.995 165.915 225.0525 ;
      RECT  29.0175 2.3325 40.0425 2.7475 ;
      RECT  40.325 1.3825 40.4575 2.3325 ;
      RECT  40.4575 1.3825 40.74 2.3325 ;
      RECT  40.4575 2.3325 40.74 2.7475 ;
      RECT  26.6825 2.7475 27.0275 22.0275 ;
      RECT  26.6825 22.0275 27.0275 22.4425 ;
      RECT  27.0275 2.7475 27.0975 22.0275 ;
      RECT  27.0975 2.7475 27.4425 22.0275 ;
      RECT  27.4425 2.7475 28.6025 22.0275 ;
      RECT  27.4425 22.0275 28.6025 22.4425 ;
      RECT  27.4425 22.4425 28.6025 45.9475 ;
      RECT  26.6825 43.3725 27.0275 45.9475 ;
      RECT  27.0275 43.3725 27.0975 45.9475 ;
      RECT  40.2875 17.015 40.325 19.0375 ;
      RECT  156.2375 17.015 156.6525 215.645 ;
      RECT  40.325 17.015 40.74 215.645 ;
      RECT  40.74 17.015 43.4725 215.645 ;
      RECT  43.4725 17.015 43.8875 215.645 ;
      RECT  43.8875 17.015 155.0075 215.645 ;
      RECT  155.0075 17.015 156.2375 215.645 ;
      RECT  157.8275 213.015 160.5325 213.3875 ;
      RECT  157.8275 213.3875 160.5325 213.8025 ;
      RECT  157.8275 213.8025 160.5325 215.645 ;
      RECT  160.5325 213.015 160.9475 213.3875 ;
      RECT  160.5325 213.8025 160.9475 215.645 ;
      RECT  160.9475 213.015 165.915 213.3875 ;
      RECT  160.9475 213.3875 165.915 213.8025 ;
      RECT  160.9475 213.8025 165.915 215.645 ;
      RECT  172.6475 25.4325 172.9925 30.9975 ;
      RECT  172.9925 25.4325 173.0625 30.9975 ;
      RECT  27.0975 34.4025 27.4425 45.9475 ;
      RECT  20.72 2.3325 25.7425 2.7475 ;
      RECT  26.1575 2.3325 28.6025 2.7475 ;
      RECT  120.5375 2.3325 131.5625 2.7475 ;
      RECT  172.9925 43.3725 173.4075 45.9475 ;
      RECT  172.6475 19.8425 172.9925 22.0275 ;
      RECT  172.6475 22.4425 172.9925 25.0175 ;
      RECT  172.9925 19.8425 173.0625 22.0275 ;
      RECT  172.9925 22.4425 173.0625 25.0175 ;
      RECT  27.0975 31.4125 27.4425 33.9875 ;
      RECT  27.0275 31.4125 27.0975 33.9875 ;
      RECT  27.0975 22.4425 27.4425 25.0175 ;
      RECT  27.0975 25.4325 27.4425 30.9975 ;
      RECT  27.0275 22.4425 27.0975 25.0175 ;
      RECT  27.0275 25.4325 27.0975 30.9975 ;
      RECT  172.6475 31.4125 172.9925 33.9875 ;
      RECT  172.6475 34.4025 172.9925 42.9575 ;
      RECT  172.9925 31.4125 173.0625 33.9875 ;
      RECT  173.0625 31.4125 173.4075 39.9675 ;
      RECT  173.0625 40.3825 173.4075 42.9575 ;
      RECT  172.9925 34.4025 173.0625 39.9675 ;
      RECT  172.9925 40.3825 173.0625 42.9575 ;
      RECT  171.4 227.475 197.725 227.8575 ;
      RECT  171.4 227.8575 197.725 227.89 ;
      RECT  197.725 227.8575 198.14 227.89 ;
      RECT  198.14 227.475 200.285 227.8575 ;
      RECT  198.14 227.8575 200.285 227.89 ;
      RECT  179.98 19.8425 197.725 227.4425 ;
      RECT  179.98 227.4425 197.725 227.475 ;
      RECT  197.725 19.8425 198.14 227.4425 ;
      RECT  198.14 19.8425 200.285 227.4425 ;
      RECT  198.14 227.4425 200.285 227.475 ;
      RECT  40.2875 222.8475 40.325 230.05 ;
      RECT  40.325 222.8475 40.74 230.05 ;
      RECT  40.74 222.8475 43.4725 225.0525 ;
      RECT  43.4725 222.8475 43.8875 225.0525 ;
      RECT  43.8875 222.8475 155.0075 225.0525 ;
      RECT  39.5575 2.7475 40.1525 7.3075 ;
      RECT  39.5575 7.3075 40.1525 7.7225 ;
      RECT  39.5575 7.7225 40.1525 8.275 ;
      RECT  40.1525 7.7225 40.2875 8.275 ;
      RECT  40.2875 7.7225 40.325 8.275 ;
      RECT  40.325 7.7225 40.4575 8.275 ;
      RECT  40.4575 7.7225 40.5675 8.275 ;
      RECT  40.5675 2.7475 40.74 7.3075 ;
      RECT  40.5675 7.3075 40.74 7.7225 ;
      RECT  40.5675 7.7225 40.74 8.275 ;
      RECT  26.6825 46.3625 27.0975 48.9375 ;
      RECT  26.6825 49.3525 27.0975 51.5375 ;
      RECT  86.2175 2.3325 97.2425 2.7475 ;
      RECT  131.9775 2.3325 143.0025 2.7475 ;
      RECT  143.4175 2.3325 154.4425 2.7475 ;
      RECT  172.9925 46.3625 173.4075 48.9375 ;
      RECT  172.9925 49.3525 173.4075 227.475 ;
      RECT  166.33 213.015 167.825 220.4775 ;
      RECT  166.33 220.4775 167.825 220.8925 ;
      RECT  166.33 220.8925 167.825 225.0525 ;
      RECT  168.24 213.015 170.985 220.4775 ;
      RECT  168.24 220.4775 170.985 220.8925 ;
      RECT  168.24 220.8925 170.985 225.0525 ;
      RECT  26.6825 22.4425 27.0275 39.9675 ;
      RECT  26.6825 40.3825 27.0275 42.9575 ;
      RECT  27.0275 34.4025 27.0975 39.9675 ;
      RECT  27.0275 40.3825 27.0975 42.9575 ;
      RECT  29.0175 19.4525 33.76 19.825 ;
      RECT  29.0175 19.825 33.76 20.24 ;
      RECT  29.0175 20.24 33.76 51.5375 ;
      RECT  33.76 19.4525 34.175 19.825 ;
      RECT  33.76 20.24 34.175 51.5375 ;
      RECT  34.175 19.4525 39.1425 19.825 ;
      RECT  34.175 19.825 39.1425 20.24 ;
      RECT  34.175 20.24 39.1425 51.5375 ;
      RECT  51.8975 2.3325 62.9225 2.7475 ;
      RECT  63.3375 2.3325 74.3625 2.7475 ;
      RECT  97.6575 2.3325 108.6825 2.7475 ;
      RECT  109.0975 2.3325 120.1225 2.7475 ;
      RECT  20.72 2.7475 24.875 44.4525 ;
      RECT  20.72 44.4525 24.875 44.8675 ;
      RECT  20.72 44.8675 24.875 45.9475 ;
      RECT  24.875 44.8675 25.29 45.9475 ;
      RECT  25.29 44.4525 26.6825 44.8675 ;
      RECT  25.29 44.8675 26.6825 45.9475 ;
      RECT  40.74 0.2775 111.5425 0.9675 ;
      RECT  111.5425 0.2775 111.9575 0.9675 ;
      RECT  111.9575 0.2775 200.285 0.9675 ;
      RECT  173.4075 43.3725 174.8 47.4425 ;
      RECT  173.4075 47.4425 174.8 47.8575 ;
      RECT  173.4075 47.8575 174.8 227.475 ;
      RECT  175.215 43.3725 179.565 47.4425 ;
      RECT  175.215 47.4425 179.565 47.8575 ;
      RECT  175.215 47.8575 179.565 227.475 ;
      RECT  100.5175 0.14 111.5425 0.2775 ;
      RECT  31.85 2.7475 32.265 9.2975 ;
      RECT  31.85 9.7125 32.265 11.7675 ;
      RECT  40.1525 2.7475 40.2875 5.4875 ;
      RECT  40.1525 5.9025 40.2875 7.3075 ;
      RECT  40.2875 2.7475 40.325 5.4875 ;
      RECT  40.2875 5.9025 40.325 7.3075 ;
      RECT  40.325 2.7475 40.4575 5.4875 ;
      RECT  40.325 5.9025 40.4575 7.3075 ;
      RECT  40.4575 2.7475 40.5675 5.4875 ;
      RECT  40.4575 5.9025 40.5675 7.3075 ;
      RECT  156.2375 215.995 156.6525 218.265 ;
      RECT  156.2375 218.615 156.6525 225.0525 ;
      RECT  156.6525 215.995 156.685 218.265 ;
      RECT  156.6525 218.615 156.685 225.0525 ;
      RECT  156.685 215.995 157.8275 218.265 ;
      RECT  156.685 218.265 157.8275 218.615 ;
      RECT  156.685 218.615 157.8275 225.0525 ;
      RECT  155.0075 215.995 156.2375 218.265 ;
      RECT  40.2875 215.995 40.325 218.265 ;
      RECT  40.325 215.995 40.74 218.265 ;
      RECT  40.74 215.995 43.4725 218.265 ;
      RECT  43.4725 215.995 43.8875 218.265 ;
      RECT  43.8875 215.995 155.0075 218.265 ;
      RECT  24.875 2.7475 25.29 38.4725 ;
      RECT  155.0075 218.615 155.0425 220.605 ;
      RECT  155.0075 220.955 155.0425 225.0525 ;
      RECT  155.0425 218.615 156.2375 220.605 ;
      RECT  155.0425 220.605 156.2375 220.955 ;
      RECT  155.0425 220.955 156.2375 225.0525 ;
      RECT  40.2875 218.615 40.325 220.605 ;
      RECT  40.2875 220.955 40.325 222.4975 ;
      RECT  40.325 218.615 40.74 220.605 ;
      RECT  40.325 220.955 40.74 222.4975 ;
      RECT  40.74 218.615 43.4725 220.605 ;
      RECT  40.74 220.955 43.4725 222.4975 ;
      RECT  43.4725 218.615 43.8875 220.605 ;
      RECT  43.4725 220.955 43.8875 222.4975 ;
      RECT  43.8875 218.615 155.0075 220.605 ;
      RECT  43.8875 220.955 155.0075 222.4975 ;
      RECT  25.29 2.7475 25.5 20.5325 ;
      RECT  25.29 20.5325 25.5 20.9475 ;
      RECT  25.29 20.9475 25.5 44.4525 ;
      RECT  25.5 2.7475 25.915 20.5325 ;
      RECT  25.915 2.7475 26.6825 20.5325 ;
      RECT  25.915 20.5325 26.6825 20.9475 ;
      RECT  25.915 20.9475 26.6825 44.4525 ;
      RECT  167.825 213.015 168.24 218.0075 ;
      RECT  167.825 218.4225 168.24 220.4775 ;
      RECT  20.72 46.3625 24.875 47.4425 ;
      RECT  20.72 47.4425 24.875 47.8575 ;
      RECT  20.72 47.8575 24.875 51.5375 ;
      RECT  24.875 46.3625 25.29 47.4425 ;
      RECT  25.29 46.3625 26.6825 47.4425 ;
      RECT  25.29 47.4425 26.6825 47.8575 ;
      RECT  25.29 47.8575 26.6825 51.5375 ;
      RECT  173.4075 19.8425 174.175 26.5125 ;
      RECT  173.4075 26.5125 174.175 26.9275 ;
      RECT  173.4075 26.9275 174.175 42.9575 ;
      RECT  174.59 19.8425 179.565 26.5125 ;
      RECT  174.59 26.5125 179.565 26.9275 ;
      RECT  169.1575 0.14 200.285 0.2775 ;
      RECT  174.59 26.9275 174.8 38.4725 ;
      RECT  174.59 38.4725 174.8 38.8875 ;
      RECT  174.59 38.8875 174.8 42.9575 ;
      RECT  174.8 26.9275 175.215 38.4725 ;
      RECT  175.215 26.9275 179.565 38.4725 ;
      RECT  175.215 38.4725 179.565 38.8875 ;
      RECT  175.215 38.8875 179.565 42.9575 ;
      RECT  156.6525 7.7225 156.685 14.045 ;
      RECT  156.6525 14.395 156.685 212.6 ;
      RECT  156.685 7.7225 165.915 14.045 ;
      RECT  156.685 14.045 165.915 14.395 ;
      RECT  156.685 14.395 165.915 212.6 ;
      RECT  40.2875 14.395 40.325 16.665 ;
      RECT  156.2375 7.7225 156.6525 14.045 ;
      RECT  156.2375 14.395 156.6525 16.665 ;
      RECT  40.325 14.395 40.74 16.665 ;
      RECT  40.74 14.395 43.4725 16.665 ;
      RECT  43.4725 14.395 43.8875 16.665 ;
      RECT  43.8875 14.395 155.0075 16.665 ;
      RECT  155.0075 8.625 156.2375 14.045 ;
      RECT  155.0075 14.395 156.2375 16.665 ;
      RECT  156.2375 1.3825 156.6525 5.4875 ;
      RECT  156.2375 5.9025 156.6525 7.3075 ;
      RECT  25.5 20.9475 25.915 23.5225 ;
      RECT  25.5 23.9375 25.915 26.5125 ;
      RECT  111.9575 0.14 122.9825 0.2775 ;
      RECT  31.85 12.1825 32.265 14.2375 ;
      RECT  31.85 14.6525 32.265 19.0375 ;
      RECT  25.5 32.9075 25.915 35.4825 ;
      RECT  25.5 35.8975 25.915 44.4525 ;
      RECT  174.8 43.3725 175.215 44.4525 ;
      RECT  174.8 44.8675 175.215 47.4425 ;
      RECT  24.875 38.8875 25.29 41.4625 ;
      RECT  24.875 41.8775 25.29 44.4525 ;
      RECT  174.175 26.9275 174.59 29.5025 ;
      RECT  174.175 29.9175 174.59 32.4925 ;
      RECT  171.4 229.2225 197.725 229.9125 ;
      RECT  171.4 229.9125 197.725 230.05 ;
      RECT  197.725 229.2225 198.14 229.9125 ;
      RECT  198.14 229.2225 199.865 229.9125 ;
      RECT  198.14 229.9125 199.865 230.05 ;
      RECT  0.14 0.2775 28.6025 0.9675 ;
      RECT  28.6025 0.2775 29.0175 0.9675 ;
      RECT  29.0175 0.2775 40.325 0.9675 ;
      RECT  40.2875 8.625 40.325 10.325 ;
      RECT  40.2875 10.675 40.325 14.045 ;
      RECT  40.325 8.625 40.74 10.325 ;
      RECT  40.325 10.675 40.74 14.045 ;
      RECT  40.74 8.625 43.4725 10.325 ;
      RECT  40.74 10.675 43.4725 14.045 ;
      RECT  43.4725 8.625 43.8875 10.325 ;
      RECT  43.4725 10.675 43.8875 14.045 ;
      RECT  43.8875 8.625 155.0075 10.325 ;
      RECT  43.8875 10.675 155.0075 14.045 ;
      RECT  40.74 227.89 168.4075 228.58 ;
      RECT  40.74 228.58 168.4075 228.995 ;
      RECT  40.74 228.995 168.4075 230.05 ;
      RECT  168.4075 227.89 168.8225 228.58 ;
      RECT  168.4075 228.995 168.8225 230.05 ;
      RECT  168.8225 227.89 170.985 228.58 ;
      RECT  168.8225 228.58 170.985 228.995 ;
      RECT  168.8225 228.995 170.985 230.05 ;
      RECT  29.0175 0.14 31.4625 0.2775 ;
      RECT  31.8775 0.14 40.325 0.2775 ;
      RECT  54.7575 0.14 65.7825 0.2775 ;
      RECT  66.1975 0.14 77.2225 0.2775 ;
      RECT  146.2775 0.14 157.3025 0.2775 ;
      RECT  157.7175 0.14 168.7425 0.2775 ;
      RECT  123.3975 0.14 134.4225 0.2775 ;
      RECT  134.8375 0.14 145.8625 0.2775 ;
      RECT  174.175 32.9075 174.59 35.4825 ;
      RECT  174.175 35.8975 174.59 42.9575 ;
      RECT  174.8 38.8875 175.215 41.4625 ;
      RECT  174.8 41.8775 175.215 42.9575 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  2.7 0.14 28.6025 0.2775 ;
      RECT  167.825 220.8925 168.24 222.9475 ;
      RECT  167.825 223.3625 168.24 225.0525 ;
      RECT  174.175 19.8425 174.59 20.5325 ;
      RECT  174.8 47.8575 175.215 50.4325 ;
      RECT  174.8 50.8475 175.215 227.475 ;
      RECT  25.5 26.9275 25.915 29.5025 ;
      RECT  25.5 29.9175 25.915 32.4925 ;
      RECT  40.74 0.14 42.9025 0.2775 ;
      RECT  43.3175 0.14 54.3425 0.2775 ;
      RECT  77.6375 0.14 88.6625 0.2775 ;
      RECT  89.0775 0.14 100.1025 0.2775 ;
      RECT  24.875 47.8575 25.29 50.4325 ;
      RECT  24.875 50.8475 25.29 51.5375 ;
      RECT  174.175 20.9475 174.59 23.5225 ;
      RECT  174.175 23.9375 174.59 26.5125 ;
   LAYER  metal4 ;
      RECT  0.14 212.52 33.0 230.05 ;
      RECT  33.0 212.52 33.7 230.05 ;
      RECT  33.7 0.14 179.705 3.035 ;
      RECT  179.705 0.14 180.405 3.035 ;
      RECT  180.405 0.14 200.285 3.035 ;
      RECT  180.405 3.035 200.285 20.39 ;
      RECT  179.705 21.09 180.405 212.52 ;
      RECT  180.405 20.39 200.285 21.09 ;
      RECT  0.14 50.29 19.88 68.345 ;
      RECT  0.14 68.345 19.88 212.52 ;
      RECT  19.88 20.39 20.58 50.29 ;
      RECT  19.88 68.345 20.58 212.52 ;
      RECT  39.0 212.45 39.7 212.52 ;
      RECT  33.7 217.42 176.985 228.0 ;
      RECT  33.7 228.0 176.985 230.05 ;
      RECT  176.985 212.52 177.685 217.42 ;
      RECT  176.985 228.0 177.685 230.05 ;
      RECT  33.7 3.035 40.08 17.22 ;
      RECT  40.08 3.035 40.78 17.22 ;
      RECT  39.7 20.39 40.08 21.09 ;
      RECT  39.7 21.09 40.08 212.45 ;
      RECT  39.7 212.45 40.08 212.52 ;
      RECT  33.7 212.52 40.08 215.37 ;
      RECT  33.7 215.37 40.08 217.42 ;
      RECT  40.08 215.37 40.78 217.42 ;
      RECT  40.78 215.37 176.985 217.42 ;
      RECT  0.14 0.14 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 20.39 ;
      RECT  0.4075 0.14 1.1075 9.5675 ;
      RECT  0.14 20.39 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 50.29 ;
      RECT  0.4075 32.53 1.1075 50.29 ;
      RECT  160.01 212.52 176.985 215.37 ;
      RECT  160.01 20.39 160.39 21.09 ;
      RECT  160.01 21.09 160.39 212.45 ;
      RECT  199.3175 21.09 200.0175 197.66 ;
      RECT  200.0175 21.09 200.285 197.66 ;
      RECT  200.0175 197.66 200.285 212.52 ;
      RECT  200.0175 212.52 200.285 217.42 ;
      RECT  199.3175 220.6225 200.0175 228.0 ;
      RECT  200.0175 217.42 200.285 220.6225 ;
      RECT  200.0175 220.6225 200.285 228.0 ;
      RECT  22.6 0.14 23.3 2.19 ;
      RECT  23.3 0.14 33.0 2.19 ;
      RECT  23.3 2.19 33.0 9.5675 ;
      RECT  22.6 17.71 23.3 20.39 ;
      RECT  23.3 9.5675 33.0 17.71 ;
      RECT  20.58 20.39 22.74 50.225 ;
      RECT  20.58 50.225 22.74 50.29 ;
      RECT  22.74 20.39 23.44 50.225 ;
      RECT  20.58 50.29 22.74 68.28 ;
      RECT  20.58 68.28 22.74 68.345 ;
      RECT  22.74 68.28 23.44 68.345 ;
      RECT  40.78 3.035 176.845 3.1 ;
      RECT  40.78 3.1 176.845 17.22 ;
      RECT  176.845 3.035 177.545 3.1 ;
      RECT  177.545 3.035 179.705 3.1 ;
      RECT  177.545 3.1 179.705 17.22 ;
      RECT  177.545 17.22 179.705 20.39 ;
      RECT  177.545 20.39 179.705 21.09 ;
      RECT  176.845 21.155 177.545 212.45 ;
      RECT  177.545 21.09 179.705 21.155 ;
      RECT  177.545 21.155 179.705 212.45 ;
      RECT  161.09 20.39 165.83 21.09 ;
      RECT  161.09 21.09 165.83 212.45 ;
      RECT  160.01 212.45 165.83 212.4825 ;
      RECT  160.01 212.4825 165.83 212.52 ;
      RECT  165.83 212.4825 166.39 212.52 ;
      RECT  160.01 17.22 165.83 20.3575 ;
      RECT  160.01 20.3575 165.83 20.39 ;
      RECT  165.83 17.22 166.53 20.3575 ;
      RECT  166.53 17.22 176.845 20.3575 ;
      RECT  177.685 228.0 193.76 230.05 ;
      RECT  194.46 228.0 200.285 230.05 ;
      RECT  177.685 212.52 193.76 214.95 ;
      RECT  177.685 214.95 193.76 217.42 ;
      RECT  193.76 212.52 194.46 214.95 ;
      RECT  177.685 217.42 193.76 220.6225 ;
      RECT  177.685 220.6225 193.76 228.0 ;
      RECT  194.46 220.6225 199.3175 228.0 ;
      RECT  20.58 68.345 31.065 212.52 ;
      RECT  31.765 68.345 33.0 212.52 ;
      RECT  23.3 17.71 31.065 20.3575 ;
      RECT  23.3 20.3575 31.065 20.39 ;
      RECT  31.065 17.71 31.765 20.3575 ;
      RECT  31.765 17.71 33.0 20.3575 ;
      RECT  31.765 20.3575 33.0 20.39 ;
      RECT  23.44 20.39 31.065 50.225 ;
      RECT  31.765 20.39 33.0 50.225 ;
      RECT  23.44 50.225 31.065 50.29 ;
      RECT  31.765 50.225 33.0 50.29 ;
      RECT  23.44 50.29 31.065 68.28 ;
      RECT  31.765 50.29 33.0 68.28 ;
      RECT  23.44 68.28 31.065 68.345 ;
      RECT  31.765 68.28 33.0 68.345 ;
      RECT  1.1075 0.14 5.825 2.19 ;
      RECT  6.525 0.14 22.6 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 22.6 9.5675 ;
      RECT  5.825 15.24 6.525 17.71 ;
      RECT  6.525 9.5675 22.6 15.24 ;
      RECT  6.525 15.24 22.6 17.71 ;
      RECT  1.1075 20.39 2.47 32.53 ;
      RECT  3.17 20.39 19.88 32.53 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 50.29 ;
      RECT  2.47 32.5625 3.17 50.29 ;
      RECT  3.17 32.53 19.88 32.5625 ;
      RECT  3.17 32.5625 19.88 50.29 ;
      RECT  1.1075 17.71 2.47 20.39 ;
      RECT  3.17 17.71 22.6 20.39 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 15.24 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  1.1075 15.24 2.47 17.71 ;
      RECT  3.17 15.24 5.825 17.71 ;
      RECT  180.405 21.09 197.255 197.6275 ;
      RECT  180.405 197.6275 197.255 197.66 ;
      RECT  197.255 21.09 197.955 197.6275 ;
      RECT  197.955 21.09 199.3175 197.6275 ;
      RECT  197.955 197.6275 199.3175 197.66 ;
      RECT  180.405 197.66 197.255 212.52 ;
      RECT  197.955 197.66 199.3175 212.52 ;
      RECT  194.46 212.52 197.255 214.95 ;
      RECT  197.955 212.52 199.3175 214.95 ;
      RECT  194.46 214.95 197.255 217.42 ;
      RECT  197.955 214.95 199.3175 217.42 ;
      RECT  194.46 217.42 197.255 220.59 ;
      RECT  194.46 220.59 197.255 220.6225 ;
      RECT  197.255 220.59 197.955 220.6225 ;
      RECT  197.955 217.42 199.3175 220.59 ;
      RECT  197.955 220.59 199.3175 220.6225 ;
      RECT  167.09 212.45 168.325 212.52 ;
      RECT  169.025 212.45 179.705 212.52 ;
      RECT  167.09 20.39 168.325 21.09 ;
      RECT  169.025 20.39 176.845 21.09 ;
      RECT  167.09 21.09 168.325 21.155 ;
      RECT  169.025 21.09 176.845 21.155 ;
      RECT  167.09 21.155 168.325 212.45 ;
      RECT  169.025 21.155 176.845 212.45 ;
      RECT  166.53 20.3575 168.325 20.39 ;
      RECT  169.025 20.3575 176.845 20.39 ;
      RECT  41.24 17.22 158.85 20.39 ;
      RECT  41.24 212.45 158.85 212.52 ;
      RECT  41.24 212.52 158.85 215.37 ;
      RECT  41.24 20.39 158.85 21.09 ;
      RECT  41.24 21.09 158.85 212.45 ;
      RECT  33.0 0.14 33.56 20.3575 ;
      RECT  33.0 20.3575 33.56 20.39 ;
      RECT  33.56 0.14 33.7 20.3575 ;
      RECT  34.26 20.39 39.0 21.09 ;
      RECT  34.26 21.09 39.0 212.45 ;
      RECT  33.7 212.4825 34.26 212.52 ;
      RECT  34.26 212.45 39.0 212.4825 ;
      RECT  34.26 212.4825 39.0 212.52 ;
      RECT  33.7 17.22 34.26 20.3575 ;
      RECT  34.26 17.22 40.08 20.3575 ;
      RECT  34.26 20.3575 40.08 20.39 ;
   END
END    freepdk45_sram_1w1r_256x48_12
END    LIBRARY
