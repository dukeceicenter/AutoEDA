../macros/freepdk45_sram_1rw0r_64x80_20/freepdk45_sram_1rw0r_64x80_20.lef