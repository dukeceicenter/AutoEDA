VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_14x128
   CLASS BLOCK ;
   SIZE 131.805 BY 88.705 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.91 1.105 24.045 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.77 1.105 26.905 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.63 1.105 29.765 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.49 1.105 32.625 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.35 1.105 35.485 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.21 1.105 38.345 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.07 1.105 41.205 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.93 1.105 44.065 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.79 1.105 46.925 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.65 1.105 49.785 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.51 1.105 52.645 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.37 1.105 55.505 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.23 1.105 58.365 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.09 1.105 61.225 1.24 ;
      END
   END din0[13]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  18.19 1.105 18.325 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.05 1.105 21.185 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.47 43.37 12.605 43.505 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.47 46.1 12.605 46.235 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.47 48.31 12.605 48.445 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.47 51.04 12.605 51.175 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.47 53.25 12.605 53.385 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.48 87.465 110.615 87.6 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.62 87.465 107.755 87.6 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.06 20.23 119.195 20.365 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.06 17.5 119.195 17.635 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.06 15.29 119.195 15.425 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.06 12.56 119.195 12.695 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.06 10.35 119.195 10.485 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.77 0.42 1.905 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.385 86.09 131.52 86.225 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.855 6.3825 1.99 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.2825 86.005 125.4175 86.14 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.8025 82.5975 32.9375 82.7325 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.5025 82.5975 37.6375 82.7325 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.2025 82.5975 42.3375 82.7325 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.9025 82.5975 47.0375 82.7325 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.6025 82.5975 51.7375 82.7325 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.3025 82.5975 56.4375 82.7325 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.0025 82.5975 61.1375 82.7325 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.7025 82.5975 65.8375 82.7325 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.4025 82.5975 70.5375 82.7325 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.1025 82.5975 75.2375 82.7325 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.8025 82.5975 79.9375 82.7325 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.5025 82.5975 84.6375 82.7325 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.2025 82.5975 89.3375 82.7325 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.9025 82.5975 94.0375 82.7325 ;
      END
   END dout1[13]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  109.055 75.32 109.195 85.34 ;
         LAYER metal4 ;
         RECT  28.47 21.3325 28.61 69.3125 ;
         LAYER metal3 ;
         RECT  112.7675 31.8 112.9025 31.935 ;
         LAYER metal3 ;
         RECT  112.4225 22.83 112.5575 22.965 ;
         LAYER metal3 ;
         RECT  112.7675 37.78 112.9025 37.915 ;
         LAYER metal4 ;
         RECT  130.9775 55.0825 131.1175 77.485 ;
         LAYER metal3 ;
         RECT  23.6275 2.47 23.7625 2.605 ;
         LAYER metal3 ;
         RECT  112.4225 25.82 112.5575 25.955 ;
         LAYER metal3 ;
         RECT  18.9125 25.82 19.0475 25.955 ;
         LAYER metal3 ;
         RECT  102.8625 70.67 102.9975 70.805 ;
         LAYER metal3 ;
         RECT  112.7675 34.79 112.9025 34.925 ;
         LAYER metal3 ;
         RECT  29.6175 17.4675 98.7025 17.5375 ;
         LAYER metal3 ;
         RECT  17.9075 2.47 18.0425 2.605 ;
         LAYER metal3 ;
         RECT  35.0675 2.47 35.2025 2.605 ;
         LAYER metal4 ;
         RECT  14.905 3.1325 15.045 18.0925 ;
         LAYER metal3 ;
         RECT  112.7675 40.77 112.9025 40.905 ;
         LAYER metal3 ;
         RECT  29.6175 8.8175 94.7075 8.8875 ;
         LAYER metal3 ;
         RECT  18.5675 34.79 18.7025 34.925 ;
         LAYER metal3 ;
         RECT  29.6175 80.04 94.7075 80.11 ;
         LAYER metal3 ;
         RECT  28.4725 19.84 28.6075 19.975 ;
         LAYER metal4 ;
         RECT  116.62 74.8425 116.76 84.8625 ;
         LAYER metal4 ;
         RECT  22.275 5.125 22.415 15.145 ;
         LAYER metal4 ;
         RECT  29.55 18.1625 29.69 72.2325 ;
         LAYER metal3 ;
         RECT  18.9125 22.83 19.0475 22.965 ;
         LAYER metal4 ;
         RECT  12.185 42.2625 12.325 54.8175 ;
         LAYER metal3 ;
         RECT  106.595 69.8825 106.73 70.0175 ;
         LAYER metal3 ;
         RECT  2.425 3.135 2.56 3.27 ;
         LAYER metal4 ;
         RECT  102.86 21.3325 103.0 69.3125 ;
         LAYER metal4 ;
         RECT  24.12 21.3325 24.26 69.3825 ;
         LAYER metal3 ;
         RECT  57.9475 2.47 58.0825 2.605 ;
         LAYER metal3 ;
         RECT  18.5675 37.78 18.7025 37.915 ;
         LAYER metal4 ;
         RECT  0.6875 10.51 0.8275 32.9125 ;
         LAYER metal4 ;
         RECT  101.78 18.1625 101.92 72.2325 ;
         LAYER metal3 ;
         RECT  29.6175 72.9275 99.8775 72.9975 ;
         LAYER metal3 ;
         RECT  18.5675 31.8 18.7025 31.935 ;
         LAYER metal3 ;
         RECT  129.245 84.725 129.38 84.86 ;
         LAYER metal4 ;
         RECT  107.21 21.3325 107.35 69.3825 ;
         LAYER metal4 ;
         RECT  119.34 8.9175 119.48 21.4725 ;
         LAYER metal3 ;
         RECT  46.5075 2.47 46.6425 2.605 ;
         LAYER metal3 ;
         RECT  18.5675 40.77 18.7025 40.905 ;
         LAYER metal3 ;
         RECT  24.74 20.6275 24.875 20.7625 ;
         LAYER metal3 ;
         RECT  110.7625 86.1 110.8975 86.235 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  49.3675 0.0 49.5025 0.135 ;
         LAYER metal3 ;
         RECT  114.575 30.305 114.71 30.44 ;
         LAYER metal4 ;
         RECT  20.6125 5.0575 20.7525 15.2125 ;
         LAYER metal3 ;
         RECT  113.95 27.315 114.085 27.45 ;
         LAYER metal4 ;
         RECT  125.42 72.3725 125.56 87.3325 ;
         LAYER metal4 ;
         RECT  22.53 21.3 22.67 69.3825 ;
         LAYER metal4 ;
         RECT  106.65 21.3 106.79 69.345 ;
         LAYER metal3 ;
         RECT  113.95 24.325 114.085 24.46 ;
         LAYER metal4 ;
         RECT  128.915 55.05 129.055 77.4525 ;
         LAYER metal3 ;
         RECT  16.76 39.275 16.895 39.41 ;
         LAYER metal3 ;
         RECT  17.385 21.335 17.52 21.47 ;
         LAYER metal3 ;
         RECT  16.76 30.305 16.895 30.44 ;
         LAYER metal3 ;
         RECT  29.6175 14.8475 98.735 14.9175 ;
         LAYER metal3 ;
         RECT  114.575 33.295 114.71 33.43 ;
         LAYER metal3 ;
         RECT  29.6175 75.5475 98.735 75.6175 ;
         LAYER metal4 ;
         RECT  110.7175 75.2525 110.8575 85.4075 ;
         LAYER metal3 ;
         RECT  17.385 24.325 17.52 24.46 ;
         LAYER metal3 ;
         RECT  26.4875 0.0 26.6225 0.135 ;
         LAYER metal3 ;
         RECT  107.9025 88.57 108.0375 88.705 ;
         LAYER metal3 ;
         RECT  29.6175 78.1475 94.7425 78.2175 ;
         LAYER metal4 ;
         RECT  15.045 42.1975 15.185 54.7525 ;
         LAYER metal4 ;
         RECT  2.75 10.5425 2.89 32.945 ;
         LAYER metal3 ;
         RECT  20.7675 0.0 20.9025 0.135 ;
         LAYER metal3 ;
         RECT  16.76 42.265 16.895 42.4 ;
         LAYER metal3 ;
         RECT  16.76 36.285 16.895 36.42 ;
         LAYER metal3 ;
         RECT  60.8075 0.0 60.9425 0.135 ;
         LAYER metal3 ;
         RECT  114.575 36.285 114.71 36.42 ;
         LAYER metal3 ;
         RECT  129.245 87.195 129.38 87.33 ;
         LAYER metal3 ;
         RECT  16.76 33.295 16.895 33.43 ;
         LAYER metal4 ;
         RECT  6.105 0.6625 6.245 15.6225 ;
         LAYER metal4 ;
         RECT  108.8 21.3 108.94 69.3825 ;
         LAYER metal3 ;
         RECT  17.385 27.315 17.52 27.45 ;
         LAYER metal3 ;
         RECT  29.6175 10.8675 94.7075 10.9375 ;
         LAYER metal4 ;
         RECT  24.68 21.3 24.82 69.345 ;
         LAYER metal3 ;
         RECT  114.575 39.275 114.71 39.41 ;
         LAYER metal4 ;
         RECT  30.01 18.1625 30.15 72.2325 ;
         LAYER metal4 ;
         RECT  101.32 18.1625 101.46 72.2325 ;
         LAYER metal4 ;
         RECT  116.48 8.9825 116.62 21.5375 ;
         LAYER metal3 ;
         RECT  113.95 21.335 114.085 21.47 ;
         LAYER metal3 ;
         RECT  2.425 0.665 2.56 0.8 ;
         LAYER metal3 ;
         RECT  114.575 42.265 114.71 42.4 ;
         LAYER metal3 ;
         RECT  37.9275 0.0 38.0625 0.135 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 131.665 88.565 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 131.665 88.565 ;
   LAYER  metal3 ;
      RECT  23.77 0.14 24.185 0.965 ;
      RECT  24.185 0.965 26.63 1.38 ;
      RECT  27.045 0.965 29.49 1.38 ;
      RECT  29.905 0.965 32.35 1.38 ;
      RECT  32.765 0.965 35.21 1.38 ;
      RECT  35.625 0.965 38.07 1.38 ;
      RECT  38.485 0.965 40.93 1.38 ;
      RECT  41.345 0.965 43.79 1.38 ;
      RECT  44.205 0.965 46.65 1.38 ;
      RECT  47.065 0.965 49.51 1.38 ;
      RECT  49.925 0.965 52.37 1.38 ;
      RECT  52.785 0.965 55.23 1.38 ;
      RECT  55.645 0.965 58.09 1.38 ;
      RECT  58.505 0.965 60.95 1.38 ;
      RECT  61.365 0.965 131.665 1.38 ;
      RECT  0.14 0.965 18.05 1.38 ;
      RECT  18.465 0.965 20.91 1.38 ;
      RECT  21.325 0.965 23.77 1.38 ;
      RECT  0.14 43.23 12.33 43.645 ;
      RECT  0.14 43.645 12.33 88.565 ;
      RECT  12.33 1.38 12.745 43.23 ;
      RECT  12.745 43.23 23.77 43.645 ;
      RECT  12.745 43.645 23.77 88.565 ;
      RECT  12.33 43.645 12.745 45.96 ;
      RECT  12.33 46.375 12.745 48.17 ;
      RECT  12.33 48.585 12.745 50.9 ;
      RECT  12.33 51.315 12.745 53.11 ;
      RECT  12.33 53.525 12.745 88.565 ;
      RECT  110.34 87.74 110.755 88.565 ;
      RECT  110.755 87.74 131.665 88.565 ;
      RECT  24.185 87.325 107.48 87.74 ;
      RECT  107.895 87.325 110.34 87.74 ;
      RECT  110.755 1.38 118.92 20.09 ;
      RECT  110.755 20.09 118.92 20.505 ;
      RECT  118.92 20.505 119.335 87.325 ;
      RECT  119.335 1.38 131.665 20.09 ;
      RECT  119.335 20.09 131.665 20.505 ;
      RECT  118.92 17.775 119.335 20.09 ;
      RECT  118.92 15.565 119.335 17.36 ;
      RECT  118.92 12.835 119.335 15.15 ;
      RECT  118.92 1.38 119.335 10.21 ;
      RECT  118.92 10.625 119.335 12.42 ;
      RECT  0.14 1.38 0.145 1.63 ;
      RECT  0.14 1.63 0.145 2.045 ;
      RECT  0.14 2.045 0.145 43.23 ;
      RECT  0.145 1.38 0.56 1.63 ;
      RECT  0.145 2.045 0.56 43.23 ;
      RECT  0.56 1.38 12.33 1.63 ;
      RECT  131.245 20.505 131.66 85.95 ;
      RECT  131.245 86.365 131.66 87.325 ;
      RECT  131.66 20.505 131.665 85.95 ;
      RECT  131.66 85.95 131.665 86.365 ;
      RECT  131.66 86.365 131.665 87.325 ;
      RECT  0.56 1.63 6.1075 1.715 ;
      RECT  0.56 1.715 6.1075 2.045 ;
      RECT  6.1075 1.63 6.5225 1.715 ;
      RECT  6.5225 1.63 12.33 1.715 ;
      RECT  6.5225 1.715 12.33 2.045 ;
      RECT  0.56 2.045 6.1075 2.13 ;
      RECT  6.1075 2.13 6.5225 43.23 ;
      RECT  6.5225 2.045 12.33 2.13 ;
      RECT  6.5225 2.13 12.33 43.23 ;
      RECT  119.335 20.505 125.1425 85.865 ;
      RECT  119.335 85.865 125.1425 85.95 ;
      RECT  125.1425 20.505 125.5575 85.865 ;
      RECT  125.5575 85.865 131.245 85.95 ;
      RECT  119.335 85.95 125.1425 86.28 ;
      RECT  119.335 86.28 125.1425 86.365 ;
      RECT  125.1425 86.28 125.5575 86.365 ;
      RECT  125.5575 85.95 131.245 86.28 ;
      RECT  125.5575 86.28 131.245 86.365 ;
      RECT  24.185 82.4575 32.6625 82.8725 ;
      RECT  24.185 82.8725 32.6625 87.325 ;
      RECT  32.6625 82.8725 33.0775 87.325 ;
      RECT  33.0775 82.8725 110.34 87.325 ;
      RECT  33.0775 82.4575 37.3625 82.8725 ;
      RECT  37.7775 82.4575 42.0625 82.8725 ;
      RECT  42.4775 82.4575 46.7625 82.8725 ;
      RECT  47.1775 82.4575 51.4625 82.8725 ;
      RECT  51.8775 82.4575 56.1625 82.8725 ;
      RECT  56.5775 82.4575 60.8625 82.8725 ;
      RECT  61.2775 82.4575 65.5625 82.8725 ;
      RECT  65.9775 82.4575 70.2625 82.8725 ;
      RECT  70.6775 82.4575 74.9625 82.8725 ;
      RECT  75.3775 82.4575 79.6625 82.8725 ;
      RECT  80.0775 82.4575 84.3625 82.8725 ;
      RECT  84.7775 82.4575 89.0625 82.8725 ;
      RECT  89.4775 82.4575 93.7625 82.8725 ;
      RECT  94.1775 82.4575 110.34 82.8725 ;
      RECT  110.755 31.66 112.6275 32.075 ;
      RECT  113.0425 31.66 118.92 32.075 ;
      RECT  110.755 20.505 112.2825 22.69 ;
      RECT  110.755 22.69 112.2825 23.105 ;
      RECT  110.755 23.105 112.2825 31.66 ;
      RECT  112.2825 20.505 112.6275 22.69 ;
      RECT  112.6275 20.505 112.6975 22.69 ;
      RECT  112.6975 20.505 113.0425 22.69 ;
      RECT  112.6975 22.69 113.0425 23.105 ;
      RECT  112.6975 23.105 113.0425 31.66 ;
      RECT  23.77 1.38 23.9025 2.33 ;
      RECT  23.77 2.745 23.9025 88.565 ;
      RECT  23.9025 1.38 24.185 2.33 ;
      RECT  23.9025 2.33 24.185 2.745 ;
      RECT  23.9025 2.745 24.185 88.565 ;
      RECT  12.745 1.38 23.4875 2.33 ;
      RECT  23.4875 1.38 23.77 2.33 ;
      RECT  23.4875 2.745 23.77 43.23 ;
      RECT  112.2825 23.105 112.6275 25.68 ;
      RECT  112.2825 26.095 112.6275 31.66 ;
      RECT  112.6275 23.105 112.6975 25.68 ;
      RECT  112.6275 26.095 112.6975 31.66 ;
      RECT  12.745 25.68 18.7725 26.095 ;
      RECT  19.1875 2.745 23.4875 25.68 ;
      RECT  19.1875 25.68 23.4875 26.095 ;
      RECT  19.1875 26.095 23.4875 43.23 ;
      RECT  33.0775 70.53 102.7225 70.945 ;
      RECT  102.7225 1.38 103.1375 70.53 ;
      RECT  102.7225 70.945 103.1375 82.4575 ;
      RECT  103.1375 70.53 110.34 70.945 ;
      RECT  103.1375 70.945 110.34 82.4575 ;
      RECT  112.6275 32.075 113.0425 34.65 ;
      RECT  112.6275 35.065 113.0425 37.64 ;
      RECT  24.185 1.38 29.4775 17.3275 ;
      RECT  24.185 17.3275 29.4775 17.6775 ;
      RECT  33.0775 17.6775 98.8425 70.53 ;
      RECT  98.8425 17.3275 102.7225 17.6775 ;
      RECT  98.8425 17.6775 102.7225 70.53 ;
      RECT  12.745 2.33 17.7675 2.745 ;
      RECT  18.1825 2.33 23.4875 2.745 ;
      RECT  33.0775 1.38 34.9275 2.33 ;
      RECT  33.0775 2.33 34.9275 2.745 ;
      RECT  34.9275 1.38 35.3425 2.33 ;
      RECT  35.3425 1.38 98.8425 2.33 ;
      RECT  112.6275 38.055 113.0425 40.63 ;
      RECT  112.6275 41.045 113.0425 87.325 ;
      RECT  29.4775 1.38 32.6625 8.6775 ;
      RECT  32.6625 1.38 33.0775 8.6775 ;
      RECT  33.0775 2.745 34.9275 8.6775 ;
      RECT  34.9275 2.745 35.3425 8.6775 ;
      RECT  35.3425 2.745 94.8475 8.6775 ;
      RECT  94.8475 2.745 98.8425 8.6775 ;
      RECT  94.8475 8.6775 98.8425 9.0275 ;
      RECT  12.745 34.65 18.4275 35.065 ;
      RECT  18.8425 26.095 19.1875 34.65 ;
      RECT  18.8425 34.65 19.1875 35.065 ;
      RECT  18.8425 35.065 19.1875 43.23 ;
      RECT  33.0775 80.25 94.8475 82.4575 ;
      RECT  94.8475 79.9 102.7225 80.25 ;
      RECT  94.8475 80.25 102.7225 82.4575 ;
      RECT  29.4775 80.25 32.6625 82.4575 ;
      RECT  32.6625 80.25 33.0775 82.4575 ;
      RECT  24.185 17.6775 28.3325 19.7 ;
      RECT  24.185 19.7 28.3325 20.115 ;
      RECT  28.3325 17.6775 28.7475 19.7 ;
      RECT  28.3325 20.115 28.7475 82.4575 ;
      RECT  28.7475 17.6775 29.4775 19.7 ;
      RECT  28.7475 19.7 29.4775 20.115 ;
      RECT  28.7475 20.115 29.4775 82.4575 ;
      RECT  18.7725 2.745 19.1875 22.69 ;
      RECT  18.7725 23.105 19.1875 25.68 ;
      RECT  103.1375 1.38 106.455 69.7425 ;
      RECT  103.1375 69.7425 106.455 70.1575 ;
      RECT  103.1375 70.1575 106.455 70.53 ;
      RECT  106.455 1.38 106.87 69.7425 ;
      RECT  106.455 70.1575 106.87 70.53 ;
      RECT  106.87 1.38 110.34 69.7425 ;
      RECT  106.87 69.7425 110.34 70.1575 ;
      RECT  106.87 70.1575 110.34 70.53 ;
      RECT  0.56 2.13 2.285 2.995 ;
      RECT  0.56 2.995 2.285 3.41 ;
      RECT  0.56 3.41 2.285 43.23 ;
      RECT  2.285 2.13 2.7 2.995 ;
      RECT  2.285 3.41 2.7 43.23 ;
      RECT  2.7 2.13 6.1075 2.995 ;
      RECT  2.7 2.995 6.1075 3.41 ;
      RECT  2.7 3.41 6.1075 43.23 ;
      RECT  58.2225 2.33 98.8425 2.745 ;
      RECT  18.4275 35.065 18.7725 37.64 ;
      RECT  18.7725 35.065 18.8425 37.64 ;
      RECT  33.0775 70.945 94.8475 72.7875 ;
      RECT  94.8475 70.945 100.0175 72.7875 ;
      RECT  100.0175 70.945 102.7225 72.7875 ;
      RECT  100.0175 72.7875 102.7225 73.1375 ;
      RECT  100.0175 73.1375 102.7225 79.9 ;
      RECT  29.4775 17.6775 32.6625 72.7875 ;
      RECT  32.6625 17.6775 33.0775 72.7875 ;
      RECT  18.4275 26.095 18.7725 31.66 ;
      RECT  18.4275 32.075 18.7725 34.65 ;
      RECT  18.7725 26.095 18.8425 31.66 ;
      RECT  18.7725 32.075 18.8425 34.65 ;
      RECT  125.5575 20.505 129.105 84.585 ;
      RECT  125.5575 84.585 129.105 85.0 ;
      RECT  125.5575 85.0 129.105 85.865 ;
      RECT  129.105 20.505 129.52 84.585 ;
      RECT  129.105 85.0 129.52 85.865 ;
      RECT  129.52 20.505 131.245 84.585 ;
      RECT  129.52 84.585 131.245 85.0 ;
      RECT  129.52 85.0 131.245 85.865 ;
      RECT  35.3425 2.33 46.3675 2.745 ;
      RECT  46.7825 2.33 57.8075 2.745 ;
      RECT  18.4275 38.055 18.7725 40.63 ;
      RECT  18.4275 41.045 18.7725 43.23 ;
      RECT  18.7725 38.055 18.8425 40.63 ;
      RECT  18.7725 41.045 18.8425 43.23 ;
      RECT  24.185 20.115 24.6 20.4875 ;
      RECT  24.185 20.4875 24.6 20.9025 ;
      RECT  24.185 20.9025 24.6 82.4575 ;
      RECT  24.6 20.115 25.015 20.4875 ;
      RECT  24.6 20.9025 25.015 82.4575 ;
      RECT  25.015 20.115 28.3325 20.4875 ;
      RECT  25.015 20.4875 28.3325 20.9025 ;
      RECT  25.015 20.9025 28.3325 82.4575 ;
      RECT  110.34 1.38 110.6225 85.96 ;
      RECT  110.34 85.96 110.6225 86.375 ;
      RECT  110.34 86.375 110.6225 87.325 ;
      RECT  110.6225 1.38 110.755 85.96 ;
      RECT  110.6225 86.375 110.755 87.325 ;
      RECT  110.755 32.075 111.0375 85.96 ;
      RECT  110.755 86.375 111.0375 87.325 ;
      RECT  111.0375 32.075 112.6275 85.96 ;
      RECT  111.0375 85.96 112.6275 86.375 ;
      RECT  111.0375 86.375 112.6275 87.325 ;
      RECT  24.185 0.275 49.2275 0.965 ;
      RECT  49.2275 0.275 49.6425 0.965 ;
      RECT  49.6425 0.275 131.665 0.965 ;
      RECT  113.0425 30.165 114.435 30.58 ;
      RECT  113.0425 30.58 114.435 31.66 ;
      RECT  114.435 20.505 114.85 30.165 ;
      RECT  114.435 30.58 114.85 31.66 ;
      RECT  114.85 20.505 118.92 30.165 ;
      RECT  114.85 30.165 118.92 30.58 ;
      RECT  114.85 30.58 118.92 31.66 ;
      RECT  113.0425 20.505 113.81 27.175 ;
      RECT  113.0425 27.175 113.81 27.59 ;
      RECT  113.0425 27.59 113.81 30.165 ;
      RECT  113.81 27.59 114.225 30.165 ;
      RECT  114.225 20.505 114.435 27.175 ;
      RECT  114.225 27.175 114.435 27.59 ;
      RECT  114.225 27.59 114.435 30.165 ;
      RECT  113.81 24.6 114.225 27.175 ;
      RECT  12.745 35.065 16.62 39.135 ;
      RECT  12.745 39.135 16.62 39.55 ;
      RECT  12.745 39.55 16.62 43.23 ;
      RECT  17.035 35.065 18.4275 39.135 ;
      RECT  17.035 39.135 18.4275 39.55 ;
      RECT  17.035 39.55 18.4275 43.23 ;
      RECT  12.745 2.745 17.245 21.195 ;
      RECT  12.745 21.195 17.245 21.61 ;
      RECT  12.745 21.61 17.245 25.68 ;
      RECT  17.245 2.745 17.66 21.195 ;
      RECT  17.66 2.745 18.7725 21.195 ;
      RECT  17.66 21.195 18.7725 21.61 ;
      RECT  17.66 21.61 18.7725 25.68 ;
      RECT  12.745 26.095 16.62 30.165 ;
      RECT  12.745 30.165 16.62 30.58 ;
      RECT  12.745 30.58 16.62 34.65 ;
      RECT  16.62 26.095 17.035 30.165 ;
      RECT  17.035 30.165 18.4275 30.58 ;
      RECT  17.035 30.58 18.4275 34.65 ;
      RECT  98.8425 1.38 98.875 14.7075 ;
      RECT  98.8425 15.0575 98.875 17.3275 ;
      RECT  98.875 1.38 102.7225 14.7075 ;
      RECT  98.875 14.7075 102.7225 15.0575 ;
      RECT  98.875 15.0575 102.7225 17.3275 ;
      RECT  29.4775 15.0575 32.6625 17.3275 ;
      RECT  32.6625 15.0575 33.0775 17.3275 ;
      RECT  33.0775 15.0575 34.9275 17.3275 ;
      RECT  34.9275 15.0575 35.3425 17.3275 ;
      RECT  35.3425 15.0575 94.8475 17.3275 ;
      RECT  94.8475 9.0275 98.8425 14.7075 ;
      RECT  94.8475 15.0575 98.8425 17.3275 ;
      RECT  113.0425 32.075 114.435 33.155 ;
      RECT  113.0425 33.155 114.435 33.57 ;
      RECT  113.0425 33.57 114.435 87.325 ;
      RECT  114.435 32.075 114.85 33.155 ;
      RECT  114.85 32.075 118.92 33.155 ;
      RECT  114.85 33.155 118.92 33.57 ;
      RECT  114.85 33.57 118.92 87.325 ;
      RECT  33.0775 73.1375 94.8475 75.4075 ;
      RECT  94.8475 73.1375 98.875 75.4075 ;
      RECT  98.875 73.1375 100.0175 75.4075 ;
      RECT  98.875 75.4075 100.0175 75.7575 ;
      RECT  98.875 75.7575 100.0175 79.9 ;
      RECT  29.4775 73.1375 32.6625 75.4075 ;
      RECT  32.6625 73.1375 33.0775 75.4075 ;
      RECT  17.245 21.61 17.66 24.185 ;
      RECT  17.245 24.6 17.66 25.68 ;
      RECT  24.185 0.14 26.3475 0.275 ;
      RECT  24.185 87.74 107.7625 88.43 ;
      RECT  24.185 88.43 107.7625 88.565 ;
      RECT  107.7625 87.74 108.1775 88.43 ;
      RECT  108.1775 87.74 110.34 88.43 ;
      RECT  108.1775 88.43 110.34 88.565 ;
      RECT  33.0775 75.7575 94.8475 78.0075 ;
      RECT  33.0775 78.3575 94.8475 79.9 ;
      RECT  94.8475 75.7575 94.8825 78.0075 ;
      RECT  94.8475 78.3575 94.8825 79.9 ;
      RECT  94.8825 75.7575 98.875 78.0075 ;
      RECT  94.8825 78.0075 98.875 78.3575 ;
      RECT  94.8825 78.3575 98.875 79.9 ;
      RECT  29.4775 75.7575 32.6625 78.0075 ;
      RECT  29.4775 78.3575 32.6625 79.9 ;
      RECT  32.6625 75.7575 33.0775 78.0075 ;
      RECT  32.6625 78.3575 33.0775 79.9 ;
      RECT  0.14 0.14 20.6275 0.275 ;
      RECT  20.6275 0.275 21.0425 0.965 ;
      RECT  21.0425 0.14 23.77 0.275 ;
      RECT  21.0425 0.275 23.77 0.965 ;
      RECT  16.62 39.55 17.035 42.125 ;
      RECT  16.62 42.54 17.035 43.23 ;
      RECT  16.62 35.065 17.035 36.145 ;
      RECT  16.62 36.56 17.035 39.135 ;
      RECT  49.6425 0.14 60.6675 0.275 ;
      RECT  61.0825 0.14 131.665 0.275 ;
      RECT  114.435 33.57 114.85 36.145 ;
      RECT  110.755 87.325 129.105 87.47 ;
      RECT  110.755 87.47 129.105 87.74 ;
      RECT  129.105 87.47 129.52 87.74 ;
      RECT  129.52 87.325 131.665 87.47 ;
      RECT  129.52 87.47 131.665 87.74 ;
      RECT  119.335 86.365 129.105 87.055 ;
      RECT  119.335 87.055 129.105 87.325 ;
      RECT  129.105 86.365 129.52 87.055 ;
      RECT  129.52 86.365 131.245 87.055 ;
      RECT  129.52 87.055 131.245 87.325 ;
      RECT  16.62 30.58 17.035 33.155 ;
      RECT  16.62 33.57 17.035 34.65 ;
      RECT  17.035 26.095 17.245 27.175 ;
      RECT  17.035 27.175 17.245 27.59 ;
      RECT  17.035 27.59 17.245 30.165 ;
      RECT  17.245 26.095 17.66 27.175 ;
      RECT  17.245 27.59 17.66 30.165 ;
      RECT  17.66 26.095 18.4275 27.175 ;
      RECT  17.66 27.175 18.4275 27.59 ;
      RECT  17.66 27.59 18.4275 30.165 ;
      RECT  29.4775 9.0275 32.6625 10.7275 ;
      RECT  29.4775 11.0775 32.6625 14.7075 ;
      RECT  32.6625 9.0275 33.0775 10.7275 ;
      RECT  32.6625 11.0775 33.0775 14.7075 ;
      RECT  33.0775 9.0275 34.9275 10.7275 ;
      RECT  33.0775 11.0775 34.9275 14.7075 ;
      RECT  34.9275 9.0275 35.3425 10.7275 ;
      RECT  34.9275 11.0775 35.3425 14.7075 ;
      RECT  35.3425 9.0275 94.8475 10.7275 ;
      RECT  35.3425 11.0775 94.8475 14.7075 ;
      RECT  114.435 36.56 114.85 39.135 ;
      RECT  113.81 20.505 114.225 21.195 ;
      RECT  113.81 21.61 114.225 24.185 ;
      RECT  0.14 0.275 2.285 0.525 ;
      RECT  0.14 0.525 2.285 0.94 ;
      RECT  0.14 0.94 2.285 0.965 ;
      RECT  2.285 0.275 2.7 0.525 ;
      RECT  2.285 0.94 2.7 0.965 ;
      RECT  2.7 0.275 20.6275 0.525 ;
      RECT  2.7 0.525 20.6275 0.94 ;
      RECT  2.7 0.94 20.6275 0.965 ;
      RECT  114.435 39.55 114.85 42.125 ;
      RECT  114.435 42.54 114.85 87.325 ;
      RECT  26.7625 0.14 37.7875 0.275 ;
      RECT  38.2025 0.14 49.2275 0.275 ;
   LAYER  metal4 ;
      RECT  0.14 75.04 108.775 85.62 ;
      RECT  0.14 85.62 108.775 88.565 ;
      RECT  108.775 85.62 109.475 88.565 ;
      RECT  28.19 0.14 28.89 21.0525 ;
      RECT  28.19 69.5925 28.89 75.04 ;
      RECT  130.6975 0.14 131.3975 54.8025 ;
      RECT  131.3975 0.14 131.665 54.8025 ;
      RECT  131.3975 54.8025 131.665 75.04 ;
      RECT  130.6975 77.765 131.3975 85.62 ;
      RECT  131.3975 75.04 131.665 77.765 ;
      RECT  131.3975 77.765 131.665 85.62 ;
      RECT  14.625 0.14 15.325 2.8525 ;
      RECT  14.625 18.3725 15.325 21.0525 ;
      RECT  15.325 0.14 28.19 2.8525 ;
      RECT  109.475 54.8025 116.34 74.5625 ;
      RECT  116.34 54.8025 117.04 74.5625 ;
      RECT  116.34 85.1425 117.04 85.62 ;
      RECT  21.995 2.8525 22.695 4.845 ;
      RECT  21.995 15.425 22.695 18.3725 ;
      RECT  22.695 2.8525 28.19 4.845 ;
      RECT  22.695 4.845 28.19 15.425 ;
      RECT  22.695 15.425 28.19 18.3725 ;
      RECT  28.89 0.14 29.27 17.8825 ;
      RECT  28.89 17.8825 29.27 21.0525 ;
      RECT  29.27 0.14 29.97 17.8825 ;
      RECT  29.97 0.14 108.775 17.8825 ;
      RECT  28.89 21.0525 29.27 69.5925 ;
      RECT  28.89 69.5925 29.27 72.5125 ;
      RECT  28.89 72.5125 29.27 75.04 ;
      RECT  29.27 72.5125 29.97 75.04 ;
      RECT  29.97 72.5125 108.775 75.04 ;
      RECT  0.14 41.9825 11.905 55.0975 ;
      RECT  0.14 55.0975 11.905 69.5925 ;
      RECT  11.905 21.0525 12.605 41.9825 ;
      RECT  11.905 55.0975 12.605 69.5925 ;
      RECT  0.14 69.6625 23.84 75.04 ;
      RECT  23.84 69.6625 24.54 75.04 ;
      RECT  24.54 69.6625 28.19 75.04 ;
      RECT  0.14 2.8525 0.4075 10.23 ;
      RECT  0.14 10.23 0.4075 18.3725 ;
      RECT  0.4075 2.8525 1.1075 10.23 ;
      RECT  0.14 18.3725 0.4075 21.0525 ;
      RECT  0.14 21.0525 0.4075 33.1925 ;
      RECT  0.14 33.1925 0.4075 41.9825 ;
      RECT  0.4075 33.1925 1.1075 41.9825 ;
      RECT  102.2 21.0525 102.58 69.5925 ;
      RECT  102.2 69.6625 106.93 72.5125 ;
      RECT  106.93 69.6625 107.63 72.5125 ;
      RECT  107.63 69.6625 108.775 72.5125 ;
      RECT  109.475 0.14 119.06 8.6375 ;
      RECT  119.06 0.14 119.76 8.6375 ;
      RECT  119.06 21.7525 119.76 54.8025 ;
      RECT  119.76 0.14 130.6975 8.6375 ;
      RECT  119.76 8.6375 130.6975 21.7525 ;
      RECT  15.325 2.8525 20.3325 4.7775 ;
      RECT  15.325 4.7775 20.3325 4.845 ;
      RECT  20.3325 2.8525 21.0325 4.7775 ;
      RECT  21.0325 2.8525 21.995 4.7775 ;
      RECT  21.0325 4.7775 21.995 4.845 ;
      RECT  15.325 4.845 20.3325 15.425 ;
      RECT  21.0325 4.845 21.995 15.425 ;
      RECT  15.325 15.425 20.3325 15.4925 ;
      RECT  15.325 15.4925 20.3325 18.3725 ;
      RECT  20.3325 15.4925 21.0325 18.3725 ;
      RECT  21.0325 15.425 21.995 15.4925 ;
      RECT  21.0325 15.4925 21.995 18.3725 ;
      RECT  109.475 87.6125 125.14 88.565 ;
      RECT  125.14 87.6125 125.84 88.565 ;
      RECT  125.84 85.62 131.665 87.6125 ;
      RECT  125.84 87.6125 131.665 88.565 ;
      RECT  117.04 54.8025 125.14 72.0925 ;
      RECT  117.04 72.0925 125.14 74.5625 ;
      RECT  125.14 54.8025 125.84 72.0925 ;
      RECT  117.04 74.5625 125.14 75.04 ;
      RECT  117.04 75.04 125.14 77.765 ;
      RECT  117.04 77.765 125.14 85.1425 ;
      RECT  125.84 77.765 130.6975 85.1425 ;
      RECT  117.04 85.1425 125.14 85.62 ;
      RECT  125.84 85.1425 130.6975 85.62 ;
      RECT  15.325 18.3725 22.25 21.02 ;
      RECT  15.325 21.02 22.25 21.0525 ;
      RECT  22.25 18.3725 22.95 21.02 ;
      RECT  22.95 18.3725 28.19 21.02 ;
      RECT  0.14 69.5925 22.25 69.6625 ;
      RECT  22.95 69.5925 23.84 69.6625 ;
      RECT  22.95 21.0525 23.84 41.9825 ;
      RECT  22.95 41.9825 23.84 55.0975 ;
      RECT  12.605 55.0975 22.25 69.5925 ;
      RECT  22.95 55.0975 23.84 69.5925 ;
      RECT  102.2 17.8825 106.37 21.02 ;
      RECT  102.2 21.02 106.37 21.0525 ;
      RECT  106.37 17.8825 107.07 21.02 ;
      RECT  107.07 17.8825 108.775 21.02 ;
      RECT  103.28 21.0525 106.37 69.5925 ;
      RECT  102.2 69.5925 106.37 69.625 ;
      RECT  102.2 69.625 106.37 69.6625 ;
      RECT  106.37 69.625 106.93 69.6625 ;
      RECT  119.76 21.7525 128.635 54.77 ;
      RECT  119.76 54.77 128.635 54.8025 ;
      RECT  128.635 21.7525 129.335 54.77 ;
      RECT  129.335 21.7525 130.6975 54.77 ;
      RECT  129.335 54.77 130.6975 54.8025 ;
      RECT  125.84 54.8025 128.635 72.0925 ;
      RECT  129.335 54.8025 130.6975 72.0925 ;
      RECT  125.84 72.0925 128.635 74.5625 ;
      RECT  129.335 72.0925 130.6975 74.5625 ;
      RECT  125.84 74.5625 128.635 75.04 ;
      RECT  129.335 74.5625 130.6975 75.04 ;
      RECT  125.84 75.04 128.635 77.7325 ;
      RECT  125.84 77.7325 128.635 77.765 ;
      RECT  128.635 77.7325 129.335 77.765 ;
      RECT  129.335 75.04 130.6975 77.7325 ;
      RECT  129.335 77.7325 130.6975 77.765 ;
      RECT  109.475 74.5625 110.4375 74.9725 ;
      RECT  109.475 74.9725 110.4375 75.04 ;
      RECT  110.4375 74.5625 111.1375 74.9725 ;
      RECT  111.1375 74.5625 116.34 74.9725 ;
      RECT  111.1375 74.9725 116.34 75.04 ;
      RECT  109.475 75.04 110.4375 77.765 ;
      RECT  111.1375 75.04 116.34 77.765 ;
      RECT  109.475 77.765 110.4375 85.1425 ;
      RECT  111.1375 77.765 116.34 85.1425 ;
      RECT  109.475 85.1425 110.4375 85.62 ;
      RECT  111.1375 85.1425 116.34 85.62 ;
      RECT  109.475 85.62 110.4375 85.6875 ;
      RECT  109.475 85.6875 110.4375 87.6125 ;
      RECT  110.4375 85.6875 111.1375 87.6125 ;
      RECT  111.1375 85.62 125.14 85.6875 ;
      RECT  111.1375 85.6875 125.14 87.6125 ;
      RECT  12.605 21.0525 14.765 41.9175 ;
      RECT  12.605 41.9175 14.765 41.9825 ;
      RECT  14.765 21.0525 15.465 41.9175 ;
      RECT  15.465 21.0525 22.25 41.9175 ;
      RECT  15.465 41.9175 22.25 41.9825 ;
      RECT  12.605 41.9825 14.765 55.0325 ;
      RECT  12.605 55.0325 14.765 55.0975 ;
      RECT  14.765 55.0325 15.465 55.0975 ;
      RECT  15.465 41.9825 22.25 55.0325 ;
      RECT  15.465 55.0325 22.25 55.0975 ;
      RECT  1.1075 10.23 2.47 10.2625 ;
      RECT  1.1075 10.2625 2.47 18.3725 ;
      RECT  2.47 10.23 3.17 10.2625 ;
      RECT  1.1075 18.3725 2.47 21.0525 ;
      RECT  3.17 18.3725 14.625 21.0525 ;
      RECT  1.1075 21.0525 2.47 33.1925 ;
      RECT  3.17 21.0525 11.905 33.1925 ;
      RECT  1.1075 33.1925 2.47 33.225 ;
      RECT  1.1075 33.225 2.47 41.9825 ;
      RECT  2.47 33.225 3.17 41.9825 ;
      RECT  3.17 33.1925 11.905 33.225 ;
      RECT  3.17 33.225 11.905 41.9825 ;
      RECT  0.14 0.14 5.825 0.3825 ;
      RECT  0.14 0.3825 5.825 2.8525 ;
      RECT  5.825 0.14 6.525 0.3825 ;
      RECT  6.525 0.14 14.625 0.3825 ;
      RECT  6.525 0.3825 14.625 2.8525 ;
      RECT  1.1075 2.8525 5.825 10.23 ;
      RECT  6.525 2.8525 14.625 10.23 ;
      RECT  3.17 10.23 5.825 10.2625 ;
      RECT  6.525 10.23 14.625 10.2625 ;
      RECT  3.17 10.2625 5.825 15.9025 ;
      RECT  3.17 15.9025 5.825 18.3725 ;
      RECT  5.825 15.9025 6.525 18.3725 ;
      RECT  6.525 10.2625 14.625 15.9025 ;
      RECT  6.525 15.9025 14.625 18.3725 ;
      RECT  108.775 0.14 109.22 21.02 ;
      RECT  108.775 69.6625 109.22 75.04 ;
      RECT  109.22 0.14 109.475 21.02 ;
      RECT  109.22 21.02 109.475 69.6625 ;
      RECT  109.22 69.6625 109.475 75.04 ;
      RECT  107.63 21.0525 108.52 69.5925 ;
      RECT  107.63 69.5925 108.52 69.6625 ;
      RECT  107.07 21.02 108.52 21.0525 ;
      RECT  24.54 69.625 25.1 69.6625 ;
      RECT  25.1 69.5925 28.19 69.625 ;
      RECT  25.1 69.625 28.19 69.6625 ;
      RECT  25.1 21.0525 28.19 41.9825 ;
      RECT  25.1 41.9825 28.19 55.0975 ;
      RECT  25.1 55.0975 28.19 69.5925 ;
      RECT  22.95 21.02 24.4 21.0525 ;
      RECT  25.1 21.02 28.19 21.0525 ;
      RECT  30.43 17.8825 101.04 21.0525 ;
      RECT  30.43 69.5925 101.04 72.5125 ;
      RECT  30.43 21.0525 101.04 69.5925 ;
      RECT  109.475 8.6375 116.2 8.7025 ;
      RECT  109.475 8.7025 116.2 21.7525 ;
      RECT  116.2 8.6375 116.9 8.7025 ;
      RECT  116.9 8.6375 119.06 8.7025 ;
      RECT  116.9 8.7025 119.06 21.7525 ;
      RECT  109.475 21.7525 116.2 21.8175 ;
      RECT  109.475 21.8175 116.2 54.8025 ;
      RECT  116.2 21.8175 116.9 54.8025 ;
      RECT  116.9 21.7525 119.06 21.8175 ;
      RECT  116.9 21.8175 119.06 54.8025 ;
   END
END    freepdk45_sram_1w1r_14x128
END    LIBRARY
