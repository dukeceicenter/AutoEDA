VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_32x32_32
   CLASS BLOCK ;
   SIZE 112.245 BY 86.67 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.94 1.1075 21.075 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.8 1.1075 23.935 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.66 1.1075 26.795 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.52 1.1075 29.655 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.38 1.1075 32.515 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.24 1.1075 35.375 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.1 1.1075 38.235 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.96 1.1075 41.095 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.82 1.1075 43.955 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.68 1.1075 46.815 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.54 1.1075 49.675 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.4 1.1075 52.535 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.26 1.1075 55.395 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.12 1.1075 58.255 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.98 1.1075 61.115 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.84 1.1075 63.975 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.7 1.1075 66.835 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.56 1.1075 69.695 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.42 1.1075 72.555 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.28 1.1075 75.415 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.14 1.1075 78.275 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.0 1.1075 81.135 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.86 1.1075 83.995 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.72 1.1075 86.855 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.58 1.1075 89.715 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.44 1.1075 92.575 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.3 1.1075 95.435 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.16 1.1075 98.295 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.02 1.1075 101.155 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.88 1.1075 104.015 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.74 1.1075 106.875 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.6 1.1075 109.735 1.2425 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 42.7075 15.355 42.8425 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 45.4375 15.355 45.5725 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 47.6475 15.355 47.7825 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 50.3775 15.355 50.5125 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 52.5875 15.355 52.7225 ;
      END
   END addr0[4]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.41 19.5675 91.545 19.7025 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.41 16.8375 91.545 16.9725 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.41 14.6275 91.545 14.7625 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.41 11.8975 91.545 12.0325 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.41 9.6875 91.545 9.8225 ;
      END
   END addr1[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.485 85.4275 106.62 85.5625 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.3825 85.3425 100.5175 85.4775 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.4525 78.72 34.5875 78.855 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.6275 78.72 35.7625 78.855 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.8025 78.72 36.9375 78.855 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.9775 78.72 38.1125 78.855 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.1525 78.72 39.2875 78.855 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.3275 78.72 40.4625 78.855 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.5025 78.72 41.6375 78.855 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.6775 78.72 42.8125 78.855 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.8525 78.72 43.9875 78.855 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.0275 78.72 45.1625 78.855 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.2025 78.72 46.3375 78.855 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.3775 78.72 47.5125 78.855 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.5525 78.72 48.6875 78.855 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.7275 78.72 49.8625 78.855 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.9025 78.72 51.0375 78.855 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.0775 78.72 52.2125 78.855 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.2525 78.72 53.3875 78.855 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.4275 78.72 54.5625 78.855 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.6025 78.72 55.7375 78.855 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.7775 78.72 56.9125 78.855 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.9525 78.72 58.0875 78.855 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.1275 78.72 59.2625 78.855 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.3025 78.72 60.4375 78.855 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.4775 78.72 61.6125 78.855 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.6525 78.72 62.7875 78.855 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.8275 78.72 63.9625 78.855 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.0025 78.72 65.1375 78.855 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.1775 78.72 66.3125 78.855 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.3525 78.72 67.4875 78.855 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.5275 78.72 68.6625 78.855 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.7025 78.72 69.8375 78.855 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.8775 78.72 71.0125 78.855 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  31.2675 76.1625 71.6825 76.2325 ;
         LAYER metal4 ;
         RECT  106.0775 54.42 106.2175 76.8225 ;
         LAYER metal3 ;
         RECT  84.7725 22.1675 84.9075 22.3025 ;
         LAYER metal3 ;
         RECT  43.5375 2.4725 43.6725 2.6075 ;
         LAYER metal4 ;
         RECT  17.655 2.47 17.795 17.43 ;
         LAYER metal3 ;
         RECT  104.345 84.0625 104.48 84.1975 ;
         LAYER metal3 ;
         RECT  85.1175 31.1375 85.2525 31.2725 ;
         LAYER metal3 ;
         RECT  85.1175 37.1175 85.2525 37.2525 ;
         LAYER metal3 ;
         RECT  30.1225 19.1775 30.2575 19.3125 ;
         LAYER metal3 ;
         RECT  21.3175 37.1175 21.4525 37.2525 ;
         LAYER metal3 ;
         RECT  100.7375 2.4725 100.8725 2.6075 ;
         LAYER metal3 ;
         RECT  21.6625 22.1675 21.7975 22.3025 ;
         LAYER metal4 ;
         RECT  88.97 74.18 89.11 84.2 ;
         LAYER metal3 ;
         RECT  20.6575 2.4725 20.7925 2.6075 ;
         LAYER metal3 ;
         RECT  21.6625 25.1575 21.7975 25.2925 ;
         LAYER metal4 ;
         RECT  79.56 20.67 79.7 68.72 ;
         LAYER metal3 ;
         RECT  89.2975 2.4725 89.4325 2.6075 ;
         LAYER metal3 ;
         RECT  77.8575 2.4725 77.9925 2.6075 ;
         LAYER metal3 ;
         RECT  85.1175 40.1075 85.2525 40.2425 ;
         LAYER metal4 ;
         RECT  30.12 20.67 30.26 68.65 ;
         LAYER metal3 ;
         RECT  54.9775 2.4725 55.1125 2.6075 ;
         LAYER metal4 ;
         RECT  26.87 20.67 27.01 68.72 ;
         LAYER metal3 ;
         RECT  66.4175 2.4725 66.5525 2.6075 ;
         LAYER metal3 ;
         RECT  78.945 69.22 79.08 69.355 ;
         LAYER metal3 ;
         RECT  31.2675 72.265 73.3275 72.335 ;
         LAYER metal4 ;
         RECT  91.69 8.255 91.83 20.81 ;
         LAYER metal4 ;
         RECT  75.23 17.5 75.37 71.57 ;
         LAYER metal3 ;
         RECT  21.3175 40.1075 21.4525 40.2425 ;
         LAYER metal3 ;
         RECT  21.3175 34.1275 21.4525 34.2625 ;
         LAYER metal4 ;
         RECT  31.2 17.5 31.34 71.57 ;
         LAYER metal3 ;
         RECT  84.7725 25.1575 84.9075 25.2925 ;
         LAYER metal3 ;
         RECT  31.2675 11.37 71.6825 11.44 ;
         LAYER metal3 ;
         RECT  76.3125 70.0075 76.4475 70.1425 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal4 ;
         RECT  14.935 41.6 15.075 54.155 ;
         LAYER metal4 ;
         RECT  76.31 20.67 76.45 68.65 ;
         LAYER metal3 ;
         RECT  31.2675 16.805 72.1525 16.875 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
         LAYER metal3 ;
         RECT  32.0975 2.4725 32.2325 2.6075 ;
         LAYER metal3 ;
         RECT  21.3175 31.1375 21.4525 31.2725 ;
         LAYER metal3 ;
         RECT  85.1175 34.1275 85.2525 34.2625 ;
         LAYER metal3 ;
         RECT  27.49 19.965 27.625 20.1 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  74.77 17.5 74.91 71.57 ;
         LAYER metal3 ;
         RECT  86.3 26.6525 86.435 26.7875 ;
         LAYER metal4 ;
         RECT  100.52 71.71 100.66 86.67 ;
         LAYER metal3 ;
         RECT  86.925 29.6425 87.06 29.7775 ;
         LAYER metal3 ;
         RECT  31.2675 74.27 71.7175 74.34 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal3 ;
         RECT  20.135 20.6725 20.27 20.8075 ;
         LAYER metal3 ;
         RECT  57.8375 0.0025 57.9725 0.1375 ;
         LAYER metal4 ;
         RECT  31.66 17.5 31.8 71.57 ;
         LAYER metal3 ;
         RECT  19.51 35.6225 19.645 35.7575 ;
         LAYER metal3 ;
         RECT  86.925 32.6325 87.06 32.7675 ;
         LAYER metal3 ;
         RECT  69.2775 0.0025 69.4125 0.1375 ;
         LAYER metal4 ;
         RECT  81.15 20.6375 81.29 68.72 ;
         LAYER metal3 ;
         RECT  103.5975 0.0025 103.7325 0.1375 ;
         LAYER metal3 ;
         RECT  86.3 20.6725 86.435 20.8075 ;
         LAYER metal3 ;
         RECT  34.9575 0.0025 35.0925 0.1375 ;
         LAYER metal4 ;
         RECT  25.28 20.6375 25.42 68.72 ;
         LAYER metal3 ;
         RECT  19.51 29.6425 19.645 29.7775 ;
         LAYER metal3 ;
         RECT  92.1575 0.0025 92.2925 0.1375 ;
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal4 ;
         RECT  17.795 41.535 17.935 54.09 ;
         LAYER metal3 ;
         RECT  80.7175 0.0025 80.8525 0.1375 ;
         LAYER metal3 ;
         RECT  46.3975 0.0025 46.5325 0.1375 ;
         LAYER metal4 ;
         RECT  104.015 54.3875 104.155 76.79 ;
         LAYER metal3 ;
         RECT  19.51 32.6325 19.645 32.7675 ;
         LAYER metal3 ;
         RECT  86.925 38.6125 87.06 38.7475 ;
         LAYER metal3 ;
         RECT  104.345 86.5325 104.48 86.6675 ;
         LAYER metal4 ;
         RECT  88.83 8.32 88.97 20.875 ;
         LAYER metal3 ;
         RECT  20.135 26.6525 20.27 26.7875 ;
         LAYER metal3 ;
         RECT  23.5175 0.0025 23.6525 0.1375 ;
         LAYER metal4 ;
         RECT  79.0 20.6375 79.14 68.6825 ;
         LAYER metal3 ;
         RECT  86.925 35.6225 87.06 35.7575 ;
         LAYER metal3 ;
         RECT  19.51 38.6125 19.645 38.7475 ;
         LAYER metal3 ;
         RECT  20.135 23.6625 20.27 23.7975 ;
         LAYER metal3 ;
         RECT  86.925 41.6025 87.06 41.7375 ;
         LAYER metal3 ;
         RECT  31.2675 13.42 71.6825 13.49 ;
         LAYER metal3 ;
         RECT  86.3 23.6625 86.435 23.7975 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal3 ;
         RECT  19.51 41.6025 19.645 41.7375 ;
         LAYER metal4 ;
         RECT  27.43 20.6375 27.57 68.6825 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 112.105 86.53 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 112.105 86.53 ;
   LAYER  metal3 ;
      RECT  20.8 0.14 21.215 0.9675 ;
      RECT  21.215 0.9675 23.66 1.3825 ;
      RECT  24.075 0.9675 26.52 1.3825 ;
      RECT  26.935 0.9675 29.38 1.3825 ;
      RECT  29.795 0.9675 32.24 1.3825 ;
      RECT  32.655 0.9675 35.1 1.3825 ;
      RECT  35.515 0.9675 37.96 1.3825 ;
      RECT  38.375 0.9675 40.82 1.3825 ;
      RECT  41.235 0.9675 43.68 1.3825 ;
      RECT  44.095 0.9675 46.54 1.3825 ;
      RECT  46.955 0.9675 49.4 1.3825 ;
      RECT  49.815 0.9675 52.26 1.3825 ;
      RECT  52.675 0.9675 55.12 1.3825 ;
      RECT  55.535 0.9675 57.98 1.3825 ;
      RECT  58.395 0.9675 60.84 1.3825 ;
      RECT  61.255 0.9675 63.7 1.3825 ;
      RECT  64.115 0.9675 66.56 1.3825 ;
      RECT  66.975 0.9675 69.42 1.3825 ;
      RECT  69.835 0.9675 72.28 1.3825 ;
      RECT  72.695 0.9675 75.14 1.3825 ;
      RECT  75.555 0.9675 78.0 1.3825 ;
      RECT  78.415 0.9675 80.86 1.3825 ;
      RECT  81.275 0.9675 83.72 1.3825 ;
      RECT  84.135 0.9675 86.58 1.3825 ;
      RECT  86.995 0.9675 89.44 1.3825 ;
      RECT  89.855 0.9675 92.3 1.3825 ;
      RECT  92.715 0.9675 95.16 1.3825 ;
      RECT  95.575 0.9675 98.02 1.3825 ;
      RECT  98.435 0.9675 100.88 1.3825 ;
      RECT  101.295 0.9675 103.74 1.3825 ;
      RECT  104.155 0.9675 106.6 1.3825 ;
      RECT  107.015 0.9675 109.46 1.3825 ;
      RECT  109.875 0.9675 112.105 1.3825 ;
      RECT  0.14 42.5675 15.08 42.9825 ;
      RECT  0.14 42.9825 15.08 86.53 ;
      RECT  15.08 1.3825 15.495 42.5675 ;
      RECT  15.495 42.5675 20.8 42.9825 ;
      RECT  15.495 42.9825 20.8 86.53 ;
      RECT  15.08 42.9825 15.495 45.2975 ;
      RECT  15.08 45.7125 15.495 47.5075 ;
      RECT  15.08 47.9225 15.495 50.2375 ;
      RECT  15.08 50.6525 15.495 52.4475 ;
      RECT  15.08 52.8625 15.495 86.53 ;
      RECT  91.27 19.8425 91.685 86.53 ;
      RECT  91.685 19.4275 112.105 19.8425 ;
      RECT  91.27 17.1125 91.685 19.4275 ;
      RECT  91.27 14.9025 91.685 16.6975 ;
      RECT  91.27 12.1725 91.685 14.4875 ;
      RECT  91.27 1.3825 91.685 9.5475 ;
      RECT  91.27 9.9625 91.685 11.7575 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  106.345 19.8425 106.76 85.2875 ;
      RECT  106.345 85.7025 106.76 86.53 ;
      RECT  106.76 19.8425 112.105 85.2875 ;
      RECT  106.76 85.2875 112.105 85.7025 ;
      RECT  106.76 85.7025 112.105 86.53 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 42.5675 ;
      RECT  6.5225 1.3825 15.08 1.4675 ;
      RECT  6.5225 1.4675 15.08 42.5675 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 20.8 1.0525 ;
      RECT  6.5225 1.0525 20.8 1.3825 ;
      RECT  91.685 19.8425 100.2425 85.2025 ;
      RECT  91.685 85.2025 100.2425 85.2875 ;
      RECT  100.2425 19.8425 100.6575 85.2025 ;
      RECT  100.6575 85.2025 106.345 85.2875 ;
      RECT  91.685 85.2875 100.2425 85.6175 ;
      RECT  91.685 85.6175 100.2425 85.7025 ;
      RECT  100.2425 85.6175 100.6575 85.7025 ;
      RECT  100.6575 85.2875 106.345 85.6175 ;
      RECT  100.6575 85.6175 106.345 85.7025 ;
      RECT  21.215 78.58 34.3125 78.995 ;
      RECT  21.215 78.995 34.3125 86.53 ;
      RECT  34.3125 78.995 34.7275 86.53 ;
      RECT  34.7275 78.995 91.27 86.53 ;
      RECT  34.7275 78.58 35.4875 78.995 ;
      RECT  35.9025 78.58 36.6625 78.995 ;
      RECT  37.0775 78.58 37.8375 78.995 ;
      RECT  38.2525 78.58 39.0125 78.995 ;
      RECT  39.4275 78.58 40.1875 78.995 ;
      RECT  40.6025 78.58 41.3625 78.995 ;
      RECT  41.7775 78.58 42.5375 78.995 ;
      RECT  42.9525 78.58 43.7125 78.995 ;
      RECT  44.1275 78.58 44.8875 78.995 ;
      RECT  45.3025 78.58 46.0625 78.995 ;
      RECT  46.4775 78.58 47.2375 78.995 ;
      RECT  47.6525 78.58 48.4125 78.995 ;
      RECT  48.8275 78.58 49.5875 78.995 ;
      RECT  50.0025 78.58 50.7625 78.995 ;
      RECT  51.1775 78.58 51.9375 78.995 ;
      RECT  52.3525 78.58 53.1125 78.995 ;
      RECT  53.5275 78.58 54.2875 78.995 ;
      RECT  54.7025 78.58 55.4625 78.995 ;
      RECT  55.8775 78.58 56.6375 78.995 ;
      RECT  57.0525 78.58 57.8125 78.995 ;
      RECT  58.2275 78.58 58.9875 78.995 ;
      RECT  59.4025 78.58 60.1625 78.995 ;
      RECT  60.5775 78.58 61.3375 78.995 ;
      RECT  61.7525 78.58 62.5125 78.995 ;
      RECT  62.9275 78.58 63.6875 78.995 ;
      RECT  64.1025 78.58 64.8625 78.995 ;
      RECT  65.2775 78.58 66.0375 78.995 ;
      RECT  66.4525 78.58 67.2125 78.995 ;
      RECT  67.6275 78.58 68.3875 78.995 ;
      RECT  68.8025 78.58 69.5625 78.995 ;
      RECT  69.9775 78.58 70.7375 78.995 ;
      RECT  71.1525 78.58 91.27 78.995 ;
      RECT  21.215 76.0225 31.1275 76.3725 ;
      RECT  21.215 76.3725 31.1275 78.58 ;
      RECT  31.1275 76.3725 34.3125 78.58 ;
      RECT  34.3125 76.3725 34.7275 78.58 ;
      RECT  34.7275 76.3725 71.8225 78.58 ;
      RECT  71.8225 76.0225 91.27 76.3725 ;
      RECT  71.8225 76.3725 91.27 78.58 ;
      RECT  71.8225 19.8425 84.6325 22.0275 ;
      RECT  71.8225 22.0275 84.6325 22.4425 ;
      RECT  84.6325 19.8425 85.0475 22.0275 ;
      RECT  85.0475 22.0275 91.27 22.4425 ;
      RECT  21.215 1.3825 43.3975 2.3325 ;
      RECT  43.3975 1.3825 43.8125 2.3325 ;
      RECT  43.8125 1.3825 91.27 2.3325 ;
      RECT  100.6575 19.8425 104.205 83.9225 ;
      RECT  100.6575 83.9225 104.205 84.3375 ;
      RECT  100.6575 84.3375 104.205 85.2025 ;
      RECT  104.205 19.8425 104.62 83.9225 ;
      RECT  104.205 84.3375 104.62 85.2025 ;
      RECT  104.62 19.8425 106.345 83.9225 ;
      RECT  104.62 83.9225 106.345 84.3375 ;
      RECT  104.62 84.3375 106.345 85.2025 ;
      RECT  84.6325 30.9975 84.9775 31.4125 ;
      RECT  84.6325 31.4125 84.9775 76.0225 ;
      RECT  85.0475 22.4425 85.3925 30.9975 ;
      RECT  85.3925 30.9975 91.27 31.4125 ;
      RECT  21.215 19.4275 29.9825 19.4525 ;
      RECT  29.9825 19.4525 30.3975 19.8425 ;
      RECT  30.3975 19.4275 91.27 19.4525 ;
      RECT  30.3975 19.4525 91.27 19.8425 ;
      RECT  21.215 2.7475 29.9825 19.0375 ;
      RECT  21.215 19.0375 29.9825 19.4275 ;
      RECT  29.9825 2.7475 30.3975 19.0375 ;
      RECT  30.3975 19.0375 43.3975 19.4275 ;
      RECT  20.8 36.9775 21.1775 37.3925 ;
      RECT  20.8 37.3925 21.1775 86.53 ;
      RECT  21.5925 36.9775 31.1275 37.3925 ;
      RECT  21.5925 37.3925 31.1275 76.0225 ;
      RECT  91.685 1.3825 100.5975 2.3325 ;
      RECT  91.685 2.3325 100.5975 2.7475 ;
      RECT  91.685 2.7475 100.5975 19.4275 ;
      RECT  100.5975 1.3825 101.0125 2.3325 ;
      RECT  100.5975 2.7475 101.0125 19.4275 ;
      RECT  101.0125 1.3825 112.105 2.3325 ;
      RECT  101.0125 2.3325 112.105 2.7475 ;
      RECT  101.0125 2.7475 112.105 19.4275 ;
      RECT  21.215 19.8425 21.5225 22.0275 ;
      RECT  21.215 22.0275 21.5225 22.4425 ;
      RECT  21.5225 19.8425 21.5925 22.0275 ;
      RECT  21.5925 19.8425 21.9375 22.0275 ;
      RECT  21.9375 22.0275 31.1275 22.4425 ;
      RECT  21.9375 22.4425 31.1275 36.9775 ;
      RECT  15.495 1.3825 20.5175 2.3325 ;
      RECT  15.495 2.3325 20.5175 2.7475 ;
      RECT  20.5175 1.3825 20.8 2.3325 ;
      RECT  20.5175 2.7475 20.8 42.5675 ;
      RECT  20.8 1.3825 20.9325 2.3325 ;
      RECT  20.8 2.7475 20.9325 36.9775 ;
      RECT  20.9325 1.3825 21.1775 2.3325 ;
      RECT  20.9325 2.3325 21.1775 2.7475 ;
      RECT  20.9325 2.7475 21.1775 36.9775 ;
      RECT  21.5225 22.4425 21.5925 25.0175 ;
      RECT  21.5925 22.4425 21.9375 25.0175 ;
      RECT  21.5925 25.4325 21.9375 36.9775 ;
      RECT  89.5725 2.3325 91.27 2.7475 ;
      RECT  78.1325 2.3325 89.1575 2.7475 ;
      RECT  84.9775 37.3925 85.0475 39.9675 ;
      RECT  84.9775 40.3825 85.0475 76.0225 ;
      RECT  85.0475 37.3925 85.3925 39.9675 ;
      RECT  85.0475 40.3825 85.3925 76.0225 ;
      RECT  43.8125 2.3325 54.8375 2.7475 ;
      RECT  55.2525 2.3325 66.2775 2.7475 ;
      RECT  66.6925 2.3325 77.7175 2.7475 ;
      RECT  71.8225 22.4425 78.805 69.08 ;
      RECT  71.8225 69.08 78.805 69.495 ;
      RECT  78.805 22.4425 79.22 69.08 ;
      RECT  78.805 69.495 79.22 76.0225 ;
      RECT  79.22 22.4425 84.6325 69.08 ;
      RECT  79.22 69.08 84.6325 69.495 ;
      RECT  79.22 69.495 84.6325 76.0225 ;
      RECT  31.1275 19.8425 34.3125 72.125 ;
      RECT  34.3125 19.8425 34.7275 72.125 ;
      RECT  34.7275 19.8425 71.8225 72.125 ;
      RECT  71.8225 69.495 73.4675 72.125 ;
      RECT  73.4675 72.125 78.805 72.475 ;
      RECT  73.4675 72.475 78.805 76.0225 ;
      RECT  21.1775 37.3925 21.215 39.9675 ;
      RECT  21.1775 40.3825 21.215 86.53 ;
      RECT  21.215 37.3925 21.5925 39.9675 ;
      RECT  21.215 40.3825 21.5925 76.0225 ;
      RECT  21.1775 34.4025 21.215 36.9775 ;
      RECT  21.215 34.4025 21.5225 36.9775 ;
      RECT  21.5225 34.4025 21.5925 36.9775 ;
      RECT  84.6325 22.4425 84.9775 25.0175 ;
      RECT  84.6325 25.4325 84.9775 30.9975 ;
      RECT  84.9775 22.4425 85.0475 25.0175 ;
      RECT  84.9775 25.4325 85.0475 30.9975 ;
      RECT  43.3975 2.7475 43.8125 11.23 ;
      RECT  43.8125 2.7475 71.8225 11.23 ;
      RECT  71.8225 2.7475 91.27 11.23 ;
      RECT  71.8225 11.23 91.27 11.58 ;
      RECT  30.3975 2.7475 31.1275 11.23 ;
      RECT  30.3975 11.23 31.1275 11.58 ;
      RECT  30.3975 11.58 31.1275 19.0375 ;
      RECT  31.1275 2.7475 43.3975 11.23 ;
      RECT  73.4675 69.495 76.1725 69.8675 ;
      RECT  73.4675 69.8675 76.1725 70.2825 ;
      RECT  73.4675 70.2825 76.1725 72.125 ;
      RECT  76.1725 69.495 76.5875 69.8675 ;
      RECT  76.1725 70.2825 76.5875 72.125 ;
      RECT  76.5875 69.495 78.805 69.8675 ;
      RECT  76.5875 69.8675 78.805 70.2825 ;
      RECT  76.5875 70.2825 78.805 72.125 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 42.5675 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 42.5675 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 42.5675 ;
      RECT  43.3975 17.015 43.8125 19.4275 ;
      RECT  43.8125 17.015 71.8225 19.4275 ;
      RECT  71.8225 11.58 72.2925 16.665 ;
      RECT  71.8225 17.015 72.2925 19.4275 ;
      RECT  72.2925 11.58 91.27 16.665 ;
      RECT  72.2925 16.665 91.27 17.015 ;
      RECT  72.2925 17.015 91.27 19.4275 ;
      RECT  31.1275 17.015 43.3975 19.0375 ;
      RECT  21.215 2.3325 31.9575 2.7475 ;
      RECT  32.3725 2.3325 43.3975 2.7475 ;
      RECT  21.1775 1.3825 21.215 30.9975 ;
      RECT  21.1775 31.4125 21.215 33.9875 ;
      RECT  21.215 22.4425 21.5225 30.9975 ;
      RECT  21.215 31.4125 21.5225 33.9875 ;
      RECT  21.5225 25.4325 21.5925 30.9975 ;
      RECT  21.5225 31.4125 21.5925 33.9875 ;
      RECT  84.9775 31.4125 85.0475 33.9875 ;
      RECT  84.9775 34.4025 85.0475 36.9775 ;
      RECT  85.0475 31.4125 85.3925 33.9875 ;
      RECT  85.0475 34.4025 85.3925 36.9775 ;
      RECT  21.215 19.4525 27.35 19.825 ;
      RECT  21.215 19.825 27.35 19.8425 ;
      RECT  27.35 19.4525 27.765 19.825 ;
      RECT  27.765 19.4525 29.9825 19.825 ;
      RECT  27.765 19.825 29.9825 19.8425 ;
      RECT  21.9375 19.8425 27.35 20.24 ;
      RECT  21.9375 20.24 27.35 22.0275 ;
      RECT  27.35 20.24 27.765 22.0275 ;
      RECT  27.765 19.8425 31.1275 20.24 ;
      RECT  27.765 20.24 31.1275 22.0275 ;
      RECT  85.3925 22.4425 86.16 26.5125 ;
      RECT  85.3925 26.5125 86.16 26.9275 ;
      RECT  85.3925 26.9275 86.16 30.9975 ;
      RECT  86.16 26.9275 86.575 30.9975 ;
      RECT  86.575 22.4425 91.27 26.5125 ;
      RECT  86.575 26.5125 91.27 26.9275 ;
      RECT  86.575 26.9275 86.785 29.5025 ;
      RECT  86.575 29.5025 86.785 29.9175 ;
      RECT  86.575 29.9175 86.785 30.9975 ;
      RECT  86.785 26.9275 87.2 29.5025 ;
      RECT  86.785 29.9175 87.2 30.9975 ;
      RECT  87.2 26.9275 91.27 29.5025 ;
      RECT  87.2 29.5025 91.27 29.9175 ;
      RECT  87.2 29.9175 91.27 30.9975 ;
      RECT  31.1275 72.475 34.3125 74.13 ;
      RECT  31.1275 74.48 34.3125 76.0225 ;
      RECT  34.3125 72.475 34.7275 74.13 ;
      RECT  34.3125 74.48 34.7275 76.0225 ;
      RECT  34.7275 72.475 71.8225 74.13 ;
      RECT  34.7275 74.48 71.8225 76.0225 ;
      RECT  71.8225 72.475 71.8575 74.13 ;
      RECT  71.8225 74.48 71.8575 76.0225 ;
      RECT  71.8575 72.475 73.4675 74.13 ;
      RECT  71.8575 74.13 73.4675 74.48 ;
      RECT  71.8575 74.48 73.4675 76.0225 ;
      RECT  15.495 2.7475 19.995 20.5325 ;
      RECT  15.495 20.5325 19.995 20.9475 ;
      RECT  19.995 2.7475 20.41 20.5325 ;
      RECT  20.41 2.7475 20.5175 20.5325 ;
      RECT  20.41 20.5325 20.5175 20.9475 ;
      RECT  20.41 20.9475 20.5175 42.5675 ;
      RECT  21.215 0.2775 57.6975 0.9675 ;
      RECT  57.6975 0.2775 58.1125 0.9675 ;
      RECT  58.1125 0.2775 112.105 0.9675 ;
      RECT  15.495 20.9475 19.37 35.4825 ;
      RECT  15.495 35.4825 19.37 35.8975 ;
      RECT  15.495 35.8975 19.37 42.5675 ;
      RECT  19.785 20.9475 19.995 35.4825 ;
      RECT  19.785 35.4825 19.995 35.8975 ;
      RECT  19.785 35.8975 19.995 42.5675 ;
      RECT  85.3925 31.4125 86.785 32.4925 ;
      RECT  85.3925 32.4925 86.785 32.9075 ;
      RECT  85.3925 32.9075 86.785 76.0225 ;
      RECT  86.785 31.4125 87.2 32.4925 ;
      RECT  87.2 31.4125 91.27 32.4925 ;
      RECT  87.2 32.4925 91.27 32.9075 ;
      RECT  87.2 32.9075 91.27 76.0225 ;
      RECT  58.1125 0.14 69.1375 0.2775 ;
      RECT  103.8725 0.14 112.105 0.2775 ;
      RECT  85.0475 19.8425 86.16 20.5325 ;
      RECT  85.0475 20.5325 86.16 20.9475 ;
      RECT  85.0475 20.9475 86.16 22.0275 ;
      RECT  86.16 19.8425 86.575 20.5325 ;
      RECT  86.16 20.9475 86.575 22.0275 ;
      RECT  86.575 19.8425 91.27 20.5325 ;
      RECT  86.575 20.5325 91.27 20.9475 ;
      RECT  86.575 20.9475 91.27 22.0275 ;
      RECT  19.37 20.9475 19.785 29.5025 ;
      RECT  92.4325 0.14 103.4575 0.2775 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  0.14 0.2775 2.285 0.9675 ;
      RECT  2.285 0.2775 2.7 0.9675 ;
      RECT  2.7 0.14 20.8 0.2775 ;
      RECT  2.7 0.2775 20.8 0.9675 ;
      RECT  69.5525 0.14 80.5775 0.2775 ;
      RECT  80.9925 0.14 92.0175 0.2775 ;
      RECT  35.2325 0.14 46.2575 0.2775 ;
      RECT  46.6725 0.14 57.6975 0.2775 ;
      RECT  19.37 29.9175 19.785 32.4925 ;
      RECT  19.37 32.9075 19.785 35.4825 ;
      RECT  91.685 85.7025 104.205 86.3925 ;
      RECT  91.685 86.3925 104.205 86.53 ;
      RECT  104.205 85.7025 104.62 86.3925 ;
      RECT  104.62 85.7025 106.345 86.3925 ;
      RECT  104.62 86.3925 106.345 86.53 ;
      RECT  19.995 26.9275 20.41 42.5675 ;
      RECT  21.215 0.14 23.3775 0.2775 ;
      RECT  23.7925 0.14 34.8175 0.2775 ;
      RECT  86.785 32.9075 87.2 35.4825 ;
      RECT  86.785 35.8975 87.2 38.4725 ;
      RECT  19.37 35.8975 19.785 38.4725 ;
      RECT  19.995 20.9475 20.41 23.5225 ;
      RECT  19.995 23.9375 20.41 26.5125 ;
      RECT  86.785 38.8875 87.2 41.4625 ;
      RECT  86.785 41.8775 87.2 76.0225 ;
      RECT  43.3975 11.58 43.8125 13.28 ;
      RECT  43.3975 13.63 43.8125 16.665 ;
      RECT  43.8125 11.58 71.8225 13.28 ;
      RECT  43.8125 13.63 71.8225 16.665 ;
      RECT  31.1275 11.58 43.3975 13.28 ;
      RECT  31.1275 13.63 43.3975 16.665 ;
      RECT  86.16 22.4425 86.575 23.5225 ;
      RECT  86.16 23.9375 86.575 26.5125 ;
      RECT  19.37 38.8875 19.785 41.4625 ;
      RECT  19.37 41.8775 19.785 42.5675 ;
   LAYER  metal4 ;
      RECT  105.7975 0.14 106.4975 54.14 ;
      RECT  105.7975 77.1025 106.4975 86.53 ;
      RECT  106.4975 0.14 112.105 54.14 ;
      RECT  106.4975 54.14 112.105 77.1025 ;
      RECT  106.4975 77.1025 112.105 86.53 ;
      RECT  17.375 0.14 18.075 2.19 ;
      RECT  18.075 0.14 105.7975 2.19 ;
      RECT  0.14 73.9 88.69 77.1025 ;
      RECT  88.69 54.14 89.39 73.9 ;
      RECT  0.14 77.1025 88.69 84.48 ;
      RECT  0.14 84.48 88.69 86.53 ;
      RECT  88.69 84.48 89.39 86.53 ;
      RECT  79.28 69.0 79.98 73.9 ;
      RECT  79.98 69.0 88.69 73.9 ;
      RECT  29.84 68.93 30.54 69.0 ;
      RECT  18.075 2.19 91.41 7.975 ;
      RECT  91.41 2.19 92.11 7.975 ;
      RECT  92.11 2.19 105.7975 7.975 ;
      RECT  92.11 7.975 105.7975 17.71 ;
      RECT  92.11 17.71 105.7975 20.39 ;
      RECT  91.41 21.09 92.11 54.14 ;
      RECT  92.11 20.39 105.7975 21.09 ;
      RECT  0.14 71.85 74.95 73.9 ;
      RECT  74.95 71.85 75.65 73.9 ;
      RECT  75.65 69.0 79.28 71.85 ;
      RECT  75.65 71.85 79.28 73.9 ;
      RECT  18.075 7.975 74.95 17.22 ;
      RECT  74.95 7.975 75.65 17.22 ;
      RECT  0.14 69.0 30.92 71.85 ;
      RECT  30.54 20.39 30.92 54.14 ;
      RECT  30.54 54.14 30.92 68.93 ;
      RECT  30.54 68.93 30.92 69.0 ;
      RECT  18.075 17.22 30.92 17.71 ;
      RECT  0.14 41.32 14.655 54.14 ;
      RECT  14.655 17.71 15.355 41.32 ;
      RECT  15.355 17.71 17.375 41.32 ;
      RECT  15.355 41.32 17.375 54.14 ;
      RECT  0.14 54.14 14.655 54.435 ;
      RECT  0.14 54.435 14.655 68.93 ;
      RECT  14.655 54.435 15.355 68.93 ;
      RECT  75.65 20.39 76.03 54.14 ;
      RECT  75.65 54.14 76.03 68.93 ;
      RECT  0.14 2.19 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 17.71 ;
      RECT  0.4075 2.19 1.1075 9.5675 ;
      RECT  0.14 17.71 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 41.32 ;
      RECT  0.4075 32.53 1.1075 41.32 ;
      RECT  89.39 54.14 100.24 71.43 ;
      RECT  89.39 71.43 100.24 73.9 ;
      RECT  100.24 54.14 100.94 71.43 ;
      RECT  89.39 73.9 100.24 77.1025 ;
      RECT  89.39 77.1025 100.24 84.48 ;
      RECT  100.94 77.1025 105.7975 84.48 ;
      RECT  89.39 84.48 100.24 86.53 ;
      RECT  100.94 84.48 105.7975 86.53 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 17.71 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  1.1075 17.71 2.47 32.53 ;
      RECT  3.17 17.71 14.655 32.53 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 41.32 ;
      RECT  2.47 32.5625 3.17 41.32 ;
      RECT  3.17 32.53 14.655 32.5625 ;
      RECT  3.17 32.5625 14.655 41.32 ;
      RECT  32.08 17.71 74.49 20.39 ;
      RECT  32.08 69.0 74.49 71.85 ;
      RECT  32.08 20.39 74.49 54.14 ;
      RECT  32.08 54.14 74.49 68.93 ;
      RECT  32.08 68.93 74.49 69.0 ;
      RECT  32.08 17.22 74.49 17.71 ;
      RECT  79.98 54.14 80.87 69.0 ;
      RECT  81.57 54.14 88.69 69.0 ;
      RECT  79.98 17.71 80.87 20.3575 ;
      RECT  79.98 20.3575 80.87 20.39 ;
      RECT  80.87 17.71 81.57 20.3575 ;
      RECT  79.98 20.39 80.87 21.09 ;
      RECT  79.98 21.09 80.87 54.14 ;
      RECT  25.7 20.39 26.59 54.14 ;
      RECT  0.14 68.93 25.0 69.0 ;
      RECT  25.7 68.93 26.59 69.0 ;
      RECT  18.075 17.71 25.0 20.3575 ;
      RECT  18.075 20.3575 25.0 20.39 ;
      RECT  25.0 17.71 25.7 20.3575 ;
      RECT  25.7 17.71 30.92 20.3575 ;
      RECT  25.7 54.14 26.59 54.435 ;
      RECT  15.355 54.435 25.0 68.93 ;
      RECT  25.7 54.435 26.59 68.93 ;
      RECT  17.375 17.71 17.515 41.255 ;
      RECT  17.375 41.255 17.515 54.14 ;
      RECT  17.515 17.71 18.075 41.255 ;
      RECT  18.075 20.39 18.215 41.255 ;
      RECT  18.215 20.39 25.0 41.255 ;
      RECT  18.215 41.255 25.0 54.14 ;
      RECT  15.355 54.14 17.515 54.37 ;
      RECT  15.355 54.37 17.515 54.435 ;
      RECT  17.515 54.37 18.215 54.435 ;
      RECT  18.215 54.14 25.0 54.37 ;
      RECT  18.215 54.37 25.0 54.435 ;
      RECT  92.11 21.09 103.735 54.1075 ;
      RECT  92.11 54.1075 103.735 54.14 ;
      RECT  103.735 21.09 104.435 54.1075 ;
      RECT  104.435 21.09 105.7975 54.1075 ;
      RECT  104.435 54.1075 105.7975 54.14 ;
      RECT  100.94 54.14 103.735 71.43 ;
      RECT  104.435 54.14 105.7975 71.43 ;
      RECT  100.94 71.43 103.735 73.9 ;
      RECT  104.435 71.43 105.7975 73.9 ;
      RECT  100.94 73.9 103.735 77.07 ;
      RECT  100.94 77.07 103.735 77.1025 ;
      RECT  103.735 77.07 104.435 77.1025 ;
      RECT  104.435 73.9 105.7975 77.07 ;
      RECT  104.435 77.07 105.7975 77.1025 ;
      RECT  75.65 7.975 88.55 8.04 ;
      RECT  75.65 8.04 88.55 17.22 ;
      RECT  88.55 7.975 89.25 8.04 ;
      RECT  89.25 7.975 91.41 8.04 ;
      RECT  89.25 8.04 91.41 17.22 ;
      RECT  75.65 17.22 88.55 17.71 ;
      RECT  89.25 17.22 91.41 17.71 ;
      RECT  81.57 17.71 88.55 20.3575 ;
      RECT  89.25 17.71 91.41 20.3575 ;
      RECT  81.57 20.3575 88.55 20.39 ;
      RECT  89.25 20.3575 91.41 20.39 ;
      RECT  81.57 20.39 88.55 21.09 ;
      RECT  89.25 20.39 91.41 21.09 ;
      RECT  81.57 21.09 88.55 21.155 ;
      RECT  81.57 21.155 88.55 54.14 ;
      RECT  88.55 21.155 89.25 54.14 ;
      RECT  89.25 21.09 91.41 21.155 ;
      RECT  89.25 21.155 91.41 54.14 ;
      RECT  79.28 17.71 79.42 20.3575 ;
      RECT  79.42 17.71 79.98 20.3575 ;
      RECT  79.42 20.3575 79.98 20.39 ;
      RECT  75.65 17.71 78.72 20.3575 ;
      RECT  75.65 20.3575 78.72 20.39 ;
      RECT  78.72 17.71 79.28 20.3575 ;
      RECT  75.65 68.93 78.72 68.9625 ;
      RECT  75.65 68.9625 78.72 69.0 ;
      RECT  78.72 68.9625 79.28 69.0 ;
      RECT  76.73 20.39 78.72 54.14 ;
      RECT  76.73 54.14 78.72 68.93 ;
      RECT  0.14 0.14 5.825 2.19 ;
      RECT  6.525 0.14 17.375 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 17.375 9.5675 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  6.525 9.5675 17.375 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  3.17 15.24 5.825 17.71 ;
      RECT  5.825 15.24 6.525 17.71 ;
      RECT  6.525 9.6 17.375 15.24 ;
      RECT  6.525 15.24 17.375 17.71 ;
      RECT  27.85 20.39 29.84 54.14 ;
      RECT  27.85 54.14 29.84 68.93 ;
      RECT  27.29 68.9625 27.85 69.0 ;
      RECT  27.85 68.93 29.84 68.9625 ;
      RECT  27.85 68.9625 29.84 69.0 ;
      RECT  25.7 20.3575 27.15 20.39 ;
      RECT  27.85 20.3575 30.92 20.39 ;
   END
END    freepdk45_sram_1w1r_32x32_32
END    LIBRARY
