VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_64x32_32
   CLASS BLOCK ;
   SIZE 147.255 BY 86.67 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.8 1.1075 23.935 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.66 1.1075 26.795 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.52 1.1075 29.655 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.38 1.1075 32.515 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.24 1.1075 35.375 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.1 1.1075 38.235 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.96 1.1075 41.095 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.82 1.1075 43.955 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.68 1.1075 46.815 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.54 1.1075 49.675 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.4 1.1075 52.535 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.26 1.1075 55.395 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.12 1.1075 58.255 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.98 1.1075 61.115 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.84 1.1075 63.975 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.7 1.1075 66.835 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.56 1.1075 69.695 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.42 1.1075 72.555 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.28 1.1075 75.415 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.14 1.1075 78.275 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.0 1.1075 81.135 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.86 1.1075 83.995 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.72 1.1075 86.855 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.58 1.1075 89.715 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.44 1.1075 92.575 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.3 1.1075 95.435 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.16 1.1075 98.295 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.02 1.1075 101.155 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.88 1.1075 104.015 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.74 1.1075 106.875 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.6 1.1075 109.735 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.46 1.1075 112.595 1.2425 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.94 1.1075 21.075 1.2425 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 42.7075 15.355 42.8425 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 45.4375 15.355 45.5725 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 47.6475 15.355 47.7825 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 50.3775 15.355 50.5125 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 52.5875 15.355 52.7225 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.18 84.1625 123.315 84.2975 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.76 19.5675 131.895 19.7025 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.76 16.8375 131.895 16.9725 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.76 14.6275 131.895 14.7625 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.76 11.8975 131.895 12.0325 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.76 9.6875 131.895 9.8225 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.835 85.4275 146.97 85.5625 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.7325 85.3425 140.8675 85.4775 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.8275 81.675 35.9625 81.81 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.1775 81.675 38.3125 81.81 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.5275 81.675 40.6625 81.81 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.8775 81.675 43.0125 81.81 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.2275 81.675 45.3625 81.81 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.5775 81.675 47.7125 81.81 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.9275 81.675 50.0625 81.81 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.2775 81.675 52.4125 81.81 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.6275 81.675 54.7625 81.81 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.9775 81.675 57.1125 81.81 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.3275 81.675 59.4625 81.81 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.6775 81.675 61.8125 81.81 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.0275 81.675 64.1625 81.81 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.3775 81.675 66.5125 81.81 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.7275 81.675 68.8625 81.81 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.0775 81.675 71.2125 81.81 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.4275 81.675 73.5625 81.81 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.7775 81.675 75.9125 81.81 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.1275 81.675 78.2625 81.81 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.4775 81.675 80.6125 81.81 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.8275 81.675 82.9625 81.81 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.1775 81.675 85.3125 81.81 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.5275 81.675 87.6625 81.81 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.8775 81.675 90.0125 81.81 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.2275 81.675 92.3625 81.81 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.5775 81.675 94.7125 81.81 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.9275 81.675 97.0625 81.81 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.2775 81.675 99.4125 81.81 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.6275 81.675 101.7625 81.81 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.9775 81.675 104.1125 81.81 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.3275 81.675 106.4625 81.81 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.6775 81.675 108.8125 81.81 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  31.495 20.67 31.635 68.65 ;
         LAYER metal4 ;
         RECT  26.87 20.67 27.01 68.72 ;
         LAYER metal3 ;
         RECT  32.6425 16.805 111.1275 16.875 ;
         LAYER metal3 ;
         RECT  125.1225 25.1575 125.2575 25.2925 ;
         LAYER metal3 ;
         RECT  121.205 77.0975 121.34 77.2325 ;
         LAYER metal3 ;
         RECT  125.4675 34.1275 125.6025 34.2625 ;
         LAYER metal4 ;
         RECT  129.32 74.18 129.46 84.2 ;
         LAYER metal4 ;
         RECT  14.935 41.6 15.075 54.155 ;
         LAYER metal3 ;
         RECT  92.1575 2.4725 92.2925 2.6075 ;
         LAYER metal4 ;
         RECT  114.205 17.5 114.345 71.57 ;
         LAYER metal4 ;
         RECT  115.285 20.67 115.425 68.65 ;
         LAYER metal3 ;
         RECT  103.5975 2.4725 103.7325 2.6075 ;
         LAYER metal3 ;
         RECT  125.1225 22.1675 125.2575 22.3025 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
         LAYER metal3 ;
         RECT  144.695 84.0625 144.83 84.1975 ;
         LAYER metal3 ;
         RECT  46.3975 2.4725 46.5325 2.6075 ;
         LAYER metal3 ;
         RECT  125.4675 40.1075 125.6025 40.2425 ;
         LAYER metal3 ;
         RECT  123.4625 82.7975 123.5975 82.9325 ;
         LAYER metal3 ;
         RECT  125.4675 37.1175 125.6025 37.2525 ;
         LAYER metal3 ;
         RECT  57.8375 2.4725 57.9725 2.6075 ;
         LAYER metal3 ;
         RECT  21.3175 31.1375 21.4525 31.2725 ;
         LAYER metal3 ;
         RECT  125.4675 31.1375 125.6025 31.2725 ;
         LAYER metal3 ;
         RECT  21.3175 37.1175 21.4525 37.2525 ;
         LAYER metal3 ;
         RECT  32.6425 72.265 112.3025 72.335 ;
         LAYER metal3 ;
         RECT  23.5175 2.4725 23.6525 2.6075 ;
         LAYER metal3 ;
         RECT  34.9575 2.4725 35.0925 2.6075 ;
         LAYER metal3 ;
         RECT  21.3175 40.1075 21.4525 40.2425 ;
         LAYER metal4 ;
         RECT  119.91 20.67 120.05 68.72 ;
         LAYER metal3 ;
         RECT  27.49 19.965 27.625 20.1 ;
         LAYER metal4 ;
         RECT  17.655 2.47 17.795 17.43 ;
         LAYER metal3 ;
         RECT  21.6625 25.1575 21.7975 25.2925 ;
         LAYER metal3 ;
         RECT  32.6425 79.1175 109.4825 79.1875 ;
         LAYER metal3 ;
         RECT  25.58 11.9075 25.715 12.0425 ;
         LAYER metal3 ;
         RECT  69.2775 2.4725 69.4125 2.6075 ;
         LAYER metal3 ;
         RECT  20.6575 2.4725 20.7925 2.6075 ;
         LAYER metal4 ;
         RECT  32.575 17.5 32.715 71.57 ;
         LAYER metal3 ;
         RECT  32.6425 8.415 109.4825 8.485 ;
         LAYER metal3 ;
         RECT  119.295 69.22 119.43 69.355 ;
         LAYER metal4 ;
         RECT  132.04 8.255 132.18 20.81 ;
         LAYER metal3 ;
         RECT  21.3175 34.1275 21.4525 34.2625 ;
         LAYER metal3 ;
         RECT  115.2875 70.0075 115.4225 70.1425 ;
         LAYER metal4 ;
         RECT  146.4275 54.42 146.5675 76.8225 ;
         LAYER metal3 ;
         RECT  31.4975 19.1775 31.6325 19.3125 ;
         LAYER metal3 ;
         RECT  80.7175 2.4725 80.8525 2.6075 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal3 ;
         RECT  21.6625 22.1675 21.7975 22.3025 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  121.205 74.6275 121.34 74.7625 ;
         LAYER metal4 ;
         RECT  119.35 20.6375 119.49 68.6825 ;
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal3 ;
         RECT  72.1375 0.0025 72.2725 0.1375 ;
         LAYER metal3 ;
         RECT  25.58 9.4375 25.715 9.5725 ;
         LAYER metal3 ;
         RECT  25.58 14.3775 25.715 14.5125 ;
         LAYER metal4 ;
         RECT  17.795 41.535 17.935 54.09 ;
         LAYER metal4 ;
         RECT  27.43 20.6375 27.57 68.6825 ;
         LAYER metal3 ;
         RECT  83.5775 0.0025 83.7125 0.1375 ;
         LAYER metal3 ;
         RECT  37.8175 0.0025 37.9525 0.1375 ;
         LAYER metal3 ;
         RECT  144.695 86.5325 144.83 86.6675 ;
         LAYER metal3 ;
         RECT  19.51 41.6025 19.645 41.7375 ;
         LAYER metal3 ;
         RECT  127.275 35.6225 127.41 35.7575 ;
         LAYER metal3 ;
         RECT  19.51 29.6425 19.645 29.7775 ;
         LAYER metal3 ;
         RECT  20.135 26.6525 20.27 26.7875 ;
         LAYER metal3 ;
         RECT  49.2575 0.0025 49.3925 0.1375 ;
         LAYER metal3 ;
         RECT  127.275 32.6325 127.41 32.7675 ;
         LAYER metal4 ;
         RECT  33.035 17.5 33.175 71.57 ;
         LAYER metal3 ;
         RECT  20.135 23.6625 20.27 23.7975 ;
         LAYER metal3 ;
         RECT  126.65 20.6725 126.785 20.8075 ;
         LAYER metal3 ;
         RECT  127.275 38.6125 127.41 38.7475 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal3 ;
         RECT  19.51 35.6225 19.645 35.7575 ;
         LAYER metal4 ;
         RECT  113.745 17.5 113.885 71.57 ;
         LAYER metal3 ;
         RECT  26.3775 0.0025 26.5125 0.1375 ;
         LAYER metal3 ;
         RECT  32.6425 74.885 111.16 74.955 ;
         LAYER metal3 ;
         RECT  19.51 38.6125 19.645 38.7475 ;
         LAYER metal4 ;
         RECT  129.18 8.32 129.32 20.875 ;
         LAYER metal3 ;
         RECT  32.6425 10.465 109.4825 10.535 ;
         LAYER metal4 ;
         RECT  25.28 20.6375 25.42 68.72 ;
         LAYER metal3 ;
         RECT  32.6425 14.185 111.16 14.255 ;
         LAYER metal3 ;
         RECT  19.51 32.6325 19.645 32.7675 ;
         LAYER metal3 ;
         RECT  95.0175 0.0025 95.1525 0.1375 ;
         LAYER metal4 ;
         RECT  140.87 71.71 141.01 86.67 ;
         LAYER metal3 ;
         RECT  106.4575 0.0025 106.5925 0.1375 ;
         LAYER metal3 ;
         RECT  120.6025 85.2675 120.7375 85.4025 ;
         LAYER metal3 ;
         RECT  126.65 26.6525 126.785 26.7875 ;
         LAYER metal3 ;
         RECT  126.65 23.6625 126.785 23.7975 ;
         LAYER metal4 ;
         RECT  144.365 54.3875 144.505 76.79 ;
         LAYER metal3 ;
         RECT  23.5175 0.0025 23.6525 0.1375 ;
         LAYER metal3 ;
         RECT  60.6975 0.0025 60.8325 0.1375 ;
         LAYER metal3 ;
         RECT  127.275 41.6025 127.41 41.7375 ;
         LAYER metal3 ;
         RECT  20.135 20.6725 20.27 20.8075 ;
         LAYER metal3 ;
         RECT  127.275 29.6425 127.41 29.7775 ;
         LAYER metal3 ;
         RECT  32.6425 77.225 109.5175 77.295 ;
         LAYER metal3 ;
         RECT  121.205 79.5675 121.34 79.7025 ;
         LAYER metal4 ;
         RECT  121.5 20.6375 121.64 68.72 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 147.115 86.53 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 147.115 86.53 ;
   LAYER  metal3 ;
      RECT  24.075 0.9675 26.52 1.3825 ;
      RECT  26.935 0.9675 29.38 1.3825 ;
      RECT  29.795 0.9675 32.24 1.3825 ;
      RECT  32.655 0.9675 35.1 1.3825 ;
      RECT  35.515 0.9675 37.96 1.3825 ;
      RECT  38.375 0.9675 40.82 1.3825 ;
      RECT  41.235 0.9675 43.68 1.3825 ;
      RECT  44.095 0.9675 46.54 1.3825 ;
      RECT  46.955 0.9675 49.4 1.3825 ;
      RECT  49.815 0.9675 52.26 1.3825 ;
      RECT  52.675 0.9675 55.12 1.3825 ;
      RECT  55.535 0.9675 57.98 1.3825 ;
      RECT  58.395 0.9675 60.84 1.3825 ;
      RECT  61.255 0.9675 63.7 1.3825 ;
      RECT  64.115 0.9675 66.56 1.3825 ;
      RECT  66.975 0.9675 69.42 1.3825 ;
      RECT  69.835 0.9675 72.28 1.3825 ;
      RECT  72.695 0.9675 75.14 1.3825 ;
      RECT  75.555 0.9675 78.0 1.3825 ;
      RECT  78.415 0.9675 80.86 1.3825 ;
      RECT  81.275 0.9675 83.72 1.3825 ;
      RECT  84.135 0.9675 86.58 1.3825 ;
      RECT  86.995 0.9675 89.44 1.3825 ;
      RECT  89.855 0.9675 92.3 1.3825 ;
      RECT  92.715 0.9675 95.16 1.3825 ;
      RECT  95.575 0.9675 98.02 1.3825 ;
      RECT  98.435 0.9675 100.88 1.3825 ;
      RECT  101.295 0.9675 103.74 1.3825 ;
      RECT  104.155 0.9675 106.6 1.3825 ;
      RECT  107.015 0.9675 109.46 1.3825 ;
      RECT  109.875 0.9675 112.32 1.3825 ;
      RECT  112.735 0.9675 147.115 1.3825 ;
      RECT  21.215 0.9675 23.66 1.3825 ;
      RECT  0.14 42.5675 15.08 42.9825 ;
      RECT  0.14 42.9825 15.08 86.53 ;
      RECT  15.08 1.3825 15.495 42.5675 ;
      RECT  15.495 42.5675 23.66 42.9825 ;
      RECT  15.495 42.9825 23.66 86.53 ;
      RECT  15.08 42.9825 15.495 45.2975 ;
      RECT  15.08 45.7125 15.495 47.5075 ;
      RECT  15.08 47.9225 15.495 50.2375 ;
      RECT  15.08 50.6525 15.495 52.4475 ;
      RECT  15.08 52.8625 15.495 86.53 ;
      RECT  24.075 84.0225 123.04 84.4375 ;
      RECT  123.04 84.4375 123.455 86.53 ;
      RECT  123.455 1.3825 131.62 19.4275 ;
      RECT  123.455 19.4275 131.62 19.8425 ;
      RECT  131.62 19.8425 132.035 84.0225 ;
      RECT  132.035 1.3825 147.115 19.4275 ;
      RECT  132.035 19.4275 147.115 19.8425 ;
      RECT  131.62 17.1125 132.035 19.4275 ;
      RECT  131.62 14.9025 132.035 16.6975 ;
      RECT  131.62 12.1725 132.035 14.4875 ;
      RECT  131.62 1.3825 132.035 9.5475 ;
      RECT  131.62 9.9625 132.035 11.7575 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  146.695 84.4375 147.11 85.2875 ;
      RECT  146.695 85.7025 147.11 86.53 ;
      RECT  147.11 84.4375 147.115 85.2875 ;
      RECT  147.11 85.2875 147.115 85.7025 ;
      RECT  147.11 85.7025 147.115 86.53 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 42.5675 ;
      RECT  6.5225 1.3825 15.08 1.4675 ;
      RECT  6.5225 1.4675 15.08 42.5675 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 20.8 1.0525 ;
      RECT  6.5225 1.0525 20.8 1.3825 ;
      RECT  123.455 84.4375 140.5925 85.2025 ;
      RECT  123.455 85.2025 140.5925 85.2875 ;
      RECT  140.5925 84.4375 141.0075 85.2025 ;
      RECT  141.0075 84.4375 146.695 85.2025 ;
      RECT  141.0075 85.2025 146.695 85.2875 ;
      RECT  123.455 85.2875 140.5925 85.6175 ;
      RECT  123.455 85.6175 140.5925 85.7025 ;
      RECT  140.5925 85.6175 141.0075 85.7025 ;
      RECT  141.0075 85.2875 146.695 85.6175 ;
      RECT  141.0075 85.6175 146.695 85.7025 ;
      RECT  24.075 81.535 35.6875 81.95 ;
      RECT  24.075 81.95 35.6875 84.0225 ;
      RECT  35.6875 81.95 36.1025 84.0225 ;
      RECT  36.1025 81.95 123.04 84.0225 ;
      RECT  36.1025 81.535 38.0375 81.95 ;
      RECT  38.4525 81.535 40.3875 81.95 ;
      RECT  40.8025 81.535 42.7375 81.95 ;
      RECT  43.1525 81.535 45.0875 81.95 ;
      RECT  45.5025 81.535 47.4375 81.95 ;
      RECT  47.8525 81.535 49.7875 81.95 ;
      RECT  50.2025 81.535 52.1375 81.95 ;
      RECT  52.5525 81.535 54.4875 81.95 ;
      RECT  54.9025 81.535 56.8375 81.95 ;
      RECT  57.2525 81.535 59.1875 81.95 ;
      RECT  59.6025 81.535 61.5375 81.95 ;
      RECT  61.9525 81.535 63.8875 81.95 ;
      RECT  64.3025 81.535 66.2375 81.95 ;
      RECT  66.6525 81.535 68.5875 81.95 ;
      RECT  69.0025 81.535 70.9375 81.95 ;
      RECT  71.3525 81.535 73.2875 81.95 ;
      RECT  73.7025 81.535 75.6375 81.95 ;
      RECT  76.0525 81.535 77.9875 81.95 ;
      RECT  78.4025 81.535 80.3375 81.95 ;
      RECT  80.7525 81.535 82.6875 81.95 ;
      RECT  83.1025 81.535 85.0375 81.95 ;
      RECT  85.4525 81.535 87.3875 81.95 ;
      RECT  87.8025 81.535 89.7375 81.95 ;
      RECT  90.1525 81.535 92.0875 81.95 ;
      RECT  92.5025 81.535 94.4375 81.95 ;
      RECT  94.8525 81.535 96.7875 81.95 ;
      RECT  97.2025 81.535 99.1375 81.95 ;
      RECT  99.5525 81.535 101.4875 81.95 ;
      RECT  101.9025 81.535 103.8375 81.95 ;
      RECT  104.2525 81.535 106.1875 81.95 ;
      RECT  106.6025 81.535 108.5375 81.95 ;
      RECT  108.9525 81.535 123.04 81.95 ;
      RECT  24.075 16.665 32.5025 17.015 ;
      RECT  111.2675 16.665 123.04 17.015 ;
      RECT  123.455 19.8425 124.9825 25.0175 ;
      RECT  123.455 25.0175 124.9825 25.4325 ;
      RECT  125.3975 25.0175 131.62 25.4325 ;
      RECT  111.2675 76.9575 121.065 77.3725 ;
      RECT  111.2675 77.3725 121.065 81.535 ;
      RECT  121.48 17.015 123.04 76.9575 ;
      RECT  121.48 76.9575 123.04 77.3725 ;
      RECT  121.48 77.3725 123.04 81.535 ;
      RECT  124.9825 25.4325 125.3275 33.9875 ;
      RECT  124.9825 33.9875 125.3275 34.4025 ;
      RECT  124.9825 34.4025 125.3275 84.0225 ;
      RECT  125.7425 33.9875 131.62 34.4025 ;
      RECT  36.1025 1.3825 92.0175 2.3325 ;
      RECT  92.0175 1.3825 92.4325 2.3325 ;
      RECT  92.4325 1.3825 111.2675 2.3325 ;
      RECT  92.4325 2.3325 103.4575 2.7475 ;
      RECT  103.8725 2.3325 111.2675 2.7475 ;
      RECT  124.9825 19.8425 125.3975 22.0275 ;
      RECT  124.9825 22.4425 125.3975 25.0175 ;
      RECT  123.455 84.0225 144.555 84.3375 ;
      RECT  123.455 84.3375 144.555 84.4375 ;
      RECT  144.555 84.3375 144.97 84.4375 ;
      RECT  144.97 84.0225 147.115 84.3375 ;
      RECT  144.97 84.3375 147.115 84.4375 ;
      RECT  132.035 19.8425 144.555 83.9225 ;
      RECT  132.035 83.9225 144.555 84.0225 ;
      RECT  144.555 19.8425 144.97 83.9225 ;
      RECT  144.97 19.8425 147.115 83.9225 ;
      RECT  144.97 83.9225 147.115 84.0225 ;
      RECT  36.1025 2.3325 46.2575 2.7475 ;
      RECT  125.3275 40.3825 125.3975 84.0225 ;
      RECT  125.3975 40.3825 125.7425 84.0225 ;
      RECT  123.04 1.3825 123.3225 82.6575 ;
      RECT  123.04 82.6575 123.3225 83.0725 ;
      RECT  123.04 83.0725 123.3225 84.0225 ;
      RECT  123.3225 1.3825 123.455 82.6575 ;
      RECT  123.3225 83.0725 123.455 84.0225 ;
      RECT  123.455 25.4325 123.7375 82.6575 ;
      RECT  123.455 83.0725 123.7375 84.0225 ;
      RECT  123.7375 25.4325 124.9825 82.6575 ;
      RECT  123.7375 82.6575 124.9825 83.0725 ;
      RECT  123.7375 83.0725 124.9825 84.0225 ;
      RECT  125.3275 34.4025 125.3975 36.9775 ;
      RECT  125.3275 37.3925 125.3975 39.9675 ;
      RECT  125.3975 34.4025 125.7425 36.9775 ;
      RECT  125.3975 37.3925 125.7425 39.9675 ;
      RECT  46.6725 2.3325 57.6975 2.7475 ;
      RECT  15.495 30.9975 21.1775 31.4125 ;
      RECT  21.5925 30.9975 23.66 31.4125 ;
      RECT  21.5925 31.4125 23.66 42.5675 ;
      RECT  125.3275 25.4325 125.3975 30.9975 ;
      RECT  125.3275 31.4125 125.3975 33.9875 ;
      RECT  125.3975 25.4325 125.7425 30.9975 ;
      RECT  125.3975 31.4125 125.7425 33.9875 ;
      RECT  32.5025 17.015 35.6875 72.125 ;
      RECT  35.6875 17.015 36.1025 72.125 ;
      RECT  36.1025 17.015 111.2675 72.125 ;
      RECT  111.2675 17.015 112.4425 72.125 ;
      RECT  112.4425 72.125 121.065 72.475 ;
      RECT  112.4425 72.475 121.065 76.9575 ;
      RECT  23.66 1.3825 23.7925 2.3325 ;
      RECT  23.66 2.7475 23.7925 86.53 ;
      RECT  23.7925 1.3825 24.075 2.3325 ;
      RECT  23.7925 2.3325 24.075 2.7475 ;
      RECT  23.7925 2.7475 24.075 86.53 ;
      RECT  21.5925 1.3825 23.3775 2.3325 ;
      RECT  21.5925 2.3325 23.3775 2.7475 ;
      RECT  23.3775 1.3825 23.66 2.3325 ;
      RECT  23.3775 2.7475 23.66 30.9975 ;
      RECT  32.5025 1.3825 34.8175 2.3325 ;
      RECT  32.5025 2.3325 34.8175 2.7475 ;
      RECT  34.8175 1.3825 35.2325 2.3325 ;
      RECT  35.2325 1.3825 35.6875 2.3325 ;
      RECT  35.2325 2.3325 35.6875 2.7475 ;
      RECT  21.1775 37.3925 21.5925 39.9675 ;
      RECT  21.1775 40.3825 21.5925 42.5675 ;
      RECT  24.075 17.015 27.35 19.825 ;
      RECT  24.075 19.825 27.35 20.24 ;
      RECT  24.075 20.24 27.35 81.535 ;
      RECT  27.35 17.015 27.765 19.825 ;
      RECT  27.35 20.24 27.765 81.535 ;
      RECT  27.765 19.825 32.5025 20.24 ;
      RECT  27.765 20.24 32.5025 81.535 ;
      RECT  21.1775 1.3825 21.5225 25.0175 ;
      RECT  21.1775 25.0175 21.5225 25.4325 ;
      RECT  21.1775 25.4325 21.5225 30.9975 ;
      RECT  21.5225 25.4325 21.5925 30.9975 ;
      RECT  21.5925 25.4325 21.9375 30.9975 ;
      RECT  21.9375 2.7475 23.3775 25.0175 ;
      RECT  21.9375 25.0175 23.3775 25.4325 ;
      RECT  21.9375 25.4325 23.3775 30.9975 ;
      RECT  32.5025 79.3275 35.6875 81.535 ;
      RECT  35.6875 79.3275 36.1025 81.535 ;
      RECT  36.1025 79.3275 109.6225 81.535 ;
      RECT  109.6225 78.9775 111.2675 79.3275 ;
      RECT  109.6225 79.3275 111.2675 81.535 ;
      RECT  24.075 1.3825 25.44 11.7675 ;
      RECT  24.075 11.7675 25.44 12.1825 ;
      RECT  24.075 12.1825 25.44 16.665 ;
      RECT  25.855 1.3825 32.5025 11.7675 ;
      RECT  25.855 11.7675 32.5025 12.1825 ;
      RECT  25.855 12.1825 32.5025 16.665 ;
      RECT  58.1125 2.3325 69.1375 2.7475 ;
      RECT  15.495 1.3825 20.5175 2.3325 ;
      RECT  15.495 2.3325 20.5175 2.7475 ;
      RECT  20.5175 1.3825 20.9325 2.3325 ;
      RECT  20.5175 2.7475 20.9325 30.9975 ;
      RECT  20.9325 1.3825 21.1775 2.3325 ;
      RECT  20.9325 2.3325 21.1775 2.7475 ;
      RECT  20.9325 2.7475 21.1775 30.9975 ;
      RECT  35.6875 1.3825 36.1025 8.275 ;
      RECT  36.1025 2.7475 92.0175 8.275 ;
      RECT  92.0175 2.7475 92.4325 8.275 ;
      RECT  92.4325 2.7475 109.6225 8.275 ;
      RECT  109.6225 2.7475 111.2675 8.275 ;
      RECT  109.6225 8.275 111.2675 8.625 ;
      RECT  32.5025 2.7475 34.8175 8.275 ;
      RECT  34.8175 2.7475 35.2325 8.275 ;
      RECT  35.2325 2.7475 35.6875 8.275 ;
      RECT  112.4425 17.015 119.155 69.08 ;
      RECT  112.4425 69.08 119.155 69.495 ;
      RECT  119.155 17.015 119.57 69.08 ;
      RECT  119.155 69.495 119.57 72.125 ;
      RECT  119.57 17.015 121.065 69.08 ;
      RECT  119.57 69.08 121.065 69.495 ;
      RECT  119.57 69.495 121.065 72.125 ;
      RECT  21.1775 31.4125 21.5925 33.9875 ;
      RECT  21.1775 34.4025 21.5925 36.9775 ;
      RECT  112.4425 69.495 115.1475 69.8675 ;
      RECT  112.4425 69.8675 115.1475 70.2825 ;
      RECT  112.4425 70.2825 115.1475 72.125 ;
      RECT  115.1475 69.495 115.5625 69.8675 ;
      RECT  115.1475 70.2825 115.5625 72.125 ;
      RECT  115.5625 69.495 119.155 69.8675 ;
      RECT  115.5625 69.8675 119.155 70.2825 ;
      RECT  115.5625 70.2825 119.155 72.125 ;
      RECT  27.765 17.015 31.3575 19.0375 ;
      RECT  27.765 19.0375 31.3575 19.4525 ;
      RECT  27.765 19.4525 31.3575 19.825 ;
      RECT  31.3575 17.015 31.7725 19.0375 ;
      RECT  31.3575 19.4525 31.7725 19.825 ;
      RECT  31.7725 17.015 32.5025 19.0375 ;
      RECT  31.7725 19.0375 32.5025 19.4525 ;
      RECT  31.7725 19.4525 32.5025 19.825 ;
      RECT  69.5525 2.3325 80.5775 2.7475 ;
      RECT  80.9925 2.3325 92.0175 2.7475 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 42.5675 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 42.5675 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 42.5675 ;
      RECT  21.5225 1.3825 21.5925 22.0275 ;
      RECT  21.5225 22.4425 21.5925 25.0175 ;
      RECT  21.5925 2.7475 21.9375 22.0275 ;
      RECT  21.5925 22.4425 21.9375 25.0175 ;
      RECT  121.065 17.015 121.48 74.4875 ;
      RECT  121.065 74.9025 121.48 76.9575 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  0.14 0.2775 2.285 0.9675 ;
      RECT  2.285 0.2775 2.7 0.9675 ;
      RECT  2.7 0.2775 23.66 0.9675 ;
      RECT  24.075 0.2775 71.9975 0.9675 ;
      RECT  71.9975 0.2775 72.4125 0.9675 ;
      RECT  72.4125 0.2775 147.115 0.9675 ;
      RECT  25.44 1.3825 25.855 9.2975 ;
      RECT  25.44 9.7125 25.855 11.7675 ;
      RECT  25.44 12.1825 25.855 14.2375 ;
      RECT  25.44 14.6525 25.855 16.665 ;
      RECT  72.4125 0.14 83.4375 0.2775 ;
      RECT  123.455 85.7025 144.555 86.3925 ;
      RECT  123.455 86.3925 144.555 86.53 ;
      RECT  144.555 85.7025 144.97 86.3925 ;
      RECT  144.97 85.7025 146.695 86.3925 ;
      RECT  144.97 86.3925 146.695 86.53 ;
      RECT  15.495 31.4125 19.37 41.4625 ;
      RECT  15.495 41.4625 19.37 41.8775 ;
      RECT  15.495 41.8775 19.37 42.5675 ;
      RECT  19.37 41.8775 19.785 42.5675 ;
      RECT  19.785 31.4125 21.1775 41.4625 ;
      RECT  19.785 41.4625 21.1775 41.8775 ;
      RECT  19.785 41.8775 21.1775 42.5675 ;
      RECT  125.7425 34.4025 127.135 35.4825 ;
      RECT  125.7425 35.4825 127.135 35.8975 ;
      RECT  125.7425 35.8975 127.135 84.0225 ;
      RECT  127.135 34.4025 127.55 35.4825 ;
      RECT  127.55 34.4025 131.62 35.4825 ;
      RECT  127.55 35.4825 131.62 35.8975 ;
      RECT  127.55 35.8975 131.62 84.0225 ;
      RECT  15.495 2.7475 19.37 29.5025 ;
      RECT  15.495 29.5025 19.37 29.9175 ;
      RECT  15.495 29.9175 19.37 30.9975 ;
      RECT  19.37 2.7475 19.785 29.5025 ;
      RECT  19.37 29.9175 19.785 30.9975 ;
      RECT  19.785 29.5025 20.5175 29.9175 ;
      RECT  19.785 29.9175 20.5175 30.9975 ;
      RECT  19.785 2.7475 19.995 26.5125 ;
      RECT  19.785 26.5125 19.995 26.9275 ;
      RECT  19.785 26.9275 19.995 29.5025 ;
      RECT  19.995 26.9275 20.41 29.5025 ;
      RECT  20.41 2.7475 20.5175 26.5125 ;
      RECT  20.41 26.5125 20.5175 26.9275 ;
      RECT  20.41 26.9275 20.5175 29.5025 ;
      RECT  38.0925 0.14 49.1175 0.2775 ;
      RECT  125.7425 32.4925 127.135 32.9075 ;
      RECT  125.7425 32.9075 127.135 33.9875 ;
      RECT  127.135 32.9075 127.55 33.9875 ;
      RECT  127.55 25.4325 131.62 32.4925 ;
      RECT  127.55 32.4925 131.62 32.9075 ;
      RECT  127.55 32.9075 131.62 33.9875 ;
      RECT  19.995 23.9375 20.41 26.5125 ;
      RECT  125.3975 19.8425 126.51 20.5325 ;
      RECT  125.3975 20.5325 126.51 20.9475 ;
      RECT  125.3975 20.9475 126.51 25.0175 ;
      RECT  126.51 19.8425 126.925 20.5325 ;
      RECT  126.925 19.8425 131.62 20.5325 ;
      RECT  126.925 20.5325 131.62 20.9475 ;
      RECT  126.925 20.9475 131.62 25.0175 ;
      RECT  127.135 35.8975 127.55 38.4725 ;
      RECT  24.075 0.14 26.2375 0.2775 ;
      RECT  26.6525 0.14 37.6775 0.2775 ;
      RECT  111.2675 72.475 111.3 74.745 ;
      RECT  111.2675 75.095 111.3 76.9575 ;
      RECT  111.3 72.475 112.4425 74.745 ;
      RECT  111.3 74.745 112.4425 75.095 ;
      RECT  111.3 75.095 112.4425 76.9575 ;
      RECT  32.5025 72.475 35.6875 74.745 ;
      RECT  35.6875 72.475 36.1025 74.745 ;
      RECT  36.1025 72.475 109.6225 74.745 ;
      RECT  109.6225 72.475 111.2675 74.745 ;
      RECT  19.37 35.8975 19.785 38.4725 ;
      RECT  19.37 38.8875 19.785 41.4625 ;
      RECT  35.6875 8.625 36.1025 10.325 ;
      RECT  36.1025 8.625 92.0175 10.325 ;
      RECT  92.0175 8.625 92.4325 10.325 ;
      RECT  92.4325 8.625 109.6225 10.325 ;
      RECT  32.5025 8.625 34.8175 10.325 ;
      RECT  34.8175 8.625 35.2325 10.325 ;
      RECT  35.2325 8.625 35.6875 10.325 ;
      RECT  111.2675 1.3825 111.3 14.045 ;
      RECT  111.2675 14.395 111.3 16.665 ;
      RECT  111.3 1.3825 123.04 14.045 ;
      RECT  111.3 14.045 123.04 14.395 ;
      RECT  111.3 14.395 123.04 16.665 ;
      RECT  109.6225 8.625 111.2675 14.045 ;
      RECT  109.6225 14.395 111.2675 16.665 ;
      RECT  35.6875 10.675 36.1025 14.045 ;
      RECT  35.6875 14.395 36.1025 16.665 ;
      RECT  36.1025 10.675 92.0175 14.045 ;
      RECT  36.1025 14.395 92.0175 16.665 ;
      RECT  92.0175 10.675 92.4325 14.045 ;
      RECT  92.0175 14.395 92.4325 16.665 ;
      RECT  92.4325 10.675 109.6225 14.045 ;
      RECT  92.4325 14.395 109.6225 16.665 ;
      RECT  32.5025 10.675 34.8175 14.045 ;
      RECT  32.5025 14.395 34.8175 16.665 ;
      RECT  34.8175 10.675 35.2325 14.045 ;
      RECT  34.8175 14.395 35.2325 16.665 ;
      RECT  35.2325 10.675 35.6875 14.045 ;
      RECT  35.2325 14.395 35.6875 16.665 ;
      RECT  19.37 31.4125 19.785 32.4925 ;
      RECT  19.37 32.9075 19.785 35.4825 ;
      RECT  83.8525 0.14 94.8775 0.2775 ;
      RECT  95.2925 0.14 106.3175 0.2775 ;
      RECT  106.7325 0.14 147.115 0.2775 ;
      RECT  24.075 84.4375 120.4625 85.1275 ;
      RECT  24.075 85.1275 120.4625 85.5425 ;
      RECT  24.075 85.5425 120.4625 86.53 ;
      RECT  120.4625 84.4375 120.8775 85.1275 ;
      RECT  120.4625 85.5425 120.8775 86.53 ;
      RECT  120.8775 84.4375 123.04 85.1275 ;
      RECT  120.8775 85.1275 123.04 85.5425 ;
      RECT  120.8775 85.5425 123.04 86.53 ;
      RECT  125.7425 25.4325 126.51 26.5125 ;
      RECT  125.7425 26.5125 126.51 26.9275 ;
      RECT  125.7425 26.9275 126.51 32.4925 ;
      RECT  126.51 25.4325 126.925 26.5125 ;
      RECT  126.51 26.9275 126.925 32.4925 ;
      RECT  126.925 25.4325 127.135 26.5125 ;
      RECT  126.925 26.5125 127.135 26.9275 ;
      RECT  126.925 26.9275 127.135 32.4925 ;
      RECT  126.51 20.9475 126.925 23.5225 ;
      RECT  126.51 23.9375 126.925 25.0175 ;
      RECT  23.66 0.2775 23.7925 0.9675 ;
      RECT  23.7925 0.14 24.075 0.2775 ;
      RECT  23.7925 0.2775 24.075 0.9675 ;
      RECT  2.7 0.14 23.3775 0.2775 ;
      RECT  49.5325 0.14 60.5575 0.2775 ;
      RECT  60.9725 0.14 71.9975 0.2775 ;
      RECT  127.135 38.8875 127.55 41.4625 ;
      RECT  127.135 41.8775 127.55 84.0225 ;
      RECT  19.995 2.7475 20.41 20.5325 ;
      RECT  19.995 20.9475 20.41 23.5225 ;
      RECT  127.135 25.4325 127.55 29.5025 ;
      RECT  127.135 29.9175 127.55 32.4925 ;
      RECT  32.5025 75.095 35.6875 77.085 ;
      RECT  32.5025 77.435 35.6875 78.9775 ;
      RECT  35.6875 75.095 36.1025 77.085 ;
      RECT  35.6875 77.435 36.1025 78.9775 ;
      RECT  36.1025 75.095 109.6225 77.085 ;
      RECT  36.1025 77.435 109.6225 78.9775 ;
      RECT  109.6225 75.095 109.6575 77.085 ;
      RECT  109.6225 77.435 109.6575 78.9775 ;
      RECT  109.6575 75.095 111.2675 77.085 ;
      RECT  109.6575 77.085 111.2675 77.435 ;
      RECT  109.6575 77.435 111.2675 78.9775 ;
      RECT  121.065 77.3725 121.48 79.4275 ;
      RECT  121.065 79.8425 121.48 81.535 ;
   LAYER  metal4 ;
      RECT  31.215 0.14 31.915 20.39 ;
      RECT  31.215 68.93 31.915 86.53 ;
      RECT  0.14 69.0 26.59 86.53 ;
      RECT  26.59 69.0 27.29 86.53 ;
      RECT  27.29 69.0 31.215 86.53 ;
      RECT  31.915 73.9 129.04 84.48 ;
      RECT  31.915 84.48 129.04 86.53 ;
      RECT  129.04 68.93 129.74 73.9 ;
      RECT  129.04 84.48 129.74 86.53 ;
      RECT  0.14 41.32 14.655 54.435 ;
      RECT  0.14 54.435 14.655 68.93 ;
      RECT  14.655 20.39 15.355 41.32 ;
      RECT  14.655 54.435 15.355 68.93 ;
      RECT  31.915 0.14 113.925 17.22 ;
      RECT  113.925 0.14 114.625 17.22 ;
      RECT  31.915 71.85 113.925 73.9 ;
      RECT  113.925 71.85 114.625 73.9 ;
      RECT  114.625 71.85 129.04 73.9 ;
      RECT  114.625 20.39 115.005 68.93 ;
      RECT  0.14 0.14 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 20.39 ;
      RECT  0.4075 0.14 1.1075 9.5675 ;
      RECT  0.14 20.39 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 41.32 ;
      RECT  0.4075 32.53 1.1075 41.32 ;
      RECT  114.625 69.0 119.63 71.85 ;
      RECT  119.63 69.0 120.33 71.85 ;
      RECT  120.33 69.0 129.04 71.85 ;
      RECT  17.375 0.14 18.075 2.19 ;
      RECT  18.075 0.14 31.215 2.19 ;
      RECT  18.075 2.19 31.215 9.5675 ;
      RECT  17.375 17.71 18.075 20.39 ;
      RECT  18.075 9.5675 31.215 17.71 ;
      RECT  31.915 17.22 32.295 20.39 ;
      RECT  31.915 20.39 32.295 68.93 ;
      RECT  31.915 68.93 32.295 71.85 ;
      RECT  114.625 0.14 131.76 7.975 ;
      RECT  131.76 0.14 132.46 7.975 ;
      RECT  132.46 0.14 147.115 7.975 ;
      RECT  132.46 7.975 147.115 17.22 ;
      RECT  132.46 17.22 147.115 20.39 ;
      RECT  131.76 21.09 132.46 68.93 ;
      RECT  132.46 20.39 147.115 21.09 ;
      RECT  146.8475 68.93 147.115 73.9 ;
      RECT  146.1475 77.1025 146.8475 84.48 ;
      RECT  146.8475 73.9 147.115 77.1025 ;
      RECT  146.8475 77.1025 147.115 84.48 ;
      RECT  146.1475 21.09 146.8475 54.14 ;
      RECT  146.8475 21.09 147.115 54.14 ;
      RECT  146.8475 54.14 147.115 68.93 ;
      RECT  114.625 68.93 119.07 68.9625 ;
      RECT  114.625 68.9625 119.07 69.0 ;
      RECT  119.07 68.9625 119.63 69.0 ;
      RECT  115.705 20.39 119.07 68.93 ;
      RECT  114.625 17.22 119.07 20.3575 ;
      RECT  114.625 20.3575 119.07 20.39 ;
      RECT  119.07 17.22 119.77 20.3575 ;
      RECT  1.1075 0.14 5.825 2.19 ;
      RECT  6.525 0.14 17.375 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 17.375 9.5675 ;
      RECT  5.825 15.24 6.525 17.71 ;
      RECT  6.525 9.5675 17.375 15.24 ;
      RECT  6.525 15.24 17.375 17.71 ;
      RECT  15.355 20.39 17.515 41.255 ;
      RECT  15.355 41.255 17.515 41.32 ;
      RECT  17.515 20.39 18.215 41.255 ;
      RECT  15.355 41.32 17.515 54.37 ;
      RECT  15.355 54.37 17.515 54.435 ;
      RECT  17.515 54.37 18.215 54.435 ;
      RECT  27.85 20.39 31.215 68.93 ;
      RECT  27.29 68.9625 27.85 69.0 ;
      RECT  27.85 68.93 31.215 68.9625 ;
      RECT  27.85 68.9625 31.215 69.0 ;
      RECT  18.075 17.71 27.15 20.3575 ;
      RECT  27.15 17.71 27.85 20.3575 ;
      RECT  27.85 17.71 31.215 20.3575 ;
      RECT  27.85 20.3575 31.215 20.39 ;
      RECT  1.1075 20.39 2.47 32.53 ;
      RECT  3.17 20.39 14.655 32.53 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 41.32 ;
      RECT  2.47 32.5625 3.17 41.32 ;
      RECT  3.17 32.53 14.655 32.5625 ;
      RECT  3.17 32.5625 14.655 41.32 ;
      RECT  1.1075 17.71 2.47 20.39 ;
      RECT  3.17 17.71 17.375 20.39 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 15.24 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  1.1075 15.24 2.47 17.71 ;
      RECT  3.17 15.24 5.825 17.71 ;
      RECT  33.455 17.22 113.465 20.39 ;
      RECT  33.455 20.39 113.465 68.93 ;
      RECT  33.455 68.93 113.465 71.85 ;
      RECT  114.625 7.975 128.9 8.04 ;
      RECT  114.625 8.04 128.9 17.22 ;
      RECT  128.9 7.975 129.6 8.04 ;
      RECT  129.6 7.975 131.76 8.04 ;
      RECT  129.6 8.04 131.76 17.22 ;
      RECT  129.6 20.39 131.76 21.09 ;
      RECT  128.9 21.155 129.6 68.93 ;
      RECT  129.6 21.09 131.76 21.155 ;
      RECT  129.6 21.155 131.76 68.93 ;
      RECT  119.77 17.22 128.9 20.3575 ;
      RECT  129.6 17.22 131.76 20.3575 ;
      RECT  129.6 20.3575 131.76 20.39 ;
      RECT  0.14 68.93 25.0 69.0 ;
      RECT  25.7 68.93 26.59 69.0 ;
      RECT  15.355 54.435 25.0 68.93 ;
      RECT  25.7 54.435 26.59 68.93 ;
      RECT  18.215 20.39 25.0 41.255 ;
      RECT  25.7 20.39 26.59 41.255 ;
      RECT  18.215 41.255 25.0 41.32 ;
      RECT  25.7 41.255 26.59 41.32 ;
      RECT  18.215 41.32 25.0 54.37 ;
      RECT  25.7 41.32 26.59 54.37 ;
      RECT  18.215 54.37 25.0 54.435 ;
      RECT  25.7 54.37 26.59 54.435 ;
      RECT  18.075 20.3575 25.0 20.39 ;
      RECT  25.7 20.3575 27.15 20.39 ;
      RECT  129.74 84.48 140.59 86.53 ;
      RECT  141.29 84.48 147.115 86.53 ;
      RECT  129.74 68.93 140.59 71.43 ;
      RECT  129.74 71.43 140.59 73.9 ;
      RECT  140.59 68.93 141.29 71.43 ;
      RECT  129.74 73.9 140.59 77.1025 ;
      RECT  129.74 77.1025 140.59 84.48 ;
      RECT  141.29 77.1025 146.1475 84.48 ;
      RECT  132.46 21.09 144.085 54.1075 ;
      RECT  132.46 54.1075 144.085 54.14 ;
      RECT  144.085 21.09 144.785 54.1075 ;
      RECT  144.785 21.09 146.1475 54.1075 ;
      RECT  144.785 54.1075 146.1475 54.14 ;
      RECT  132.46 54.14 144.085 68.93 ;
      RECT  144.785 54.14 146.1475 68.93 ;
      RECT  141.29 68.93 144.085 71.43 ;
      RECT  144.785 68.93 146.1475 71.43 ;
      RECT  141.29 71.43 144.085 73.9 ;
      RECT  144.785 71.43 146.1475 73.9 ;
      RECT  141.29 73.9 144.085 77.07 ;
      RECT  141.29 77.07 144.085 77.1025 ;
      RECT  144.085 77.07 144.785 77.1025 ;
      RECT  144.785 73.9 146.1475 77.07 ;
      RECT  144.785 77.07 146.1475 77.1025 ;
      RECT  120.33 68.93 121.22 69.0 ;
      RECT  121.92 68.93 129.04 69.0 ;
      RECT  120.33 20.39 121.22 21.09 ;
      RECT  121.92 20.39 128.9 21.09 ;
      RECT  120.33 21.09 121.22 21.155 ;
      RECT  121.92 21.09 128.9 21.155 ;
      RECT  120.33 21.155 121.22 68.93 ;
      RECT  121.92 21.155 128.9 68.93 ;
      RECT  119.77 20.3575 121.22 20.39 ;
      RECT  121.92 20.3575 128.9 20.39 ;
   END
END    freepdk45_sram_1w1r_64x32_32
END    LIBRARY
