../macros/freepdk45_sram_1w1r_96x32_32/freepdk45_sram_1w1r_96x32_32.lef