../macros/freepdk45_sram_1w1r_512x64_64/freepdk45_sram_1w1r_512x64_64.lef