VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1rw0r_45x512
   CLASS BLOCK ;
   SIZE 1593.62 BY 218.82 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.345 4.2375 126.48 4.3725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.205 4.2375 129.34 4.3725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.065 4.2375 132.2 4.3725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.925 4.2375 135.06 4.3725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.785 4.2375 137.92 4.3725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.645 4.2375 140.78 4.3725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.505 4.2375 143.64 4.3725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.365 4.2375 146.5 4.3725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.225 4.2375 149.36 4.3725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.085 4.2375 152.22 4.3725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.945 4.2375 155.08 4.3725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.805 4.2375 157.94 4.3725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.665 4.2375 160.8 4.3725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.525 4.2375 163.66 4.3725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.385 4.2375 166.52 4.3725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.245 4.2375 169.38 4.3725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.105 4.2375 172.24 4.3725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.965 4.2375 175.1 4.3725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.825 4.2375 177.96 4.3725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.685 4.2375 180.82 4.3725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.545 4.2375 183.68 4.3725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.405 4.2375 186.54 4.3725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.265 4.2375 189.4 4.3725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.125 4.2375 192.26 4.3725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.985 4.2375 195.12 4.3725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.845 4.2375 197.98 4.3725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.705 4.2375 200.84 4.3725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.565 4.2375 203.7 4.3725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.425 4.2375 206.56 4.3725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.285 4.2375 209.42 4.3725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.145 4.2375 212.28 4.3725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.005 4.2375 215.14 4.3725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.865 4.2375 218.0 4.3725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.725 4.2375 220.86 4.3725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.585 4.2375 223.72 4.3725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.445 4.2375 226.58 4.3725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.305 4.2375 229.44 4.3725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.165 4.2375 232.3 4.3725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.025 4.2375 235.16 4.3725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.885 4.2375 238.02 4.3725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.745 4.2375 240.88 4.3725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.605 4.2375 243.74 4.3725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.465 4.2375 246.6 4.3725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.325 4.2375 249.46 4.3725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.185 4.2375 252.32 4.3725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.045 4.2375 255.18 4.3725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.905 4.2375 258.04 4.3725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.765 4.2375 260.9 4.3725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.625 4.2375 263.76 4.3725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.485 4.2375 266.62 4.3725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.345 4.2375 269.48 4.3725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.205 4.2375 272.34 4.3725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.065 4.2375 275.2 4.3725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.925 4.2375 278.06 4.3725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.785 4.2375 280.92 4.3725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.645 4.2375 283.78 4.3725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.505 4.2375 286.64 4.3725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.365 4.2375 289.5 4.3725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.225 4.2375 292.36 4.3725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.085 4.2375 295.22 4.3725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.945 4.2375 298.08 4.3725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.805 4.2375 300.94 4.3725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.665 4.2375 303.8 4.3725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.525 4.2375 306.66 4.3725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.385 4.2375 309.52 4.3725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.245 4.2375 312.38 4.3725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.105 4.2375 315.24 4.3725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.965 4.2375 318.1 4.3725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.825 4.2375 320.96 4.3725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.685 4.2375 323.82 4.3725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.545 4.2375 326.68 4.3725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.405 4.2375 329.54 4.3725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.265 4.2375 332.4 4.3725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.125 4.2375 335.26 4.3725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.985 4.2375 338.12 4.3725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.845 4.2375 340.98 4.3725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.705 4.2375 343.84 4.3725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.565 4.2375 346.7 4.3725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.425 4.2375 349.56 4.3725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.285 4.2375 352.42 4.3725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.145 4.2375 355.28 4.3725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.005 4.2375 358.14 4.3725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.865 4.2375 361.0 4.3725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.725 4.2375 363.86 4.3725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.585 4.2375 366.72 4.3725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.445 4.2375 369.58 4.3725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.305 4.2375 372.44 4.3725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.165 4.2375 375.3 4.3725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.025 4.2375 378.16 4.3725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.885 4.2375 381.02 4.3725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.745 4.2375 383.88 4.3725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.605 4.2375 386.74 4.3725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.465 4.2375 389.6 4.3725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.325 4.2375 392.46 4.3725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.185 4.2375 395.32 4.3725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.045 4.2375 398.18 4.3725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.905 4.2375 401.04 4.3725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.765 4.2375 403.9 4.3725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.625 4.2375 406.76 4.3725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.485 4.2375 409.62 4.3725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.345 4.2375 412.48 4.3725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.205 4.2375 415.34 4.3725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.065 4.2375 418.2 4.3725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.925 4.2375 421.06 4.3725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.785 4.2375 423.92 4.3725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.645 4.2375 426.78 4.3725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.505 4.2375 429.64 4.3725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.365 4.2375 432.5 4.3725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.225 4.2375 435.36 4.3725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.085 4.2375 438.22 4.3725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.945 4.2375 441.08 4.3725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.805 4.2375 443.94 4.3725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.665 4.2375 446.8 4.3725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.525 4.2375 449.66 4.3725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.385 4.2375 452.52 4.3725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.245 4.2375 455.38 4.3725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.105 4.2375 458.24 4.3725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  460.965 4.2375 461.1 4.3725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  463.825 4.2375 463.96 4.3725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.685 4.2375 466.82 4.3725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.545 4.2375 469.68 4.3725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.405 4.2375 472.54 4.3725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.265 4.2375 475.4 4.3725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.125 4.2375 478.26 4.3725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  480.985 4.2375 481.12 4.3725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  483.845 4.2375 483.98 4.3725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.705 4.2375 486.84 4.3725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.565 4.2375 489.7 4.3725 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.425 4.2375 492.56 4.3725 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.285 4.2375 495.42 4.3725 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.145 4.2375 498.28 4.3725 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.005 4.2375 501.14 4.3725 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  503.865 4.2375 504.0 4.3725 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  506.725 4.2375 506.86 4.3725 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.585 4.2375 509.72 4.3725 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.445 4.2375 512.58 4.3725 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.305 4.2375 515.44 4.3725 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.165 4.2375 518.3 4.3725 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.025 4.2375 521.16 4.3725 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  523.885 4.2375 524.02 4.3725 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  526.745 4.2375 526.88 4.3725 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  529.605 4.2375 529.74 4.3725 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  532.465 4.2375 532.6 4.3725 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  535.325 4.2375 535.46 4.3725 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  538.185 4.2375 538.32 4.3725 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  541.045 4.2375 541.18 4.3725 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  543.905 4.2375 544.04 4.3725 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  546.765 4.2375 546.9 4.3725 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  549.625 4.2375 549.76 4.3725 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  552.485 4.2375 552.62 4.3725 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  555.345 4.2375 555.48 4.3725 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  558.205 4.2375 558.34 4.3725 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  561.065 4.2375 561.2 4.3725 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  563.925 4.2375 564.06 4.3725 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  566.785 4.2375 566.92 4.3725 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  569.645 4.2375 569.78 4.3725 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  572.505 4.2375 572.64 4.3725 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  575.365 4.2375 575.5 4.3725 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  578.225 4.2375 578.36 4.3725 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  581.085 4.2375 581.22 4.3725 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  583.945 4.2375 584.08 4.3725 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  586.805 4.2375 586.94 4.3725 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  589.665 4.2375 589.8 4.3725 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  592.525 4.2375 592.66 4.3725 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  595.385 4.2375 595.52 4.3725 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  598.245 4.2375 598.38 4.3725 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  601.105 4.2375 601.24 4.3725 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  603.965 4.2375 604.1 4.3725 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  606.825 4.2375 606.96 4.3725 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  609.685 4.2375 609.82 4.3725 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  612.545 4.2375 612.68 4.3725 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  615.405 4.2375 615.54 4.3725 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  618.265 4.2375 618.4 4.3725 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  621.125 4.2375 621.26 4.3725 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  623.985 4.2375 624.12 4.3725 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  626.845 4.2375 626.98 4.3725 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  629.705 4.2375 629.84 4.3725 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  632.565 4.2375 632.7 4.3725 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  635.425 4.2375 635.56 4.3725 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  638.285 4.2375 638.42 4.3725 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  641.145 4.2375 641.28 4.3725 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  644.005 4.2375 644.14 4.3725 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  646.865 4.2375 647.0 4.3725 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  649.725 4.2375 649.86 4.3725 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  652.585 4.2375 652.72 4.3725 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  655.445 4.2375 655.58 4.3725 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  658.305 4.2375 658.44 4.3725 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  661.165 4.2375 661.3 4.3725 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  664.025 4.2375 664.16 4.3725 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  666.885 4.2375 667.02 4.3725 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  669.745 4.2375 669.88 4.3725 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  672.605 4.2375 672.74 4.3725 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  675.465 4.2375 675.6 4.3725 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  678.325 4.2375 678.46 4.3725 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  681.185 4.2375 681.32 4.3725 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  684.045 4.2375 684.18 4.3725 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  686.905 4.2375 687.04 4.3725 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  689.765 4.2375 689.9 4.3725 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  692.625 4.2375 692.76 4.3725 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  695.485 4.2375 695.62 4.3725 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  698.345 4.2375 698.48 4.3725 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  701.205 4.2375 701.34 4.3725 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  704.065 4.2375 704.2 4.3725 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  706.925 4.2375 707.06 4.3725 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  709.785 4.2375 709.92 4.3725 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  712.645 4.2375 712.78 4.3725 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  715.505 4.2375 715.64 4.3725 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  718.365 4.2375 718.5 4.3725 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  721.225 4.2375 721.36 4.3725 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  724.085 4.2375 724.22 4.3725 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  726.945 4.2375 727.08 4.3725 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  729.805 4.2375 729.94 4.3725 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  732.665 4.2375 732.8 4.3725 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  735.525 4.2375 735.66 4.3725 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  738.385 4.2375 738.52 4.3725 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  741.245 4.2375 741.38 4.3725 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  744.105 4.2375 744.24 4.3725 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  746.965 4.2375 747.1 4.3725 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  749.825 4.2375 749.96 4.3725 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  752.685 4.2375 752.82 4.3725 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  755.545 4.2375 755.68 4.3725 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  758.405 4.2375 758.54 4.3725 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  761.265 4.2375 761.4 4.3725 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  764.125 4.2375 764.26 4.3725 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  766.985 4.2375 767.12 4.3725 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  769.845 4.2375 769.98 4.3725 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  772.705 4.2375 772.84 4.3725 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  775.565 4.2375 775.7 4.3725 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  778.425 4.2375 778.56 4.3725 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  781.285 4.2375 781.42 4.3725 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  784.145 4.2375 784.28 4.3725 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  787.005 4.2375 787.14 4.3725 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  789.865 4.2375 790.0 4.3725 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  792.725 4.2375 792.86 4.3725 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  795.585 4.2375 795.72 4.3725 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  798.445 4.2375 798.58 4.3725 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.305 4.2375 801.44 4.3725 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  804.165 4.2375 804.3 4.3725 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  807.025 4.2375 807.16 4.3725 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  809.885 4.2375 810.02 4.3725 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  812.745 4.2375 812.88 4.3725 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  815.605 4.2375 815.74 4.3725 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  818.465 4.2375 818.6 4.3725 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  821.325 4.2375 821.46 4.3725 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  824.185 4.2375 824.32 4.3725 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  827.045 4.2375 827.18 4.3725 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  829.905 4.2375 830.04 4.3725 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  832.765 4.2375 832.9 4.3725 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  835.625 4.2375 835.76 4.3725 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  838.485 4.2375 838.62 4.3725 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  841.345 4.2375 841.48 4.3725 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  844.205 4.2375 844.34 4.3725 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  847.065 4.2375 847.2 4.3725 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  849.925 4.2375 850.06 4.3725 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  852.785 4.2375 852.92 4.3725 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  855.645 4.2375 855.78 4.3725 ;
      END
   END din0[255]
   PIN din0[256]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  858.505 4.2375 858.64 4.3725 ;
      END
   END din0[256]
   PIN din0[257]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  861.365 4.2375 861.5 4.3725 ;
      END
   END din0[257]
   PIN din0[258]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  864.225 4.2375 864.36 4.3725 ;
      END
   END din0[258]
   PIN din0[259]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  867.085 4.2375 867.22 4.3725 ;
      END
   END din0[259]
   PIN din0[260]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  869.945 4.2375 870.08 4.3725 ;
      END
   END din0[260]
   PIN din0[261]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  872.805 4.2375 872.94 4.3725 ;
      END
   END din0[261]
   PIN din0[262]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  875.665 4.2375 875.8 4.3725 ;
      END
   END din0[262]
   PIN din0[263]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  878.525 4.2375 878.66 4.3725 ;
      END
   END din0[263]
   PIN din0[264]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  881.385 4.2375 881.52 4.3725 ;
      END
   END din0[264]
   PIN din0[265]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  884.245 4.2375 884.38 4.3725 ;
      END
   END din0[265]
   PIN din0[266]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  887.105 4.2375 887.24 4.3725 ;
      END
   END din0[266]
   PIN din0[267]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  889.965 4.2375 890.1 4.3725 ;
      END
   END din0[267]
   PIN din0[268]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  892.825 4.2375 892.96 4.3725 ;
      END
   END din0[268]
   PIN din0[269]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  895.685 4.2375 895.82 4.3725 ;
      END
   END din0[269]
   PIN din0[270]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  898.545 4.2375 898.68 4.3725 ;
      END
   END din0[270]
   PIN din0[271]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  901.405 4.2375 901.54 4.3725 ;
      END
   END din0[271]
   PIN din0[272]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  904.265 4.2375 904.4 4.3725 ;
      END
   END din0[272]
   PIN din0[273]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  907.125 4.2375 907.26 4.3725 ;
      END
   END din0[273]
   PIN din0[274]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  909.985 4.2375 910.12 4.3725 ;
      END
   END din0[274]
   PIN din0[275]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  912.845 4.2375 912.98 4.3725 ;
      END
   END din0[275]
   PIN din0[276]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  915.705 4.2375 915.84 4.3725 ;
      END
   END din0[276]
   PIN din0[277]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  918.565 4.2375 918.7 4.3725 ;
      END
   END din0[277]
   PIN din0[278]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  921.425 4.2375 921.56 4.3725 ;
      END
   END din0[278]
   PIN din0[279]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  924.285 4.2375 924.42 4.3725 ;
      END
   END din0[279]
   PIN din0[280]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  927.145 4.2375 927.28 4.3725 ;
      END
   END din0[280]
   PIN din0[281]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  930.005 4.2375 930.14 4.3725 ;
      END
   END din0[281]
   PIN din0[282]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  932.865 4.2375 933.0 4.3725 ;
      END
   END din0[282]
   PIN din0[283]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  935.725 4.2375 935.86 4.3725 ;
      END
   END din0[283]
   PIN din0[284]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  938.585 4.2375 938.72 4.3725 ;
      END
   END din0[284]
   PIN din0[285]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  941.445 4.2375 941.58 4.3725 ;
      END
   END din0[285]
   PIN din0[286]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  944.305 4.2375 944.44 4.3725 ;
      END
   END din0[286]
   PIN din0[287]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  947.165 4.2375 947.3 4.3725 ;
      END
   END din0[287]
   PIN din0[288]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  950.025 4.2375 950.16 4.3725 ;
      END
   END din0[288]
   PIN din0[289]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  952.885 4.2375 953.02 4.3725 ;
      END
   END din0[289]
   PIN din0[290]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  955.745 4.2375 955.88 4.3725 ;
      END
   END din0[290]
   PIN din0[291]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  958.605 4.2375 958.74 4.3725 ;
      END
   END din0[291]
   PIN din0[292]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  961.465 4.2375 961.6 4.3725 ;
      END
   END din0[292]
   PIN din0[293]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  964.325 4.2375 964.46 4.3725 ;
      END
   END din0[293]
   PIN din0[294]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  967.185 4.2375 967.32 4.3725 ;
      END
   END din0[294]
   PIN din0[295]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  970.045 4.2375 970.18 4.3725 ;
      END
   END din0[295]
   PIN din0[296]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  972.905 4.2375 973.04 4.3725 ;
      END
   END din0[296]
   PIN din0[297]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  975.765 4.2375 975.9 4.3725 ;
      END
   END din0[297]
   PIN din0[298]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  978.625 4.2375 978.76 4.3725 ;
      END
   END din0[298]
   PIN din0[299]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  981.485 4.2375 981.62 4.3725 ;
      END
   END din0[299]
   PIN din0[300]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  984.345 4.2375 984.48 4.3725 ;
      END
   END din0[300]
   PIN din0[301]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  987.205 4.2375 987.34 4.3725 ;
      END
   END din0[301]
   PIN din0[302]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  990.065 4.2375 990.2 4.3725 ;
      END
   END din0[302]
   PIN din0[303]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  992.925 4.2375 993.06 4.3725 ;
      END
   END din0[303]
   PIN din0[304]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  995.785 4.2375 995.92 4.3725 ;
      END
   END din0[304]
   PIN din0[305]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  998.645 4.2375 998.78 4.3725 ;
      END
   END din0[305]
   PIN din0[306]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1001.505 4.2375 1001.64 4.3725 ;
      END
   END din0[306]
   PIN din0[307]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1004.365 4.2375 1004.5 4.3725 ;
      END
   END din0[307]
   PIN din0[308]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1007.225 4.2375 1007.36 4.3725 ;
      END
   END din0[308]
   PIN din0[309]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1010.085 4.2375 1010.22 4.3725 ;
      END
   END din0[309]
   PIN din0[310]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1012.945 4.2375 1013.08 4.3725 ;
      END
   END din0[310]
   PIN din0[311]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1015.805 4.2375 1015.94 4.3725 ;
      END
   END din0[311]
   PIN din0[312]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1018.665 4.2375 1018.8 4.3725 ;
      END
   END din0[312]
   PIN din0[313]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1021.525 4.2375 1021.66 4.3725 ;
      END
   END din0[313]
   PIN din0[314]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1024.385 4.2375 1024.52 4.3725 ;
      END
   END din0[314]
   PIN din0[315]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1027.245 4.2375 1027.38 4.3725 ;
      END
   END din0[315]
   PIN din0[316]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1030.105 4.2375 1030.24 4.3725 ;
      END
   END din0[316]
   PIN din0[317]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1032.965 4.2375 1033.1 4.3725 ;
      END
   END din0[317]
   PIN din0[318]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1035.825 4.2375 1035.96 4.3725 ;
      END
   END din0[318]
   PIN din0[319]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1038.685 4.2375 1038.82 4.3725 ;
      END
   END din0[319]
   PIN din0[320]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1041.545 4.2375 1041.68 4.3725 ;
      END
   END din0[320]
   PIN din0[321]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1044.405 4.2375 1044.54 4.3725 ;
      END
   END din0[321]
   PIN din0[322]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1047.265 4.2375 1047.4 4.3725 ;
      END
   END din0[322]
   PIN din0[323]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1050.125 4.2375 1050.26 4.3725 ;
      END
   END din0[323]
   PIN din0[324]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1052.985 4.2375 1053.12 4.3725 ;
      END
   END din0[324]
   PIN din0[325]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1055.845 4.2375 1055.98 4.3725 ;
      END
   END din0[325]
   PIN din0[326]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1058.705 4.2375 1058.84 4.3725 ;
      END
   END din0[326]
   PIN din0[327]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1061.565 4.2375 1061.7 4.3725 ;
      END
   END din0[327]
   PIN din0[328]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1064.425 4.2375 1064.56 4.3725 ;
      END
   END din0[328]
   PIN din0[329]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1067.285 4.2375 1067.42 4.3725 ;
      END
   END din0[329]
   PIN din0[330]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1070.145 4.2375 1070.28 4.3725 ;
      END
   END din0[330]
   PIN din0[331]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1073.005 4.2375 1073.14 4.3725 ;
      END
   END din0[331]
   PIN din0[332]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1075.865 4.2375 1076.0 4.3725 ;
      END
   END din0[332]
   PIN din0[333]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1078.725 4.2375 1078.86 4.3725 ;
      END
   END din0[333]
   PIN din0[334]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1081.585 4.2375 1081.72 4.3725 ;
      END
   END din0[334]
   PIN din0[335]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1084.445 4.2375 1084.58 4.3725 ;
      END
   END din0[335]
   PIN din0[336]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1087.305 4.2375 1087.44 4.3725 ;
      END
   END din0[336]
   PIN din0[337]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1090.165 4.2375 1090.3 4.3725 ;
      END
   END din0[337]
   PIN din0[338]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1093.025 4.2375 1093.16 4.3725 ;
      END
   END din0[338]
   PIN din0[339]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1095.885 4.2375 1096.02 4.3725 ;
      END
   END din0[339]
   PIN din0[340]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1098.745 4.2375 1098.88 4.3725 ;
      END
   END din0[340]
   PIN din0[341]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1101.605 4.2375 1101.74 4.3725 ;
      END
   END din0[341]
   PIN din0[342]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1104.465 4.2375 1104.6 4.3725 ;
      END
   END din0[342]
   PIN din0[343]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1107.325 4.2375 1107.46 4.3725 ;
      END
   END din0[343]
   PIN din0[344]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1110.185 4.2375 1110.32 4.3725 ;
      END
   END din0[344]
   PIN din0[345]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1113.045 4.2375 1113.18 4.3725 ;
      END
   END din0[345]
   PIN din0[346]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1115.905 4.2375 1116.04 4.3725 ;
      END
   END din0[346]
   PIN din0[347]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1118.765 4.2375 1118.9 4.3725 ;
      END
   END din0[347]
   PIN din0[348]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1121.625 4.2375 1121.76 4.3725 ;
      END
   END din0[348]
   PIN din0[349]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1124.485 4.2375 1124.62 4.3725 ;
      END
   END din0[349]
   PIN din0[350]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1127.345 4.2375 1127.48 4.3725 ;
      END
   END din0[350]
   PIN din0[351]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1130.205 4.2375 1130.34 4.3725 ;
      END
   END din0[351]
   PIN din0[352]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1133.065 4.2375 1133.2 4.3725 ;
      END
   END din0[352]
   PIN din0[353]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1135.925 4.2375 1136.06 4.3725 ;
      END
   END din0[353]
   PIN din0[354]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1138.785 4.2375 1138.92 4.3725 ;
      END
   END din0[354]
   PIN din0[355]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1141.645 4.2375 1141.78 4.3725 ;
      END
   END din0[355]
   PIN din0[356]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1144.505 4.2375 1144.64 4.3725 ;
      END
   END din0[356]
   PIN din0[357]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1147.365 4.2375 1147.5 4.3725 ;
      END
   END din0[357]
   PIN din0[358]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1150.225 4.2375 1150.36 4.3725 ;
      END
   END din0[358]
   PIN din0[359]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1153.085 4.2375 1153.22 4.3725 ;
      END
   END din0[359]
   PIN din0[360]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1155.945 4.2375 1156.08 4.3725 ;
      END
   END din0[360]
   PIN din0[361]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1158.805 4.2375 1158.94 4.3725 ;
      END
   END din0[361]
   PIN din0[362]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1161.665 4.2375 1161.8 4.3725 ;
      END
   END din0[362]
   PIN din0[363]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1164.525 4.2375 1164.66 4.3725 ;
      END
   END din0[363]
   PIN din0[364]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1167.385 4.2375 1167.52 4.3725 ;
      END
   END din0[364]
   PIN din0[365]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1170.245 4.2375 1170.38 4.3725 ;
      END
   END din0[365]
   PIN din0[366]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1173.105 4.2375 1173.24 4.3725 ;
      END
   END din0[366]
   PIN din0[367]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1175.965 4.2375 1176.1 4.3725 ;
      END
   END din0[367]
   PIN din0[368]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1178.825 4.2375 1178.96 4.3725 ;
      END
   END din0[368]
   PIN din0[369]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1181.685 4.2375 1181.82 4.3725 ;
      END
   END din0[369]
   PIN din0[370]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1184.545 4.2375 1184.68 4.3725 ;
      END
   END din0[370]
   PIN din0[371]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1187.405 4.2375 1187.54 4.3725 ;
      END
   END din0[371]
   PIN din0[372]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1190.265 4.2375 1190.4 4.3725 ;
      END
   END din0[372]
   PIN din0[373]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1193.125 4.2375 1193.26 4.3725 ;
      END
   END din0[373]
   PIN din0[374]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1195.985 4.2375 1196.12 4.3725 ;
      END
   END din0[374]
   PIN din0[375]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1198.845 4.2375 1198.98 4.3725 ;
      END
   END din0[375]
   PIN din0[376]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1201.705 4.2375 1201.84 4.3725 ;
      END
   END din0[376]
   PIN din0[377]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1204.565 4.2375 1204.7 4.3725 ;
      END
   END din0[377]
   PIN din0[378]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1207.425 4.2375 1207.56 4.3725 ;
      END
   END din0[378]
   PIN din0[379]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1210.285 4.2375 1210.42 4.3725 ;
      END
   END din0[379]
   PIN din0[380]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1213.145 4.2375 1213.28 4.3725 ;
      END
   END din0[380]
   PIN din0[381]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1216.005 4.2375 1216.14 4.3725 ;
      END
   END din0[381]
   PIN din0[382]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1218.865 4.2375 1219.0 4.3725 ;
      END
   END din0[382]
   PIN din0[383]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1221.725 4.2375 1221.86 4.3725 ;
      END
   END din0[383]
   PIN din0[384]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1224.585 4.2375 1224.72 4.3725 ;
      END
   END din0[384]
   PIN din0[385]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1227.445 4.2375 1227.58 4.3725 ;
      END
   END din0[385]
   PIN din0[386]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1230.305 4.2375 1230.44 4.3725 ;
      END
   END din0[386]
   PIN din0[387]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1233.165 4.2375 1233.3 4.3725 ;
      END
   END din0[387]
   PIN din0[388]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1236.025 4.2375 1236.16 4.3725 ;
      END
   END din0[388]
   PIN din0[389]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1238.885 4.2375 1239.02 4.3725 ;
      END
   END din0[389]
   PIN din0[390]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1241.745 4.2375 1241.88 4.3725 ;
      END
   END din0[390]
   PIN din0[391]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1244.605 4.2375 1244.74 4.3725 ;
      END
   END din0[391]
   PIN din0[392]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1247.465 4.2375 1247.6 4.3725 ;
      END
   END din0[392]
   PIN din0[393]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1250.325 4.2375 1250.46 4.3725 ;
      END
   END din0[393]
   PIN din0[394]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1253.185 4.2375 1253.32 4.3725 ;
      END
   END din0[394]
   PIN din0[395]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1256.045 4.2375 1256.18 4.3725 ;
      END
   END din0[395]
   PIN din0[396]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1258.905 4.2375 1259.04 4.3725 ;
      END
   END din0[396]
   PIN din0[397]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1261.765 4.2375 1261.9 4.3725 ;
      END
   END din0[397]
   PIN din0[398]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1264.625 4.2375 1264.76 4.3725 ;
      END
   END din0[398]
   PIN din0[399]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1267.485 4.2375 1267.62 4.3725 ;
      END
   END din0[399]
   PIN din0[400]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1270.345 4.2375 1270.48 4.3725 ;
      END
   END din0[400]
   PIN din0[401]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1273.205 4.2375 1273.34 4.3725 ;
      END
   END din0[401]
   PIN din0[402]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1276.065 4.2375 1276.2 4.3725 ;
      END
   END din0[402]
   PIN din0[403]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1278.925 4.2375 1279.06 4.3725 ;
      END
   END din0[403]
   PIN din0[404]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1281.785 4.2375 1281.92 4.3725 ;
      END
   END din0[404]
   PIN din0[405]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1284.645 4.2375 1284.78 4.3725 ;
      END
   END din0[405]
   PIN din0[406]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1287.505 4.2375 1287.64 4.3725 ;
      END
   END din0[406]
   PIN din0[407]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1290.365 4.2375 1290.5 4.3725 ;
      END
   END din0[407]
   PIN din0[408]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1293.225 4.2375 1293.36 4.3725 ;
      END
   END din0[408]
   PIN din0[409]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1296.085 4.2375 1296.22 4.3725 ;
      END
   END din0[409]
   PIN din0[410]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1298.945 4.2375 1299.08 4.3725 ;
      END
   END din0[410]
   PIN din0[411]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1301.805 4.2375 1301.94 4.3725 ;
      END
   END din0[411]
   PIN din0[412]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1304.665 4.2375 1304.8 4.3725 ;
      END
   END din0[412]
   PIN din0[413]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1307.525 4.2375 1307.66 4.3725 ;
      END
   END din0[413]
   PIN din0[414]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1310.385 4.2375 1310.52 4.3725 ;
      END
   END din0[414]
   PIN din0[415]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1313.245 4.2375 1313.38 4.3725 ;
      END
   END din0[415]
   PIN din0[416]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1316.105 4.2375 1316.24 4.3725 ;
      END
   END din0[416]
   PIN din0[417]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1318.965 4.2375 1319.1 4.3725 ;
      END
   END din0[417]
   PIN din0[418]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1321.825 4.2375 1321.96 4.3725 ;
      END
   END din0[418]
   PIN din0[419]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1324.685 4.2375 1324.82 4.3725 ;
      END
   END din0[419]
   PIN din0[420]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1327.545 4.2375 1327.68 4.3725 ;
      END
   END din0[420]
   PIN din0[421]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1330.405 4.2375 1330.54 4.3725 ;
      END
   END din0[421]
   PIN din0[422]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1333.265 4.2375 1333.4 4.3725 ;
      END
   END din0[422]
   PIN din0[423]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1336.125 4.2375 1336.26 4.3725 ;
      END
   END din0[423]
   PIN din0[424]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1338.985 4.2375 1339.12 4.3725 ;
      END
   END din0[424]
   PIN din0[425]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1341.845 4.2375 1341.98 4.3725 ;
      END
   END din0[425]
   PIN din0[426]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1344.705 4.2375 1344.84 4.3725 ;
      END
   END din0[426]
   PIN din0[427]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1347.565 4.2375 1347.7 4.3725 ;
      END
   END din0[427]
   PIN din0[428]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1350.425 4.2375 1350.56 4.3725 ;
      END
   END din0[428]
   PIN din0[429]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1353.285 4.2375 1353.42 4.3725 ;
      END
   END din0[429]
   PIN din0[430]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1356.145 4.2375 1356.28 4.3725 ;
      END
   END din0[430]
   PIN din0[431]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1359.005 4.2375 1359.14 4.3725 ;
      END
   END din0[431]
   PIN din0[432]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1361.865 4.2375 1362.0 4.3725 ;
      END
   END din0[432]
   PIN din0[433]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1364.725 4.2375 1364.86 4.3725 ;
      END
   END din0[433]
   PIN din0[434]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1367.585 4.2375 1367.72 4.3725 ;
      END
   END din0[434]
   PIN din0[435]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1370.445 4.2375 1370.58 4.3725 ;
      END
   END din0[435]
   PIN din0[436]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1373.305 4.2375 1373.44 4.3725 ;
      END
   END din0[436]
   PIN din0[437]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1376.165 4.2375 1376.3 4.3725 ;
      END
   END din0[437]
   PIN din0[438]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1379.025 4.2375 1379.16 4.3725 ;
      END
   END din0[438]
   PIN din0[439]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1381.885 4.2375 1382.02 4.3725 ;
      END
   END din0[439]
   PIN din0[440]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1384.745 4.2375 1384.88 4.3725 ;
      END
   END din0[440]
   PIN din0[441]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1387.605 4.2375 1387.74 4.3725 ;
      END
   END din0[441]
   PIN din0[442]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1390.465 4.2375 1390.6 4.3725 ;
      END
   END din0[442]
   PIN din0[443]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1393.325 4.2375 1393.46 4.3725 ;
      END
   END din0[443]
   PIN din0[444]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1396.185 4.2375 1396.32 4.3725 ;
      END
   END din0[444]
   PIN din0[445]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1399.045 4.2375 1399.18 4.3725 ;
      END
   END din0[445]
   PIN din0[446]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1401.905 4.2375 1402.04 4.3725 ;
      END
   END din0[446]
   PIN din0[447]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1404.765 4.2375 1404.9 4.3725 ;
      END
   END din0[447]
   PIN din0[448]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1407.625 4.2375 1407.76 4.3725 ;
      END
   END din0[448]
   PIN din0[449]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1410.485 4.2375 1410.62 4.3725 ;
      END
   END din0[449]
   PIN din0[450]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1413.345 4.2375 1413.48 4.3725 ;
      END
   END din0[450]
   PIN din0[451]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1416.205 4.2375 1416.34 4.3725 ;
      END
   END din0[451]
   PIN din0[452]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1419.065 4.2375 1419.2 4.3725 ;
      END
   END din0[452]
   PIN din0[453]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1421.925 4.2375 1422.06 4.3725 ;
      END
   END din0[453]
   PIN din0[454]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1424.785 4.2375 1424.92 4.3725 ;
      END
   END din0[454]
   PIN din0[455]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1427.645 4.2375 1427.78 4.3725 ;
      END
   END din0[455]
   PIN din0[456]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1430.505 4.2375 1430.64 4.3725 ;
      END
   END din0[456]
   PIN din0[457]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1433.365 4.2375 1433.5 4.3725 ;
      END
   END din0[457]
   PIN din0[458]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1436.225 4.2375 1436.36 4.3725 ;
      END
   END din0[458]
   PIN din0[459]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1439.085 4.2375 1439.22 4.3725 ;
      END
   END din0[459]
   PIN din0[460]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1441.945 4.2375 1442.08 4.3725 ;
      END
   END din0[460]
   PIN din0[461]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1444.805 4.2375 1444.94 4.3725 ;
      END
   END din0[461]
   PIN din0[462]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1447.665 4.2375 1447.8 4.3725 ;
      END
   END din0[462]
   PIN din0[463]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1450.525 4.2375 1450.66 4.3725 ;
      END
   END din0[463]
   PIN din0[464]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1453.385 4.2375 1453.52 4.3725 ;
      END
   END din0[464]
   PIN din0[465]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1456.245 4.2375 1456.38 4.3725 ;
      END
   END din0[465]
   PIN din0[466]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1459.105 4.2375 1459.24 4.3725 ;
      END
   END din0[466]
   PIN din0[467]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1461.965 4.2375 1462.1 4.3725 ;
      END
   END din0[467]
   PIN din0[468]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1464.825 4.2375 1464.96 4.3725 ;
      END
   END din0[468]
   PIN din0[469]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1467.685 4.2375 1467.82 4.3725 ;
      END
   END din0[469]
   PIN din0[470]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1470.545 4.2375 1470.68 4.3725 ;
      END
   END din0[470]
   PIN din0[471]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1473.405 4.2375 1473.54 4.3725 ;
      END
   END din0[471]
   PIN din0[472]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1476.265 4.2375 1476.4 4.3725 ;
      END
   END din0[472]
   PIN din0[473]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1479.125 4.2375 1479.26 4.3725 ;
      END
   END din0[473]
   PIN din0[474]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1481.985 4.2375 1482.12 4.3725 ;
      END
   END din0[474]
   PIN din0[475]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1484.845 4.2375 1484.98 4.3725 ;
      END
   END din0[475]
   PIN din0[476]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1487.705 4.2375 1487.84 4.3725 ;
      END
   END din0[476]
   PIN din0[477]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1490.565 4.2375 1490.7 4.3725 ;
      END
   END din0[477]
   PIN din0[478]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1493.425 4.2375 1493.56 4.3725 ;
      END
   END din0[478]
   PIN din0[479]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1496.285 4.2375 1496.42 4.3725 ;
      END
   END din0[479]
   PIN din0[480]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1499.145 4.2375 1499.28 4.3725 ;
      END
   END din0[480]
   PIN din0[481]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1502.005 4.2375 1502.14 4.3725 ;
      END
   END din0[481]
   PIN din0[482]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1504.865 4.2375 1505.0 4.3725 ;
      END
   END din0[482]
   PIN din0[483]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1507.725 4.2375 1507.86 4.3725 ;
      END
   END din0[483]
   PIN din0[484]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1510.585 4.2375 1510.72 4.3725 ;
      END
   END din0[484]
   PIN din0[485]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1513.445 4.2375 1513.58 4.3725 ;
      END
   END din0[485]
   PIN din0[486]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1516.305 4.2375 1516.44 4.3725 ;
      END
   END din0[486]
   PIN din0[487]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1519.165 4.2375 1519.3 4.3725 ;
      END
   END din0[487]
   PIN din0[488]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1522.025 4.2375 1522.16 4.3725 ;
      END
   END din0[488]
   PIN din0[489]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1524.885 4.2375 1525.02 4.3725 ;
      END
   END din0[489]
   PIN din0[490]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1527.745 4.2375 1527.88 4.3725 ;
      END
   END din0[490]
   PIN din0[491]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1530.605 4.2375 1530.74 4.3725 ;
      END
   END din0[491]
   PIN din0[492]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1533.465 4.2375 1533.6 4.3725 ;
      END
   END din0[492]
   PIN din0[493]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1536.325 4.2375 1536.46 4.3725 ;
      END
   END din0[493]
   PIN din0[494]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1539.185 4.2375 1539.32 4.3725 ;
      END
   END din0[494]
   PIN din0[495]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1542.045 4.2375 1542.18 4.3725 ;
      END
   END din0[495]
   PIN din0[496]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1544.905 4.2375 1545.04 4.3725 ;
      END
   END din0[496]
   PIN din0[497]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1547.765 4.2375 1547.9 4.3725 ;
      END
   END din0[497]
   PIN din0[498]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1550.625 4.2375 1550.76 4.3725 ;
      END
   END din0[498]
   PIN din0[499]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1553.485 4.2375 1553.62 4.3725 ;
      END
   END din0[499]
   PIN din0[500]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1556.345 4.2375 1556.48 4.3725 ;
      END
   END din0[500]
   PIN din0[501]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1559.205 4.2375 1559.34 4.3725 ;
      END
   END din0[501]
   PIN din0[502]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1562.065 4.2375 1562.2 4.3725 ;
      END
   END din0[502]
   PIN din0[503]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1564.925 4.2375 1565.06 4.3725 ;
      END
   END din0[503]
   PIN din0[504]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1567.785 4.2375 1567.92 4.3725 ;
      END
   END din0[504]
   PIN din0[505]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1570.645 4.2375 1570.78 4.3725 ;
      END
   END din0[505]
   PIN din0[506]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1573.505 4.2375 1573.64 4.3725 ;
      END
   END din0[506]
   PIN din0[507]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1576.365 4.2375 1576.5 4.3725 ;
      END
   END din0[507]
   PIN din0[508]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1579.225 4.2375 1579.36 4.3725 ;
      END
   END din0[508]
   PIN din0[509]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1582.085 4.2375 1582.22 4.3725 ;
      END
   END din0[509]
   PIN din0[510]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1584.945 4.2375 1585.08 4.3725 ;
      END
   END din0[510]
   PIN din0[511]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1587.805 4.2375 1587.94 4.3725 ;
      END
   END din0[511]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.625 148.7225 120.76 148.8575 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.625 151.4525 120.76 151.5875 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.625 153.6625 120.76 153.7975 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.625 156.3925 120.76 156.5275 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.625 158.6025 120.76 158.7375 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.625 161.3325 120.76 161.4675 ;
      END
   END addr0[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  3.385 104.0025 3.52 104.1375 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  3.385 106.7325 3.52 106.8675 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.6275 104.0875 9.7625 104.2225 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.1125 115.65 163.2475 115.785 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.8175 115.65 163.9525 115.785 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.5225 115.65 164.6575 115.785 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.2275 115.65 165.3625 115.785 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.9325 115.65 166.0675 115.785 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.6375 115.65 166.7725 115.785 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.3425 115.65 167.4775 115.785 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.0475 115.65 168.1825 115.785 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.7525 115.65 168.8875 115.785 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.4575 115.65 169.5925 115.785 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.1625 115.65 170.2975 115.785 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.8675 115.65 171.0025 115.785 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.5725 115.65 171.7075 115.785 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.2775 115.65 172.4125 115.785 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.9825 115.65 173.1175 115.785 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.6875 115.65 173.8225 115.785 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.3925 115.65 174.5275 115.785 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.0975 115.65 175.2325 115.785 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.8025 115.65 175.9375 115.785 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.5075 115.65 176.6425 115.785 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.2125 115.65 177.3475 115.785 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.9175 115.65 178.0525 115.785 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.6225 115.65 178.7575 115.785 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.3275 115.65 179.4625 115.785 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.0325 115.65 180.1675 115.785 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.7375 115.65 180.8725 115.785 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.4425 115.65 181.5775 115.785 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.1475 115.65 182.2825 115.785 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.8525 115.65 182.9875 115.785 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.5575 115.65 183.6925 115.785 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.2625 115.65 184.3975 115.785 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.9675 115.65 185.1025 115.785 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.6725 115.65 185.8075 115.785 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.3775 115.65 186.5125 115.785 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.0825 115.65 187.2175 115.785 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.7875 115.65 187.9225 115.785 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.4925 115.65 188.6275 115.785 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.1975 115.65 189.3325 115.785 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.9025 115.65 190.0375 115.785 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.6075 115.65 190.7425 115.785 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.3125 115.65 191.4475 115.785 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.0175 115.65 192.1525 115.785 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.7225 115.65 192.8575 115.785 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.4275 115.65 193.5625 115.785 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.1325 115.65 194.2675 115.785 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.8375 115.65 194.9725 115.785 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.5425 115.65 195.6775 115.785 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.2475 115.65 196.3825 115.785 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.9525 115.65 197.0875 115.785 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.6575 115.65 197.7925 115.785 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.3625 115.65 198.4975 115.785 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.0675 115.65 199.2025 115.785 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.7725 115.65 199.9075 115.785 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.4775 115.65 200.6125 115.785 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.1825 115.65 201.3175 115.785 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.8875 115.65 202.0225 115.785 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.5925 115.65 202.7275 115.785 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.2975 115.65 203.4325 115.785 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.0025 115.65 204.1375 115.785 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.7075 115.65 204.8425 115.785 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.4125 115.65 205.5475 115.785 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.1175 115.65 206.2525 115.785 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.8225 115.65 206.9575 115.785 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.5275 115.65 207.6625 115.785 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.2325 115.65 208.3675 115.785 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.9375 115.65 209.0725 115.785 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.6425 115.65 209.7775 115.785 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.3475 115.65 210.4825 115.785 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.0525 115.65 211.1875 115.785 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.7575 115.65 211.8925 115.785 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.4625 115.65 212.5975 115.785 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.1675 115.65 213.3025 115.785 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.8725 115.65 214.0075 115.785 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.5775 115.65 214.7125 115.785 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.2825 115.65 215.4175 115.785 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.9875 115.65 216.1225 115.785 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.6925 115.65 216.8275 115.785 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.3975 115.65 217.5325 115.785 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.1025 115.65 218.2375 115.785 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.8075 115.65 218.9425 115.785 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.5125 115.65 219.6475 115.785 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.2175 115.65 220.3525 115.785 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.9225 115.65 221.0575 115.785 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.6275 115.65 221.7625 115.785 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.3325 115.65 222.4675 115.785 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.0375 115.65 223.1725 115.785 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.7425 115.65 223.8775 115.785 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.4475 115.65 224.5825 115.785 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.1525 115.65 225.2875 115.785 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.8575 115.65 225.9925 115.785 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.5625 115.65 226.6975 115.785 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.2675 115.65 227.4025 115.785 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.9725 115.65 228.1075 115.785 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.6775 115.65 228.8125 115.785 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.3825 115.65 229.5175 115.785 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.0875 115.65 230.2225 115.785 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.7925 115.65 230.9275 115.785 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.4975 115.65 231.6325 115.785 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.2025 115.65 232.3375 115.785 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.9075 115.65 233.0425 115.785 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.6125 115.65 233.7475 115.785 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.3175 115.65 234.4525 115.785 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.0225 115.65 235.1575 115.785 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.7275 115.65 235.8625 115.785 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.4325 115.65 236.5675 115.785 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.1375 115.65 237.2725 115.785 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.8425 115.65 237.9775 115.785 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.5475 115.65 238.6825 115.785 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.2525 115.65 239.3875 115.785 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.9575 115.65 240.0925 115.785 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.6625 115.65 240.7975 115.785 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.3675 115.65 241.5025 115.785 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.0725 115.65 242.2075 115.785 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.7775 115.65 242.9125 115.785 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.4825 115.65 243.6175 115.785 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.1875 115.65 244.3225 115.785 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.8925 115.65 245.0275 115.785 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.5975 115.65 245.7325 115.785 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.3025 115.65 246.4375 115.785 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.0075 115.65 247.1425 115.785 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.7125 115.65 247.8475 115.785 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.4175 115.65 248.5525 115.785 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.1225 115.65 249.2575 115.785 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.8275 115.65 249.9625 115.785 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.5325 115.65 250.6675 115.785 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.2375 115.65 251.3725 115.785 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.9425 115.65 252.0775 115.785 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.6475 115.65 252.7825 115.785 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.3525 115.65 253.4875 115.785 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.0575 115.65 254.1925 115.785 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.7625 115.65 254.8975 115.785 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.4675 115.65 255.6025 115.785 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.1725 115.65 256.3075 115.785 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.8775 115.65 257.0125 115.785 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.5825 115.65 257.7175 115.785 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.2875 115.65 258.4225 115.785 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.9925 115.65 259.1275 115.785 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.6975 115.65 259.8325 115.785 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.4025 115.65 260.5375 115.785 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.1075 115.65 261.2425 115.785 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.8125 115.65 261.9475 115.785 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.5175 115.65 262.6525 115.785 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.2225 115.65 263.3575 115.785 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.9275 115.65 264.0625 115.785 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.6325 115.65 264.7675 115.785 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.3375 115.65 265.4725 115.785 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.0425 115.65 266.1775 115.785 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.7475 115.65 266.8825 115.785 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.4525 115.65 267.5875 115.785 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.1575 115.65 268.2925 115.785 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.8625 115.65 268.9975 115.785 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.5675 115.65 269.7025 115.785 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.2725 115.65 270.4075 115.785 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.9775 115.65 271.1125 115.785 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.6825 115.65 271.8175 115.785 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.3875 115.65 272.5225 115.785 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.0925 115.65 273.2275 115.785 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.7975 115.65 273.9325 115.785 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.5025 115.65 274.6375 115.785 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.2075 115.65 275.3425 115.785 ;
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.9125 115.65 276.0475 115.785 ;
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.6175 115.65 276.7525 115.785 ;
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.3225 115.65 277.4575 115.785 ;
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.0275 115.65 278.1625 115.785 ;
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.7325 115.65 278.8675 115.785 ;
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.4375 115.65 279.5725 115.785 ;
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.1425 115.65 280.2775 115.785 ;
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.8475 115.65 280.9825 115.785 ;
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.5525 115.65 281.6875 115.785 ;
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  282.2575 115.65 282.3925 115.785 ;
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  282.9625 115.65 283.0975 115.785 ;
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.6675 115.65 283.8025 115.785 ;
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.3725 115.65 284.5075 115.785 ;
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.0775 115.65 285.2125 115.785 ;
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.7825 115.65 285.9175 115.785 ;
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.4875 115.65 286.6225 115.785 ;
      END
   END dout0[175]
   PIN dout0[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.1925 115.65 287.3275 115.785 ;
      END
   END dout0[176]
   PIN dout0[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.8975 115.65 288.0325 115.785 ;
      END
   END dout0[177]
   PIN dout0[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.6025 115.65 288.7375 115.785 ;
      END
   END dout0[178]
   PIN dout0[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.3075 115.65 289.4425 115.785 ;
      END
   END dout0[179]
   PIN dout0[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.0125 115.65 290.1475 115.785 ;
      END
   END dout0[180]
   PIN dout0[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.7175 115.65 290.8525 115.785 ;
      END
   END dout0[181]
   PIN dout0[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.4225 115.65 291.5575 115.785 ;
      END
   END dout0[182]
   PIN dout0[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.1275 115.65 292.2625 115.785 ;
      END
   END dout0[183]
   PIN dout0[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.8325 115.65 292.9675 115.785 ;
      END
   END dout0[184]
   PIN dout0[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.5375 115.65 293.6725 115.785 ;
      END
   END dout0[185]
   PIN dout0[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.2425 115.65 294.3775 115.785 ;
      END
   END dout0[186]
   PIN dout0[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.9475 115.65 295.0825 115.785 ;
      END
   END dout0[187]
   PIN dout0[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.6525 115.65 295.7875 115.785 ;
      END
   END dout0[188]
   PIN dout0[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.3575 115.65 296.4925 115.785 ;
      END
   END dout0[189]
   PIN dout0[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.0625 115.65 297.1975 115.785 ;
      END
   END dout0[190]
   PIN dout0[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.7675 115.65 297.9025 115.785 ;
      END
   END dout0[191]
   PIN dout0[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.4725 115.65 298.6075 115.785 ;
      END
   END dout0[192]
   PIN dout0[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.1775 115.65 299.3125 115.785 ;
      END
   END dout0[193]
   PIN dout0[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.8825 115.65 300.0175 115.785 ;
      END
   END dout0[194]
   PIN dout0[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.5875 115.65 300.7225 115.785 ;
      END
   END dout0[195]
   PIN dout0[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.2925 115.65 301.4275 115.785 ;
      END
   END dout0[196]
   PIN dout0[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.9975 115.65 302.1325 115.785 ;
      END
   END dout0[197]
   PIN dout0[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  302.7025 115.65 302.8375 115.785 ;
      END
   END dout0[198]
   PIN dout0[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.4075 115.65 303.5425 115.785 ;
      END
   END dout0[199]
   PIN dout0[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.1125 115.65 304.2475 115.785 ;
      END
   END dout0[200]
   PIN dout0[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.8175 115.65 304.9525 115.785 ;
      END
   END dout0[201]
   PIN dout0[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.5225 115.65 305.6575 115.785 ;
      END
   END dout0[202]
   PIN dout0[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.2275 115.65 306.3625 115.785 ;
      END
   END dout0[203]
   PIN dout0[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.9325 115.65 307.0675 115.785 ;
      END
   END dout0[204]
   PIN dout0[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.6375 115.65 307.7725 115.785 ;
      END
   END dout0[205]
   PIN dout0[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.3425 115.65 308.4775 115.785 ;
      END
   END dout0[206]
   PIN dout0[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.0475 115.65 309.1825 115.785 ;
      END
   END dout0[207]
   PIN dout0[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.7525 115.65 309.8875 115.785 ;
      END
   END dout0[208]
   PIN dout0[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.4575 115.65 310.5925 115.785 ;
      END
   END dout0[209]
   PIN dout0[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.1625 115.65 311.2975 115.785 ;
      END
   END dout0[210]
   PIN dout0[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.8675 115.65 312.0025 115.785 ;
      END
   END dout0[211]
   PIN dout0[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.5725 115.65 312.7075 115.785 ;
      END
   END dout0[212]
   PIN dout0[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.2775 115.65 313.4125 115.785 ;
      END
   END dout0[213]
   PIN dout0[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.9825 115.65 314.1175 115.785 ;
      END
   END dout0[214]
   PIN dout0[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.6875 115.65 314.8225 115.785 ;
      END
   END dout0[215]
   PIN dout0[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.3925 115.65 315.5275 115.785 ;
      END
   END dout0[216]
   PIN dout0[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.0975 115.65 316.2325 115.785 ;
      END
   END dout0[217]
   PIN dout0[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.8025 115.65 316.9375 115.785 ;
      END
   END dout0[218]
   PIN dout0[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.5075 115.65 317.6425 115.785 ;
      END
   END dout0[219]
   PIN dout0[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.2125 115.65 318.3475 115.785 ;
      END
   END dout0[220]
   PIN dout0[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.9175 115.65 319.0525 115.785 ;
      END
   END dout0[221]
   PIN dout0[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.6225 115.65 319.7575 115.785 ;
      END
   END dout0[222]
   PIN dout0[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.3275 115.65 320.4625 115.785 ;
      END
   END dout0[223]
   PIN dout0[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.0325 115.65 321.1675 115.785 ;
      END
   END dout0[224]
   PIN dout0[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.7375 115.65 321.8725 115.785 ;
      END
   END dout0[225]
   PIN dout0[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  322.4425 115.65 322.5775 115.785 ;
      END
   END dout0[226]
   PIN dout0[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.1475 115.65 323.2825 115.785 ;
      END
   END dout0[227]
   PIN dout0[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.8525 115.65 323.9875 115.785 ;
      END
   END dout0[228]
   PIN dout0[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.5575 115.65 324.6925 115.785 ;
      END
   END dout0[229]
   PIN dout0[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.2625 115.65 325.3975 115.785 ;
      END
   END dout0[230]
   PIN dout0[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.9675 115.65 326.1025 115.785 ;
      END
   END dout0[231]
   PIN dout0[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.6725 115.65 326.8075 115.785 ;
      END
   END dout0[232]
   PIN dout0[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.3775 115.65 327.5125 115.785 ;
      END
   END dout0[233]
   PIN dout0[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.0825 115.65 328.2175 115.785 ;
      END
   END dout0[234]
   PIN dout0[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.7875 115.65 328.9225 115.785 ;
      END
   END dout0[235]
   PIN dout0[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.4925 115.65 329.6275 115.785 ;
      END
   END dout0[236]
   PIN dout0[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.1975 115.65 330.3325 115.785 ;
      END
   END dout0[237]
   PIN dout0[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.9025 115.65 331.0375 115.785 ;
      END
   END dout0[238]
   PIN dout0[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.6075 115.65 331.7425 115.785 ;
      END
   END dout0[239]
   PIN dout0[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.3125 115.65 332.4475 115.785 ;
      END
   END dout0[240]
   PIN dout0[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.0175 115.65 333.1525 115.785 ;
      END
   END dout0[241]
   PIN dout0[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.7225 115.65 333.8575 115.785 ;
      END
   END dout0[242]
   PIN dout0[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.4275 115.65 334.5625 115.785 ;
      END
   END dout0[243]
   PIN dout0[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.1325 115.65 335.2675 115.785 ;
      END
   END dout0[244]
   PIN dout0[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.8375 115.65 335.9725 115.785 ;
      END
   END dout0[245]
   PIN dout0[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.5425 115.65 336.6775 115.785 ;
      END
   END dout0[246]
   PIN dout0[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.2475 115.65 337.3825 115.785 ;
      END
   END dout0[247]
   PIN dout0[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.9525 115.65 338.0875 115.785 ;
      END
   END dout0[248]
   PIN dout0[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.6575 115.65 338.7925 115.785 ;
      END
   END dout0[249]
   PIN dout0[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.3625 115.65 339.4975 115.785 ;
      END
   END dout0[250]
   PIN dout0[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.0675 115.65 340.2025 115.785 ;
      END
   END dout0[251]
   PIN dout0[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.7725 115.65 340.9075 115.785 ;
      END
   END dout0[252]
   PIN dout0[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.4775 115.65 341.6125 115.785 ;
      END
   END dout0[253]
   PIN dout0[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.1825 115.65 342.3175 115.785 ;
      END
   END dout0[254]
   PIN dout0[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.8875 115.65 343.0225 115.785 ;
      END
   END dout0[255]
   PIN dout0[256]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.5925 115.65 343.7275 115.785 ;
      END
   END dout0[256]
   PIN dout0[257]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.2975 115.65 344.4325 115.785 ;
      END
   END dout0[257]
   PIN dout0[258]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.0025 115.65 345.1375 115.785 ;
      END
   END dout0[258]
   PIN dout0[259]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.7075 115.65 345.8425 115.785 ;
      END
   END dout0[259]
   PIN dout0[260]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.4125 115.65 346.5475 115.785 ;
      END
   END dout0[260]
   PIN dout0[261]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.1175 115.65 347.2525 115.785 ;
      END
   END dout0[261]
   PIN dout0[262]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.8225 115.65 347.9575 115.785 ;
      END
   END dout0[262]
   PIN dout0[263]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.5275 115.65 348.6625 115.785 ;
      END
   END dout0[263]
   PIN dout0[264]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.2325 115.65 349.3675 115.785 ;
      END
   END dout0[264]
   PIN dout0[265]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.9375 115.65 350.0725 115.785 ;
      END
   END dout0[265]
   PIN dout0[266]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.6425 115.65 350.7775 115.785 ;
      END
   END dout0[266]
   PIN dout0[267]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  351.3475 115.65 351.4825 115.785 ;
      END
   END dout0[267]
   PIN dout0[268]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.0525 115.65 352.1875 115.785 ;
      END
   END dout0[268]
   PIN dout0[269]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.7575 115.65 352.8925 115.785 ;
      END
   END dout0[269]
   PIN dout0[270]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.4625 115.65 353.5975 115.785 ;
      END
   END dout0[270]
   PIN dout0[271]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.1675 115.65 354.3025 115.785 ;
      END
   END dout0[271]
   PIN dout0[272]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.8725 115.65 355.0075 115.785 ;
      END
   END dout0[272]
   PIN dout0[273]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.5775 115.65 355.7125 115.785 ;
      END
   END dout0[273]
   PIN dout0[274]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.2825 115.65 356.4175 115.785 ;
      END
   END dout0[274]
   PIN dout0[275]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.9875 115.65 357.1225 115.785 ;
      END
   END dout0[275]
   PIN dout0[276]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.6925 115.65 357.8275 115.785 ;
      END
   END dout0[276]
   PIN dout0[277]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.3975 115.65 358.5325 115.785 ;
      END
   END dout0[277]
   PIN dout0[278]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.1025 115.65 359.2375 115.785 ;
      END
   END dout0[278]
   PIN dout0[279]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.8075 115.65 359.9425 115.785 ;
      END
   END dout0[279]
   PIN dout0[280]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.5125 115.65 360.6475 115.785 ;
      END
   END dout0[280]
   PIN dout0[281]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.2175 115.65 361.3525 115.785 ;
      END
   END dout0[281]
   PIN dout0[282]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.9225 115.65 362.0575 115.785 ;
      END
   END dout0[282]
   PIN dout0[283]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.6275 115.65 362.7625 115.785 ;
      END
   END dout0[283]
   PIN dout0[284]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.3325 115.65 363.4675 115.785 ;
      END
   END dout0[284]
   PIN dout0[285]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.0375 115.65 364.1725 115.785 ;
      END
   END dout0[285]
   PIN dout0[286]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.7425 115.65 364.8775 115.785 ;
      END
   END dout0[286]
   PIN dout0[287]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.4475 115.65 365.5825 115.785 ;
      END
   END dout0[287]
   PIN dout0[288]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.1525 115.65 366.2875 115.785 ;
      END
   END dout0[288]
   PIN dout0[289]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.8575 115.65 366.9925 115.785 ;
      END
   END dout0[289]
   PIN dout0[290]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.5625 115.65 367.6975 115.785 ;
      END
   END dout0[290]
   PIN dout0[291]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.2675 115.65 368.4025 115.785 ;
      END
   END dout0[291]
   PIN dout0[292]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.9725 115.65 369.1075 115.785 ;
      END
   END dout0[292]
   PIN dout0[293]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.6775 115.65 369.8125 115.785 ;
      END
   END dout0[293]
   PIN dout0[294]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.3825 115.65 370.5175 115.785 ;
      END
   END dout0[294]
   PIN dout0[295]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  371.0875 115.65 371.2225 115.785 ;
      END
   END dout0[295]
   PIN dout0[296]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  371.7925 115.65 371.9275 115.785 ;
      END
   END dout0[296]
   PIN dout0[297]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.4975 115.65 372.6325 115.785 ;
      END
   END dout0[297]
   PIN dout0[298]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.2025 115.65 373.3375 115.785 ;
      END
   END dout0[298]
   PIN dout0[299]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.9075 115.65 374.0425 115.785 ;
      END
   END dout0[299]
   PIN dout0[300]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.6125 115.65 374.7475 115.785 ;
      END
   END dout0[300]
   PIN dout0[301]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.3175 115.65 375.4525 115.785 ;
      END
   END dout0[301]
   PIN dout0[302]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  376.0225 115.65 376.1575 115.785 ;
      END
   END dout0[302]
   PIN dout0[303]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  376.7275 115.65 376.8625 115.785 ;
      END
   END dout0[303]
   PIN dout0[304]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.4325 115.65 377.5675 115.785 ;
      END
   END dout0[304]
   PIN dout0[305]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.1375 115.65 378.2725 115.785 ;
      END
   END dout0[305]
   PIN dout0[306]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.8425 115.65 378.9775 115.785 ;
      END
   END dout0[306]
   PIN dout0[307]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  379.5475 115.65 379.6825 115.785 ;
      END
   END dout0[307]
   PIN dout0[308]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.2525 115.65 380.3875 115.785 ;
      END
   END dout0[308]
   PIN dout0[309]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.9575 115.65 381.0925 115.785 ;
      END
   END dout0[309]
   PIN dout0[310]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.6625 115.65 381.7975 115.785 ;
      END
   END dout0[310]
   PIN dout0[311]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  382.3675 115.65 382.5025 115.785 ;
      END
   END dout0[311]
   PIN dout0[312]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.0725 115.65 383.2075 115.785 ;
      END
   END dout0[312]
   PIN dout0[313]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.7775 115.65 383.9125 115.785 ;
      END
   END dout0[313]
   PIN dout0[314]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.4825 115.65 384.6175 115.785 ;
      END
   END dout0[314]
   PIN dout0[315]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  385.1875 115.65 385.3225 115.785 ;
      END
   END dout0[315]
   PIN dout0[316]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  385.8925 115.65 386.0275 115.785 ;
      END
   END dout0[316]
   PIN dout0[317]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.5975 115.65 386.7325 115.785 ;
      END
   END dout0[317]
   PIN dout0[318]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  387.3025 115.65 387.4375 115.785 ;
      END
   END dout0[318]
   PIN dout0[319]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  388.0075 115.65 388.1425 115.785 ;
      END
   END dout0[319]
   PIN dout0[320]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  388.7125 115.65 388.8475 115.785 ;
      END
   END dout0[320]
   PIN dout0[321]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.4175 115.65 389.5525 115.785 ;
      END
   END dout0[321]
   PIN dout0[322]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  390.1225 115.65 390.2575 115.785 ;
      END
   END dout0[322]
   PIN dout0[323]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  390.8275 115.65 390.9625 115.785 ;
      END
   END dout0[323]
   PIN dout0[324]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  391.5325 115.65 391.6675 115.785 ;
      END
   END dout0[324]
   PIN dout0[325]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.2375 115.65 392.3725 115.785 ;
      END
   END dout0[325]
   PIN dout0[326]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.9425 115.65 393.0775 115.785 ;
      END
   END dout0[326]
   PIN dout0[327]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.6475 115.65 393.7825 115.785 ;
      END
   END dout0[327]
   PIN dout0[328]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.3525 115.65 394.4875 115.785 ;
      END
   END dout0[328]
   PIN dout0[329]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.0575 115.65 395.1925 115.785 ;
      END
   END dout0[329]
   PIN dout0[330]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.7625 115.65 395.8975 115.785 ;
      END
   END dout0[330]
   PIN dout0[331]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.4675 115.65 396.6025 115.785 ;
      END
   END dout0[331]
   PIN dout0[332]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.1725 115.65 397.3075 115.785 ;
      END
   END dout0[332]
   PIN dout0[333]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.8775 115.65 398.0125 115.785 ;
      END
   END dout0[333]
   PIN dout0[334]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.5825 115.65 398.7175 115.785 ;
      END
   END dout0[334]
   PIN dout0[335]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.2875 115.65 399.4225 115.785 ;
      END
   END dout0[335]
   PIN dout0[336]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.9925 115.65 400.1275 115.785 ;
      END
   END dout0[336]
   PIN dout0[337]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.6975 115.65 400.8325 115.785 ;
      END
   END dout0[337]
   PIN dout0[338]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.4025 115.65 401.5375 115.785 ;
      END
   END dout0[338]
   PIN dout0[339]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  402.1075 115.65 402.2425 115.785 ;
      END
   END dout0[339]
   PIN dout0[340]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  402.8125 115.65 402.9475 115.785 ;
      END
   END dout0[340]
   PIN dout0[341]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.5175 115.65 403.6525 115.785 ;
      END
   END dout0[341]
   PIN dout0[342]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.2225 115.65 404.3575 115.785 ;
      END
   END dout0[342]
   PIN dout0[343]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.9275 115.65 405.0625 115.785 ;
      END
   END dout0[343]
   PIN dout0[344]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  405.6325 115.65 405.7675 115.785 ;
      END
   END dout0[344]
   PIN dout0[345]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.3375 115.65 406.4725 115.785 ;
      END
   END dout0[345]
   PIN dout0[346]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.0425 115.65 407.1775 115.785 ;
      END
   END dout0[346]
   PIN dout0[347]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.7475 115.65 407.8825 115.785 ;
      END
   END dout0[347]
   PIN dout0[348]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  408.4525 115.65 408.5875 115.785 ;
      END
   END dout0[348]
   PIN dout0[349]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.1575 115.65 409.2925 115.785 ;
      END
   END dout0[349]
   PIN dout0[350]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.8625 115.65 409.9975 115.785 ;
      END
   END dout0[350]
   PIN dout0[351]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.5675 115.65 410.7025 115.785 ;
      END
   END dout0[351]
   PIN dout0[352]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  411.2725 115.65 411.4075 115.785 ;
      END
   END dout0[352]
   PIN dout0[353]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  411.9775 115.65 412.1125 115.785 ;
      END
   END dout0[353]
   PIN dout0[354]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.6825 115.65 412.8175 115.785 ;
      END
   END dout0[354]
   PIN dout0[355]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  413.3875 115.65 413.5225 115.785 ;
      END
   END dout0[355]
   PIN dout0[356]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  414.0925 115.65 414.2275 115.785 ;
      END
   END dout0[356]
   PIN dout0[357]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  414.7975 115.65 414.9325 115.785 ;
      END
   END dout0[357]
   PIN dout0[358]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.5025 115.65 415.6375 115.785 ;
      END
   END dout0[358]
   PIN dout0[359]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  416.2075 115.65 416.3425 115.785 ;
      END
   END dout0[359]
   PIN dout0[360]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  416.9125 115.65 417.0475 115.785 ;
      END
   END dout0[360]
   PIN dout0[361]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.6175 115.65 417.7525 115.785 ;
      END
   END dout0[361]
   PIN dout0[362]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.3225 115.65 418.4575 115.785 ;
      END
   END dout0[362]
   PIN dout0[363]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  419.0275 115.65 419.1625 115.785 ;
      END
   END dout0[363]
   PIN dout0[364]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  419.7325 115.65 419.8675 115.785 ;
      END
   END dout0[364]
   PIN dout0[365]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.4375 115.65 420.5725 115.785 ;
      END
   END dout0[365]
   PIN dout0[366]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.1425 115.65 421.2775 115.785 ;
      END
   END dout0[366]
   PIN dout0[367]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.8475 115.65 421.9825 115.785 ;
      END
   END dout0[367]
   PIN dout0[368]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  422.5525 115.65 422.6875 115.785 ;
      END
   END dout0[368]
   PIN dout0[369]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.2575 115.65 423.3925 115.785 ;
      END
   END dout0[369]
   PIN dout0[370]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.9625 115.65 424.0975 115.785 ;
      END
   END dout0[370]
   PIN dout0[371]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.6675 115.65 424.8025 115.785 ;
      END
   END dout0[371]
   PIN dout0[372]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  425.3725 115.65 425.5075 115.785 ;
      END
   END dout0[372]
   PIN dout0[373]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.0775 115.65 426.2125 115.785 ;
      END
   END dout0[373]
   PIN dout0[374]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.7825 115.65 426.9175 115.785 ;
      END
   END dout0[374]
   PIN dout0[375]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.4875 115.65 427.6225 115.785 ;
      END
   END dout0[375]
   PIN dout0[376]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  428.1925 115.65 428.3275 115.785 ;
      END
   END dout0[376]
   PIN dout0[377]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  428.8975 115.65 429.0325 115.785 ;
      END
   END dout0[377]
   PIN dout0[378]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.6025 115.65 429.7375 115.785 ;
      END
   END dout0[378]
   PIN dout0[379]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  430.3075 115.65 430.4425 115.785 ;
      END
   END dout0[379]
   PIN dout0[380]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  431.0125 115.65 431.1475 115.785 ;
      END
   END dout0[380]
   PIN dout0[381]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  431.7175 115.65 431.8525 115.785 ;
      END
   END dout0[381]
   PIN dout0[382]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.4225 115.65 432.5575 115.785 ;
      END
   END dout0[382]
   PIN dout0[383]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  433.1275 115.65 433.2625 115.785 ;
      END
   END dout0[383]
   PIN dout0[384]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  433.8325 115.65 433.9675 115.785 ;
      END
   END dout0[384]
   PIN dout0[385]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  434.5375 115.65 434.6725 115.785 ;
      END
   END dout0[385]
   PIN dout0[386]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.2425 115.65 435.3775 115.785 ;
      END
   END dout0[386]
   PIN dout0[387]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.9475 115.65 436.0825 115.785 ;
      END
   END dout0[387]
   PIN dout0[388]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  436.6525 115.65 436.7875 115.785 ;
      END
   END dout0[388]
   PIN dout0[389]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  437.3575 115.65 437.4925 115.785 ;
      END
   END dout0[389]
   PIN dout0[390]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.0625 115.65 438.1975 115.785 ;
      END
   END dout0[390]
   PIN dout0[391]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.7675 115.65 438.9025 115.785 ;
      END
   END dout0[391]
   PIN dout0[392]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  439.4725 115.65 439.6075 115.785 ;
      END
   END dout0[392]
   PIN dout0[393]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.1775 115.65 440.3125 115.785 ;
      END
   END dout0[393]
   PIN dout0[394]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.8825 115.65 441.0175 115.785 ;
      END
   END dout0[394]
   PIN dout0[395]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.5875 115.65 441.7225 115.785 ;
      END
   END dout0[395]
   PIN dout0[396]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  442.2925 115.65 442.4275 115.785 ;
      END
   END dout0[396]
   PIN dout0[397]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  442.9975 115.65 443.1325 115.785 ;
      END
   END dout0[397]
   PIN dout0[398]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.7025 115.65 443.8375 115.785 ;
      END
   END dout0[398]
   PIN dout0[399]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.4075 115.65 444.5425 115.785 ;
      END
   END dout0[399]
   PIN dout0[400]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  445.1125 115.65 445.2475 115.785 ;
      END
   END dout0[400]
   PIN dout0[401]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  445.8175 115.65 445.9525 115.785 ;
      END
   END dout0[401]
   PIN dout0[402]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.5225 115.65 446.6575 115.785 ;
      END
   END dout0[402]
   PIN dout0[403]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.2275 115.65 447.3625 115.785 ;
      END
   END dout0[403]
   PIN dout0[404]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.9325 115.65 448.0675 115.785 ;
      END
   END dout0[404]
   PIN dout0[405]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  448.6375 115.65 448.7725 115.785 ;
      END
   END dout0[405]
   PIN dout0[406]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.3425 115.65 449.4775 115.785 ;
      END
   END dout0[406]
   PIN dout0[407]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  450.0475 115.65 450.1825 115.785 ;
      END
   END dout0[407]
   PIN dout0[408]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  450.7525 115.65 450.8875 115.785 ;
      END
   END dout0[408]
   PIN dout0[409]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  451.4575 115.65 451.5925 115.785 ;
      END
   END dout0[409]
   PIN dout0[410]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.1625 115.65 452.2975 115.785 ;
      END
   END dout0[410]
   PIN dout0[411]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.8675 115.65 453.0025 115.785 ;
      END
   END dout0[411]
   PIN dout0[412]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.5725 115.65 453.7075 115.785 ;
      END
   END dout0[412]
   PIN dout0[413]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  454.2775 115.65 454.4125 115.785 ;
      END
   END dout0[413]
   PIN dout0[414]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  454.9825 115.65 455.1175 115.785 ;
      END
   END dout0[414]
   PIN dout0[415]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.6875 115.65 455.8225 115.785 ;
      END
   END dout0[415]
   PIN dout0[416]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  456.3925 115.65 456.5275 115.785 ;
      END
   END dout0[416]
   PIN dout0[417]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  457.0975 115.65 457.2325 115.785 ;
      END
   END dout0[417]
   PIN dout0[418]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  457.8025 115.65 457.9375 115.785 ;
      END
   END dout0[418]
   PIN dout0[419]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.5075 115.65 458.6425 115.785 ;
      END
   END dout0[419]
   PIN dout0[420]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  459.2125 115.65 459.3475 115.785 ;
      END
   END dout0[420]
   PIN dout0[421]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  459.9175 115.65 460.0525 115.785 ;
      END
   END dout0[421]
   PIN dout0[422]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  460.6225 115.65 460.7575 115.785 ;
      END
   END dout0[422]
   PIN dout0[423]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.3275 115.65 461.4625 115.785 ;
      END
   END dout0[423]
   PIN dout0[424]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  462.0325 115.65 462.1675 115.785 ;
      END
   END dout0[424]
   PIN dout0[425]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  462.7375 115.65 462.8725 115.785 ;
      END
   END dout0[425]
   PIN dout0[426]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  463.4425 115.65 463.5775 115.785 ;
      END
   END dout0[426]
   PIN dout0[427]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.1475 115.65 464.2825 115.785 ;
      END
   END dout0[427]
   PIN dout0[428]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.8525 115.65 464.9875 115.785 ;
      END
   END dout0[428]
   PIN dout0[429]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  465.5575 115.65 465.6925 115.785 ;
      END
   END dout0[429]
   PIN dout0[430]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.2625 115.65 466.3975 115.785 ;
      END
   END dout0[430]
   PIN dout0[431]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.9675 115.65 467.1025 115.785 ;
      END
   END dout0[431]
   PIN dout0[432]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.6725 115.65 467.8075 115.785 ;
      END
   END dout0[432]
   PIN dout0[433]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  468.3775 115.65 468.5125 115.785 ;
      END
   END dout0[433]
   PIN dout0[434]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.0825 115.65 469.2175 115.785 ;
      END
   END dout0[434]
   PIN dout0[435]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.7875 115.65 469.9225 115.785 ;
      END
   END dout0[435]
   PIN dout0[436]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.4925 115.65 470.6275 115.785 ;
      END
   END dout0[436]
   PIN dout0[437]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  471.1975 115.65 471.3325 115.785 ;
      END
   END dout0[437]
   PIN dout0[438]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  471.9025 115.65 472.0375 115.785 ;
      END
   END dout0[438]
   PIN dout0[439]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.6075 115.65 472.7425 115.785 ;
      END
   END dout0[439]
   PIN dout0[440]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  473.3125 115.65 473.4475 115.785 ;
      END
   END dout0[440]
   PIN dout0[441]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  474.0175 115.65 474.1525 115.785 ;
      END
   END dout0[441]
   PIN dout0[442]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  474.7225 115.65 474.8575 115.785 ;
      END
   END dout0[442]
   PIN dout0[443]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.4275 115.65 475.5625 115.785 ;
      END
   END dout0[443]
   PIN dout0[444]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  476.1325 115.65 476.2675 115.785 ;
      END
   END dout0[444]
   PIN dout0[445]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  476.8375 115.65 476.9725 115.785 ;
      END
   END dout0[445]
   PIN dout0[446]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  477.5425 115.65 477.6775 115.785 ;
      END
   END dout0[446]
   PIN dout0[447]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.2475 115.65 478.3825 115.785 ;
      END
   END dout0[447]
   PIN dout0[448]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.9525 115.65 479.0875 115.785 ;
      END
   END dout0[448]
   PIN dout0[449]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  479.6575 115.65 479.7925 115.785 ;
      END
   END dout0[449]
   PIN dout0[450]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  480.3625 115.65 480.4975 115.785 ;
      END
   END dout0[450]
   PIN dout0[451]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.0675 115.65 481.2025 115.785 ;
      END
   END dout0[451]
   PIN dout0[452]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.7725 115.65 481.9075 115.785 ;
      END
   END dout0[452]
   PIN dout0[453]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.4775 115.65 482.6125 115.785 ;
      END
   END dout0[453]
   PIN dout0[454]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  483.1825 115.65 483.3175 115.785 ;
      END
   END dout0[454]
   PIN dout0[455]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  483.8875 115.65 484.0225 115.785 ;
      END
   END dout0[455]
   PIN dout0[456]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.5925 115.65 484.7275 115.785 ;
      END
   END dout0[456]
   PIN dout0[457]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  485.2975 115.65 485.4325 115.785 ;
      END
   END dout0[457]
   PIN dout0[458]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.0025 115.65 486.1375 115.785 ;
      END
   END dout0[458]
   PIN dout0[459]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.7075 115.65 486.8425 115.785 ;
      END
   END dout0[459]
   PIN dout0[460]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.4125 115.65 487.5475 115.785 ;
      END
   END dout0[460]
   PIN dout0[461]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  488.1175 115.65 488.2525 115.785 ;
      END
   END dout0[461]
   PIN dout0[462]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  488.8225 115.65 488.9575 115.785 ;
      END
   END dout0[462]
   PIN dout0[463]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.5275 115.65 489.6625 115.785 ;
      END
   END dout0[463]
   PIN dout0[464]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  490.2325 115.65 490.3675 115.785 ;
      END
   END dout0[464]
   PIN dout0[465]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  490.9375 115.65 491.0725 115.785 ;
      END
   END dout0[465]
   PIN dout0[466]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  491.6425 115.65 491.7775 115.785 ;
      END
   END dout0[466]
   PIN dout0[467]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.3475 115.65 492.4825 115.785 ;
      END
   END dout0[467]
   PIN dout0[468]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  493.0525 115.65 493.1875 115.785 ;
      END
   END dout0[468]
   PIN dout0[469]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  493.7575 115.65 493.8925 115.785 ;
      END
   END dout0[469]
   PIN dout0[470]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  494.4625 115.65 494.5975 115.785 ;
      END
   END dout0[470]
   PIN dout0[471]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.1675 115.65 495.3025 115.785 ;
      END
   END dout0[471]
   PIN dout0[472]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.8725 115.65 496.0075 115.785 ;
      END
   END dout0[472]
   PIN dout0[473]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  496.5775 115.65 496.7125 115.785 ;
      END
   END dout0[473]
   PIN dout0[474]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  497.2825 115.65 497.4175 115.785 ;
      END
   END dout0[474]
   PIN dout0[475]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  497.9875 115.65 498.1225 115.785 ;
      END
   END dout0[475]
   PIN dout0[476]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.6925 115.65 498.8275 115.785 ;
      END
   END dout0[476]
   PIN dout0[477]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  499.3975 115.65 499.5325 115.785 ;
      END
   END dout0[477]
   PIN dout0[478]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  500.1025 115.65 500.2375 115.785 ;
      END
   END dout0[478]
   PIN dout0[479]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  500.8075 115.65 500.9425 115.785 ;
      END
   END dout0[479]
   PIN dout0[480]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.5125 115.65 501.6475 115.785 ;
      END
   END dout0[480]
   PIN dout0[481]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  502.2175 115.65 502.3525 115.785 ;
      END
   END dout0[481]
   PIN dout0[482]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  502.9225 115.65 503.0575 115.785 ;
      END
   END dout0[482]
   PIN dout0[483]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  503.6275 115.65 503.7625 115.785 ;
      END
   END dout0[483]
   PIN dout0[484]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.3325 115.65 504.4675 115.785 ;
      END
   END dout0[484]
   PIN dout0[485]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  505.0375 115.65 505.1725 115.785 ;
      END
   END dout0[485]
   PIN dout0[486]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  505.7425 115.65 505.8775 115.785 ;
      END
   END dout0[486]
   PIN dout0[487]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  506.4475 115.65 506.5825 115.785 ;
      END
   END dout0[487]
   PIN dout0[488]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.1525 115.65 507.2875 115.785 ;
      END
   END dout0[488]
   PIN dout0[489]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.8575 115.65 507.9925 115.785 ;
      END
   END dout0[489]
   PIN dout0[490]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  508.5625 115.65 508.6975 115.785 ;
      END
   END dout0[490]
   PIN dout0[491]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.2675 115.65 509.4025 115.785 ;
      END
   END dout0[491]
   PIN dout0[492]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.9725 115.65 510.1075 115.785 ;
      END
   END dout0[492]
   PIN dout0[493]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.6775 115.65 510.8125 115.785 ;
      END
   END dout0[493]
   PIN dout0[494]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  511.3825 115.65 511.5175 115.785 ;
      END
   END dout0[494]
   PIN dout0[495]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.0875 115.65 512.2225 115.785 ;
      END
   END dout0[495]
   PIN dout0[496]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.7925 115.65 512.9275 115.785 ;
      END
   END dout0[496]
   PIN dout0[497]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  513.4975 115.65 513.6325 115.785 ;
      END
   END dout0[497]
   PIN dout0[498]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.2025 115.65 514.3375 115.785 ;
      END
   END dout0[498]
   PIN dout0[499]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.9075 115.65 515.0425 115.785 ;
      END
   END dout0[499]
   PIN dout0[500]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.6125 115.65 515.7475 115.785 ;
      END
   END dout0[500]
   PIN dout0[501]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  516.3175 115.65 516.4525 115.785 ;
      END
   END dout0[501]
   PIN dout0[502]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  517.0225 115.65 517.1575 115.785 ;
      END
   END dout0[502]
   PIN dout0[503]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  517.7275 115.65 517.8625 115.785 ;
      END
   END dout0[503]
   PIN dout0[504]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.4325 115.65 518.5675 115.785 ;
      END
   END dout0[504]
   PIN dout0[505]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  519.1375 115.65 519.2725 115.785 ;
      END
   END dout0[505]
   PIN dout0[506]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  519.8425 115.65 519.9775 115.785 ;
      END
   END dout0[506]
   PIN dout0[507]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  520.5475 115.65 520.6825 115.785 ;
      END
   END dout0[507]
   PIN dout0[508]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.2525 115.65 521.3875 115.785 ;
      END
   END dout0[508]
   PIN dout0[509]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.9575 115.65 522.0925 115.785 ;
      END
   END dout0[509]
   PIN dout0[510]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  522.6625 115.65 522.7975 115.785 ;
      END
   END dout0[510]
   PIN dout0[511]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  523.3675 115.65 523.5025 115.785 ;
      END
   END dout0[511]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  1591.52 1.4 1592.22 217.42 ;
         LAYER metal3 ;
         RECT  1.4 1.4 1592.22 2.1 ;
         LAYER metal3 ;
         RECT  1.4 216.72 1592.22 217.42 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 217.42 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 0.0 1593.62 0.7 ;
         LAYER metal4 ;
         RECT  1592.92 0.0 1593.62 218.82 ;
         LAYER metal3 ;
         RECT  0.0 218.12 1593.62 218.82 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 218.82 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 1593.48 218.68 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 1593.48 218.68 ;
   LAYER  metal3 ;
      RECT  0.14 4.0975 126.205 4.5125 ;
      RECT  126.62 4.0975 129.065 4.5125 ;
      RECT  129.48 4.0975 131.925 4.5125 ;
      RECT  132.34 4.0975 134.785 4.5125 ;
      RECT  135.2 4.0975 137.645 4.5125 ;
      RECT  138.06 4.0975 140.505 4.5125 ;
      RECT  140.92 4.0975 143.365 4.5125 ;
      RECT  143.78 4.0975 146.225 4.5125 ;
      RECT  146.64 4.0975 149.085 4.5125 ;
      RECT  149.5 4.0975 151.945 4.5125 ;
      RECT  152.36 4.0975 154.805 4.5125 ;
      RECT  155.22 4.0975 157.665 4.5125 ;
      RECT  158.08 4.0975 160.525 4.5125 ;
      RECT  160.94 4.0975 163.385 4.5125 ;
      RECT  163.8 4.0975 166.245 4.5125 ;
      RECT  166.66 4.0975 169.105 4.5125 ;
      RECT  169.52 4.0975 171.965 4.5125 ;
      RECT  172.38 4.0975 174.825 4.5125 ;
      RECT  175.24 4.0975 177.685 4.5125 ;
      RECT  178.1 4.0975 180.545 4.5125 ;
      RECT  180.96 4.0975 183.405 4.5125 ;
      RECT  183.82 4.0975 186.265 4.5125 ;
      RECT  186.68 4.0975 189.125 4.5125 ;
      RECT  189.54 4.0975 191.985 4.5125 ;
      RECT  192.4 4.0975 194.845 4.5125 ;
      RECT  195.26 4.0975 197.705 4.5125 ;
      RECT  198.12 4.0975 200.565 4.5125 ;
      RECT  200.98 4.0975 203.425 4.5125 ;
      RECT  203.84 4.0975 206.285 4.5125 ;
      RECT  206.7 4.0975 209.145 4.5125 ;
      RECT  209.56 4.0975 212.005 4.5125 ;
      RECT  212.42 4.0975 214.865 4.5125 ;
      RECT  215.28 4.0975 217.725 4.5125 ;
      RECT  218.14 4.0975 220.585 4.5125 ;
      RECT  221.0 4.0975 223.445 4.5125 ;
      RECT  223.86 4.0975 226.305 4.5125 ;
      RECT  226.72 4.0975 229.165 4.5125 ;
      RECT  229.58 4.0975 232.025 4.5125 ;
      RECT  232.44 4.0975 234.885 4.5125 ;
      RECT  235.3 4.0975 237.745 4.5125 ;
      RECT  238.16 4.0975 240.605 4.5125 ;
      RECT  241.02 4.0975 243.465 4.5125 ;
      RECT  243.88 4.0975 246.325 4.5125 ;
      RECT  246.74 4.0975 249.185 4.5125 ;
      RECT  249.6 4.0975 252.045 4.5125 ;
      RECT  252.46 4.0975 254.905 4.5125 ;
      RECT  255.32 4.0975 257.765 4.5125 ;
      RECT  258.18 4.0975 260.625 4.5125 ;
      RECT  261.04 4.0975 263.485 4.5125 ;
      RECT  263.9 4.0975 266.345 4.5125 ;
      RECT  266.76 4.0975 269.205 4.5125 ;
      RECT  269.62 4.0975 272.065 4.5125 ;
      RECT  272.48 4.0975 274.925 4.5125 ;
      RECT  275.34 4.0975 277.785 4.5125 ;
      RECT  278.2 4.0975 280.645 4.5125 ;
      RECT  281.06 4.0975 283.505 4.5125 ;
      RECT  283.92 4.0975 286.365 4.5125 ;
      RECT  286.78 4.0975 289.225 4.5125 ;
      RECT  289.64 4.0975 292.085 4.5125 ;
      RECT  292.5 4.0975 294.945 4.5125 ;
      RECT  295.36 4.0975 297.805 4.5125 ;
      RECT  298.22 4.0975 300.665 4.5125 ;
      RECT  301.08 4.0975 303.525 4.5125 ;
      RECT  303.94 4.0975 306.385 4.5125 ;
      RECT  306.8 4.0975 309.245 4.5125 ;
      RECT  309.66 4.0975 312.105 4.5125 ;
      RECT  312.52 4.0975 314.965 4.5125 ;
      RECT  315.38 4.0975 317.825 4.5125 ;
      RECT  318.24 4.0975 320.685 4.5125 ;
      RECT  321.1 4.0975 323.545 4.5125 ;
      RECT  323.96 4.0975 326.405 4.5125 ;
      RECT  326.82 4.0975 329.265 4.5125 ;
      RECT  329.68 4.0975 332.125 4.5125 ;
      RECT  332.54 4.0975 334.985 4.5125 ;
      RECT  335.4 4.0975 337.845 4.5125 ;
      RECT  338.26 4.0975 340.705 4.5125 ;
      RECT  341.12 4.0975 343.565 4.5125 ;
      RECT  343.98 4.0975 346.425 4.5125 ;
      RECT  346.84 4.0975 349.285 4.5125 ;
      RECT  349.7 4.0975 352.145 4.5125 ;
      RECT  352.56 4.0975 355.005 4.5125 ;
      RECT  355.42 4.0975 357.865 4.5125 ;
      RECT  358.28 4.0975 360.725 4.5125 ;
      RECT  361.14 4.0975 363.585 4.5125 ;
      RECT  364.0 4.0975 366.445 4.5125 ;
      RECT  366.86 4.0975 369.305 4.5125 ;
      RECT  369.72 4.0975 372.165 4.5125 ;
      RECT  372.58 4.0975 375.025 4.5125 ;
      RECT  375.44 4.0975 377.885 4.5125 ;
      RECT  378.3 4.0975 380.745 4.5125 ;
      RECT  381.16 4.0975 383.605 4.5125 ;
      RECT  384.02 4.0975 386.465 4.5125 ;
      RECT  386.88 4.0975 389.325 4.5125 ;
      RECT  389.74 4.0975 392.185 4.5125 ;
      RECT  392.6 4.0975 395.045 4.5125 ;
      RECT  395.46 4.0975 397.905 4.5125 ;
      RECT  398.32 4.0975 400.765 4.5125 ;
      RECT  401.18 4.0975 403.625 4.5125 ;
      RECT  404.04 4.0975 406.485 4.5125 ;
      RECT  406.9 4.0975 409.345 4.5125 ;
      RECT  409.76 4.0975 412.205 4.5125 ;
      RECT  412.62 4.0975 415.065 4.5125 ;
      RECT  415.48 4.0975 417.925 4.5125 ;
      RECT  418.34 4.0975 420.785 4.5125 ;
      RECT  421.2 4.0975 423.645 4.5125 ;
      RECT  424.06 4.0975 426.505 4.5125 ;
      RECT  426.92 4.0975 429.365 4.5125 ;
      RECT  429.78 4.0975 432.225 4.5125 ;
      RECT  432.64 4.0975 435.085 4.5125 ;
      RECT  435.5 4.0975 437.945 4.5125 ;
      RECT  438.36 4.0975 440.805 4.5125 ;
      RECT  441.22 4.0975 443.665 4.5125 ;
      RECT  444.08 4.0975 446.525 4.5125 ;
      RECT  446.94 4.0975 449.385 4.5125 ;
      RECT  449.8 4.0975 452.245 4.5125 ;
      RECT  452.66 4.0975 455.105 4.5125 ;
      RECT  455.52 4.0975 457.965 4.5125 ;
      RECT  458.38 4.0975 460.825 4.5125 ;
      RECT  461.24 4.0975 463.685 4.5125 ;
      RECT  464.1 4.0975 466.545 4.5125 ;
      RECT  466.96 4.0975 469.405 4.5125 ;
      RECT  469.82 4.0975 472.265 4.5125 ;
      RECT  472.68 4.0975 475.125 4.5125 ;
      RECT  475.54 4.0975 477.985 4.5125 ;
      RECT  478.4 4.0975 480.845 4.5125 ;
      RECT  481.26 4.0975 483.705 4.5125 ;
      RECT  484.12 4.0975 486.565 4.5125 ;
      RECT  486.98 4.0975 489.425 4.5125 ;
      RECT  489.84 4.0975 492.285 4.5125 ;
      RECT  492.7 4.0975 495.145 4.5125 ;
      RECT  495.56 4.0975 498.005 4.5125 ;
      RECT  498.42 4.0975 500.865 4.5125 ;
      RECT  501.28 4.0975 503.725 4.5125 ;
      RECT  504.14 4.0975 506.585 4.5125 ;
      RECT  507.0 4.0975 509.445 4.5125 ;
      RECT  509.86 4.0975 512.305 4.5125 ;
      RECT  512.72 4.0975 515.165 4.5125 ;
      RECT  515.58 4.0975 518.025 4.5125 ;
      RECT  518.44 4.0975 520.885 4.5125 ;
      RECT  521.3 4.0975 523.745 4.5125 ;
      RECT  524.16 4.0975 526.605 4.5125 ;
      RECT  527.02 4.0975 529.465 4.5125 ;
      RECT  529.88 4.0975 532.325 4.5125 ;
      RECT  532.74 4.0975 535.185 4.5125 ;
      RECT  535.6 4.0975 538.045 4.5125 ;
      RECT  538.46 4.0975 540.905 4.5125 ;
      RECT  541.32 4.0975 543.765 4.5125 ;
      RECT  544.18 4.0975 546.625 4.5125 ;
      RECT  547.04 4.0975 549.485 4.5125 ;
      RECT  549.9 4.0975 552.345 4.5125 ;
      RECT  552.76 4.0975 555.205 4.5125 ;
      RECT  555.62 4.0975 558.065 4.5125 ;
      RECT  558.48 4.0975 560.925 4.5125 ;
      RECT  561.34 4.0975 563.785 4.5125 ;
      RECT  564.2 4.0975 566.645 4.5125 ;
      RECT  567.06 4.0975 569.505 4.5125 ;
      RECT  569.92 4.0975 572.365 4.5125 ;
      RECT  572.78 4.0975 575.225 4.5125 ;
      RECT  575.64 4.0975 578.085 4.5125 ;
      RECT  578.5 4.0975 580.945 4.5125 ;
      RECT  581.36 4.0975 583.805 4.5125 ;
      RECT  584.22 4.0975 586.665 4.5125 ;
      RECT  587.08 4.0975 589.525 4.5125 ;
      RECT  589.94 4.0975 592.385 4.5125 ;
      RECT  592.8 4.0975 595.245 4.5125 ;
      RECT  595.66 4.0975 598.105 4.5125 ;
      RECT  598.52 4.0975 600.965 4.5125 ;
      RECT  601.38 4.0975 603.825 4.5125 ;
      RECT  604.24 4.0975 606.685 4.5125 ;
      RECT  607.1 4.0975 609.545 4.5125 ;
      RECT  609.96 4.0975 612.405 4.5125 ;
      RECT  612.82 4.0975 615.265 4.5125 ;
      RECT  615.68 4.0975 618.125 4.5125 ;
      RECT  618.54 4.0975 620.985 4.5125 ;
      RECT  621.4 4.0975 623.845 4.5125 ;
      RECT  624.26 4.0975 626.705 4.5125 ;
      RECT  627.12 4.0975 629.565 4.5125 ;
      RECT  629.98 4.0975 632.425 4.5125 ;
      RECT  632.84 4.0975 635.285 4.5125 ;
      RECT  635.7 4.0975 638.145 4.5125 ;
      RECT  638.56 4.0975 641.005 4.5125 ;
      RECT  641.42 4.0975 643.865 4.5125 ;
      RECT  644.28 4.0975 646.725 4.5125 ;
      RECT  647.14 4.0975 649.585 4.5125 ;
      RECT  650.0 4.0975 652.445 4.5125 ;
      RECT  652.86 4.0975 655.305 4.5125 ;
      RECT  655.72 4.0975 658.165 4.5125 ;
      RECT  658.58 4.0975 661.025 4.5125 ;
      RECT  661.44 4.0975 663.885 4.5125 ;
      RECT  664.3 4.0975 666.745 4.5125 ;
      RECT  667.16 4.0975 669.605 4.5125 ;
      RECT  670.02 4.0975 672.465 4.5125 ;
      RECT  672.88 4.0975 675.325 4.5125 ;
      RECT  675.74 4.0975 678.185 4.5125 ;
      RECT  678.6 4.0975 681.045 4.5125 ;
      RECT  681.46 4.0975 683.905 4.5125 ;
      RECT  684.32 4.0975 686.765 4.5125 ;
      RECT  687.18 4.0975 689.625 4.5125 ;
      RECT  690.04 4.0975 692.485 4.5125 ;
      RECT  692.9 4.0975 695.345 4.5125 ;
      RECT  695.76 4.0975 698.205 4.5125 ;
      RECT  698.62 4.0975 701.065 4.5125 ;
      RECT  701.48 4.0975 703.925 4.5125 ;
      RECT  704.34 4.0975 706.785 4.5125 ;
      RECT  707.2 4.0975 709.645 4.5125 ;
      RECT  710.06 4.0975 712.505 4.5125 ;
      RECT  712.92 4.0975 715.365 4.5125 ;
      RECT  715.78 4.0975 718.225 4.5125 ;
      RECT  718.64 4.0975 721.085 4.5125 ;
      RECT  721.5 4.0975 723.945 4.5125 ;
      RECT  724.36 4.0975 726.805 4.5125 ;
      RECT  727.22 4.0975 729.665 4.5125 ;
      RECT  730.08 4.0975 732.525 4.5125 ;
      RECT  732.94 4.0975 735.385 4.5125 ;
      RECT  735.8 4.0975 738.245 4.5125 ;
      RECT  738.66 4.0975 741.105 4.5125 ;
      RECT  741.52 4.0975 743.965 4.5125 ;
      RECT  744.38 4.0975 746.825 4.5125 ;
      RECT  747.24 4.0975 749.685 4.5125 ;
      RECT  750.1 4.0975 752.545 4.5125 ;
      RECT  752.96 4.0975 755.405 4.5125 ;
      RECT  755.82 4.0975 758.265 4.5125 ;
      RECT  758.68 4.0975 761.125 4.5125 ;
      RECT  761.54 4.0975 763.985 4.5125 ;
      RECT  764.4 4.0975 766.845 4.5125 ;
      RECT  767.26 4.0975 769.705 4.5125 ;
      RECT  770.12 4.0975 772.565 4.5125 ;
      RECT  772.98 4.0975 775.425 4.5125 ;
      RECT  775.84 4.0975 778.285 4.5125 ;
      RECT  778.7 4.0975 781.145 4.5125 ;
      RECT  781.56 4.0975 784.005 4.5125 ;
      RECT  784.42 4.0975 786.865 4.5125 ;
      RECT  787.28 4.0975 789.725 4.5125 ;
      RECT  790.14 4.0975 792.585 4.5125 ;
      RECT  793.0 4.0975 795.445 4.5125 ;
      RECT  795.86 4.0975 798.305 4.5125 ;
      RECT  798.72 4.0975 801.165 4.5125 ;
      RECT  801.58 4.0975 804.025 4.5125 ;
      RECT  804.44 4.0975 806.885 4.5125 ;
      RECT  807.3 4.0975 809.745 4.5125 ;
      RECT  810.16 4.0975 812.605 4.5125 ;
      RECT  813.02 4.0975 815.465 4.5125 ;
      RECT  815.88 4.0975 818.325 4.5125 ;
      RECT  818.74 4.0975 821.185 4.5125 ;
      RECT  821.6 4.0975 824.045 4.5125 ;
      RECT  824.46 4.0975 826.905 4.5125 ;
      RECT  827.32 4.0975 829.765 4.5125 ;
      RECT  830.18 4.0975 832.625 4.5125 ;
      RECT  833.04 4.0975 835.485 4.5125 ;
      RECT  835.9 4.0975 838.345 4.5125 ;
      RECT  838.76 4.0975 841.205 4.5125 ;
      RECT  841.62 4.0975 844.065 4.5125 ;
      RECT  844.48 4.0975 846.925 4.5125 ;
      RECT  847.34 4.0975 849.785 4.5125 ;
      RECT  850.2 4.0975 852.645 4.5125 ;
      RECT  853.06 4.0975 855.505 4.5125 ;
      RECT  855.92 4.0975 858.365 4.5125 ;
      RECT  858.78 4.0975 861.225 4.5125 ;
      RECT  861.64 4.0975 864.085 4.5125 ;
      RECT  864.5 4.0975 866.945 4.5125 ;
      RECT  867.36 4.0975 869.805 4.5125 ;
      RECT  870.22 4.0975 872.665 4.5125 ;
      RECT  873.08 4.0975 875.525 4.5125 ;
      RECT  875.94 4.0975 878.385 4.5125 ;
      RECT  878.8 4.0975 881.245 4.5125 ;
      RECT  881.66 4.0975 884.105 4.5125 ;
      RECT  884.52 4.0975 886.965 4.5125 ;
      RECT  887.38 4.0975 889.825 4.5125 ;
      RECT  890.24 4.0975 892.685 4.5125 ;
      RECT  893.1 4.0975 895.545 4.5125 ;
      RECT  895.96 4.0975 898.405 4.5125 ;
      RECT  898.82 4.0975 901.265 4.5125 ;
      RECT  901.68 4.0975 904.125 4.5125 ;
      RECT  904.54 4.0975 906.985 4.5125 ;
      RECT  907.4 4.0975 909.845 4.5125 ;
      RECT  910.26 4.0975 912.705 4.5125 ;
      RECT  913.12 4.0975 915.565 4.5125 ;
      RECT  915.98 4.0975 918.425 4.5125 ;
      RECT  918.84 4.0975 921.285 4.5125 ;
      RECT  921.7 4.0975 924.145 4.5125 ;
      RECT  924.56 4.0975 927.005 4.5125 ;
      RECT  927.42 4.0975 929.865 4.5125 ;
      RECT  930.28 4.0975 932.725 4.5125 ;
      RECT  933.14 4.0975 935.585 4.5125 ;
      RECT  936.0 4.0975 938.445 4.5125 ;
      RECT  938.86 4.0975 941.305 4.5125 ;
      RECT  941.72 4.0975 944.165 4.5125 ;
      RECT  944.58 4.0975 947.025 4.5125 ;
      RECT  947.44 4.0975 949.885 4.5125 ;
      RECT  950.3 4.0975 952.745 4.5125 ;
      RECT  953.16 4.0975 955.605 4.5125 ;
      RECT  956.02 4.0975 958.465 4.5125 ;
      RECT  958.88 4.0975 961.325 4.5125 ;
      RECT  961.74 4.0975 964.185 4.5125 ;
      RECT  964.6 4.0975 967.045 4.5125 ;
      RECT  967.46 4.0975 969.905 4.5125 ;
      RECT  970.32 4.0975 972.765 4.5125 ;
      RECT  973.18 4.0975 975.625 4.5125 ;
      RECT  976.04 4.0975 978.485 4.5125 ;
      RECT  978.9 4.0975 981.345 4.5125 ;
      RECT  981.76 4.0975 984.205 4.5125 ;
      RECT  984.62 4.0975 987.065 4.5125 ;
      RECT  987.48 4.0975 989.925 4.5125 ;
      RECT  990.34 4.0975 992.785 4.5125 ;
      RECT  993.2 4.0975 995.645 4.5125 ;
      RECT  996.06 4.0975 998.505 4.5125 ;
      RECT  998.92 4.0975 1001.365 4.5125 ;
      RECT  1001.78 4.0975 1004.225 4.5125 ;
      RECT  1004.64 4.0975 1007.085 4.5125 ;
      RECT  1007.5 4.0975 1009.945 4.5125 ;
      RECT  1010.36 4.0975 1012.805 4.5125 ;
      RECT  1013.22 4.0975 1015.665 4.5125 ;
      RECT  1016.08 4.0975 1018.525 4.5125 ;
      RECT  1018.94 4.0975 1021.385 4.5125 ;
      RECT  1021.8 4.0975 1024.245 4.5125 ;
      RECT  1024.66 4.0975 1027.105 4.5125 ;
      RECT  1027.52 4.0975 1029.965 4.5125 ;
      RECT  1030.38 4.0975 1032.825 4.5125 ;
      RECT  1033.24 4.0975 1035.685 4.5125 ;
      RECT  1036.1 4.0975 1038.545 4.5125 ;
      RECT  1038.96 4.0975 1041.405 4.5125 ;
      RECT  1041.82 4.0975 1044.265 4.5125 ;
      RECT  1044.68 4.0975 1047.125 4.5125 ;
      RECT  1047.54 4.0975 1049.985 4.5125 ;
      RECT  1050.4 4.0975 1052.845 4.5125 ;
      RECT  1053.26 4.0975 1055.705 4.5125 ;
      RECT  1056.12 4.0975 1058.565 4.5125 ;
      RECT  1058.98 4.0975 1061.425 4.5125 ;
      RECT  1061.84 4.0975 1064.285 4.5125 ;
      RECT  1064.7 4.0975 1067.145 4.5125 ;
      RECT  1067.56 4.0975 1070.005 4.5125 ;
      RECT  1070.42 4.0975 1072.865 4.5125 ;
      RECT  1073.28 4.0975 1075.725 4.5125 ;
      RECT  1076.14 4.0975 1078.585 4.5125 ;
      RECT  1079.0 4.0975 1081.445 4.5125 ;
      RECT  1081.86 4.0975 1084.305 4.5125 ;
      RECT  1084.72 4.0975 1087.165 4.5125 ;
      RECT  1087.58 4.0975 1090.025 4.5125 ;
      RECT  1090.44 4.0975 1092.885 4.5125 ;
      RECT  1093.3 4.0975 1095.745 4.5125 ;
      RECT  1096.16 4.0975 1098.605 4.5125 ;
      RECT  1099.02 4.0975 1101.465 4.5125 ;
      RECT  1101.88 4.0975 1104.325 4.5125 ;
      RECT  1104.74 4.0975 1107.185 4.5125 ;
      RECT  1107.6 4.0975 1110.045 4.5125 ;
      RECT  1110.46 4.0975 1112.905 4.5125 ;
      RECT  1113.32 4.0975 1115.765 4.5125 ;
      RECT  1116.18 4.0975 1118.625 4.5125 ;
      RECT  1119.04 4.0975 1121.485 4.5125 ;
      RECT  1121.9 4.0975 1124.345 4.5125 ;
      RECT  1124.76 4.0975 1127.205 4.5125 ;
      RECT  1127.62 4.0975 1130.065 4.5125 ;
      RECT  1130.48 4.0975 1132.925 4.5125 ;
      RECT  1133.34 4.0975 1135.785 4.5125 ;
      RECT  1136.2 4.0975 1138.645 4.5125 ;
      RECT  1139.06 4.0975 1141.505 4.5125 ;
      RECT  1141.92 4.0975 1144.365 4.5125 ;
      RECT  1144.78 4.0975 1147.225 4.5125 ;
      RECT  1147.64 4.0975 1150.085 4.5125 ;
      RECT  1150.5 4.0975 1152.945 4.5125 ;
      RECT  1153.36 4.0975 1155.805 4.5125 ;
      RECT  1156.22 4.0975 1158.665 4.5125 ;
      RECT  1159.08 4.0975 1161.525 4.5125 ;
      RECT  1161.94 4.0975 1164.385 4.5125 ;
      RECT  1164.8 4.0975 1167.245 4.5125 ;
      RECT  1167.66 4.0975 1170.105 4.5125 ;
      RECT  1170.52 4.0975 1172.965 4.5125 ;
      RECT  1173.38 4.0975 1175.825 4.5125 ;
      RECT  1176.24 4.0975 1178.685 4.5125 ;
      RECT  1179.1 4.0975 1181.545 4.5125 ;
      RECT  1181.96 4.0975 1184.405 4.5125 ;
      RECT  1184.82 4.0975 1187.265 4.5125 ;
      RECT  1187.68 4.0975 1190.125 4.5125 ;
      RECT  1190.54 4.0975 1192.985 4.5125 ;
      RECT  1193.4 4.0975 1195.845 4.5125 ;
      RECT  1196.26 4.0975 1198.705 4.5125 ;
      RECT  1199.12 4.0975 1201.565 4.5125 ;
      RECT  1201.98 4.0975 1204.425 4.5125 ;
      RECT  1204.84 4.0975 1207.285 4.5125 ;
      RECT  1207.7 4.0975 1210.145 4.5125 ;
      RECT  1210.56 4.0975 1213.005 4.5125 ;
      RECT  1213.42 4.0975 1215.865 4.5125 ;
      RECT  1216.28 4.0975 1218.725 4.5125 ;
      RECT  1219.14 4.0975 1221.585 4.5125 ;
      RECT  1222.0 4.0975 1224.445 4.5125 ;
      RECT  1224.86 4.0975 1227.305 4.5125 ;
      RECT  1227.72 4.0975 1230.165 4.5125 ;
      RECT  1230.58 4.0975 1233.025 4.5125 ;
      RECT  1233.44 4.0975 1235.885 4.5125 ;
      RECT  1236.3 4.0975 1238.745 4.5125 ;
      RECT  1239.16 4.0975 1241.605 4.5125 ;
      RECT  1242.02 4.0975 1244.465 4.5125 ;
      RECT  1244.88 4.0975 1247.325 4.5125 ;
      RECT  1247.74 4.0975 1250.185 4.5125 ;
      RECT  1250.6 4.0975 1253.045 4.5125 ;
      RECT  1253.46 4.0975 1255.905 4.5125 ;
      RECT  1256.32 4.0975 1258.765 4.5125 ;
      RECT  1259.18 4.0975 1261.625 4.5125 ;
      RECT  1262.04 4.0975 1264.485 4.5125 ;
      RECT  1264.9 4.0975 1267.345 4.5125 ;
      RECT  1267.76 4.0975 1270.205 4.5125 ;
      RECT  1270.62 4.0975 1273.065 4.5125 ;
      RECT  1273.48 4.0975 1275.925 4.5125 ;
      RECT  1276.34 4.0975 1278.785 4.5125 ;
      RECT  1279.2 4.0975 1281.645 4.5125 ;
      RECT  1282.06 4.0975 1284.505 4.5125 ;
      RECT  1284.92 4.0975 1287.365 4.5125 ;
      RECT  1287.78 4.0975 1290.225 4.5125 ;
      RECT  1290.64 4.0975 1293.085 4.5125 ;
      RECT  1293.5 4.0975 1295.945 4.5125 ;
      RECT  1296.36 4.0975 1298.805 4.5125 ;
      RECT  1299.22 4.0975 1301.665 4.5125 ;
      RECT  1302.08 4.0975 1304.525 4.5125 ;
      RECT  1304.94 4.0975 1307.385 4.5125 ;
      RECT  1307.8 4.0975 1310.245 4.5125 ;
      RECT  1310.66 4.0975 1313.105 4.5125 ;
      RECT  1313.52 4.0975 1315.965 4.5125 ;
      RECT  1316.38 4.0975 1318.825 4.5125 ;
      RECT  1319.24 4.0975 1321.685 4.5125 ;
      RECT  1322.1 4.0975 1324.545 4.5125 ;
      RECT  1324.96 4.0975 1327.405 4.5125 ;
      RECT  1327.82 4.0975 1330.265 4.5125 ;
      RECT  1330.68 4.0975 1333.125 4.5125 ;
      RECT  1333.54 4.0975 1335.985 4.5125 ;
      RECT  1336.4 4.0975 1338.845 4.5125 ;
      RECT  1339.26 4.0975 1341.705 4.5125 ;
      RECT  1342.12 4.0975 1344.565 4.5125 ;
      RECT  1344.98 4.0975 1347.425 4.5125 ;
      RECT  1347.84 4.0975 1350.285 4.5125 ;
      RECT  1350.7 4.0975 1353.145 4.5125 ;
      RECT  1353.56 4.0975 1356.005 4.5125 ;
      RECT  1356.42 4.0975 1358.865 4.5125 ;
      RECT  1359.28 4.0975 1361.725 4.5125 ;
      RECT  1362.14 4.0975 1364.585 4.5125 ;
      RECT  1365.0 4.0975 1367.445 4.5125 ;
      RECT  1367.86 4.0975 1370.305 4.5125 ;
      RECT  1370.72 4.0975 1373.165 4.5125 ;
      RECT  1373.58 4.0975 1376.025 4.5125 ;
      RECT  1376.44 4.0975 1378.885 4.5125 ;
      RECT  1379.3 4.0975 1381.745 4.5125 ;
      RECT  1382.16 4.0975 1384.605 4.5125 ;
      RECT  1385.02 4.0975 1387.465 4.5125 ;
      RECT  1387.88 4.0975 1390.325 4.5125 ;
      RECT  1390.74 4.0975 1393.185 4.5125 ;
      RECT  1393.6 4.0975 1396.045 4.5125 ;
      RECT  1396.46 4.0975 1398.905 4.5125 ;
      RECT  1399.32 4.0975 1401.765 4.5125 ;
      RECT  1402.18 4.0975 1404.625 4.5125 ;
      RECT  1405.04 4.0975 1407.485 4.5125 ;
      RECT  1407.9 4.0975 1410.345 4.5125 ;
      RECT  1410.76 4.0975 1413.205 4.5125 ;
      RECT  1413.62 4.0975 1416.065 4.5125 ;
      RECT  1416.48 4.0975 1418.925 4.5125 ;
      RECT  1419.34 4.0975 1421.785 4.5125 ;
      RECT  1422.2 4.0975 1424.645 4.5125 ;
      RECT  1425.06 4.0975 1427.505 4.5125 ;
      RECT  1427.92 4.0975 1430.365 4.5125 ;
      RECT  1430.78 4.0975 1433.225 4.5125 ;
      RECT  1433.64 4.0975 1436.085 4.5125 ;
      RECT  1436.5 4.0975 1438.945 4.5125 ;
      RECT  1439.36 4.0975 1441.805 4.5125 ;
      RECT  1442.22 4.0975 1444.665 4.5125 ;
      RECT  1445.08 4.0975 1447.525 4.5125 ;
      RECT  1447.94 4.0975 1450.385 4.5125 ;
      RECT  1450.8 4.0975 1453.245 4.5125 ;
      RECT  1453.66 4.0975 1456.105 4.5125 ;
      RECT  1456.52 4.0975 1458.965 4.5125 ;
      RECT  1459.38 4.0975 1461.825 4.5125 ;
      RECT  1462.24 4.0975 1464.685 4.5125 ;
      RECT  1465.1 4.0975 1467.545 4.5125 ;
      RECT  1467.96 4.0975 1470.405 4.5125 ;
      RECT  1470.82 4.0975 1473.265 4.5125 ;
      RECT  1473.68 4.0975 1476.125 4.5125 ;
      RECT  1476.54 4.0975 1478.985 4.5125 ;
      RECT  1479.4 4.0975 1481.845 4.5125 ;
      RECT  1482.26 4.0975 1484.705 4.5125 ;
      RECT  1485.12 4.0975 1487.565 4.5125 ;
      RECT  1487.98 4.0975 1490.425 4.5125 ;
      RECT  1490.84 4.0975 1493.285 4.5125 ;
      RECT  1493.7 4.0975 1496.145 4.5125 ;
      RECT  1496.56 4.0975 1499.005 4.5125 ;
      RECT  1499.42 4.0975 1501.865 4.5125 ;
      RECT  1502.28 4.0975 1504.725 4.5125 ;
      RECT  1505.14 4.0975 1507.585 4.5125 ;
      RECT  1508.0 4.0975 1510.445 4.5125 ;
      RECT  1510.86 4.0975 1513.305 4.5125 ;
      RECT  1513.72 4.0975 1516.165 4.5125 ;
      RECT  1516.58 4.0975 1519.025 4.5125 ;
      RECT  1519.44 4.0975 1521.885 4.5125 ;
      RECT  1522.3 4.0975 1524.745 4.5125 ;
      RECT  1525.16 4.0975 1527.605 4.5125 ;
      RECT  1528.02 4.0975 1530.465 4.5125 ;
      RECT  1530.88 4.0975 1533.325 4.5125 ;
      RECT  1533.74 4.0975 1536.185 4.5125 ;
      RECT  1536.6 4.0975 1539.045 4.5125 ;
      RECT  1539.46 4.0975 1541.905 4.5125 ;
      RECT  1542.32 4.0975 1544.765 4.5125 ;
      RECT  1545.18 4.0975 1547.625 4.5125 ;
      RECT  1548.04 4.0975 1550.485 4.5125 ;
      RECT  1550.9 4.0975 1553.345 4.5125 ;
      RECT  1553.76 4.0975 1556.205 4.5125 ;
      RECT  1556.62 4.0975 1559.065 4.5125 ;
      RECT  1559.48 4.0975 1561.925 4.5125 ;
      RECT  1562.34 4.0975 1564.785 4.5125 ;
      RECT  1565.2 4.0975 1567.645 4.5125 ;
      RECT  1568.06 4.0975 1570.505 4.5125 ;
      RECT  1570.92 4.0975 1573.365 4.5125 ;
      RECT  1573.78 4.0975 1576.225 4.5125 ;
      RECT  1576.64 4.0975 1579.085 4.5125 ;
      RECT  1579.5 4.0975 1581.945 4.5125 ;
      RECT  1582.36 4.0975 1584.805 4.5125 ;
      RECT  1585.22 4.0975 1587.665 4.5125 ;
      RECT  1588.08 4.0975 1593.48 4.5125 ;
      RECT  0.14 148.5825 120.485 148.9975 ;
      RECT  120.485 4.5125 120.9 148.5825 ;
      RECT  120.9 4.5125 126.205 148.5825 ;
      RECT  120.9 148.5825 126.205 148.9975 ;
      RECT  120.485 148.9975 120.9 151.3125 ;
      RECT  120.485 151.7275 120.9 153.5225 ;
      RECT  120.485 153.9375 120.9 156.2525 ;
      RECT  120.485 156.6675 120.9 158.4625 ;
      RECT  120.485 158.8775 120.9 161.1925 ;
      RECT  0.14 4.5125 3.245 103.8625 ;
      RECT  0.14 103.8625 3.245 104.2775 ;
      RECT  0.14 104.2775 3.245 148.5825 ;
      RECT  3.245 4.5125 3.66 103.8625 ;
      RECT  3.66 4.5125 120.485 103.8625 ;
      RECT  3.245 104.2775 3.66 106.5925 ;
      RECT  3.245 107.0075 3.66 148.5825 ;
      RECT  3.66 103.8625 9.4875 103.9475 ;
      RECT  3.66 103.9475 9.4875 104.2775 ;
      RECT  9.4875 103.8625 9.9025 103.9475 ;
      RECT  9.9025 103.8625 120.485 103.9475 ;
      RECT  9.9025 103.9475 120.485 104.2775 ;
      RECT  3.66 104.2775 9.4875 104.3625 ;
      RECT  3.66 104.3625 9.4875 148.5825 ;
      RECT  9.4875 104.3625 9.9025 148.5825 ;
      RECT  9.9025 104.2775 120.485 104.3625 ;
      RECT  9.9025 104.3625 120.485 148.5825 ;
      RECT  126.62 4.5125 162.9725 115.51 ;
      RECT  126.62 115.51 162.9725 115.925 ;
      RECT  162.9725 4.5125 163.3875 115.51 ;
      RECT  163.3875 4.5125 1593.48 115.51 ;
      RECT  163.3875 115.51 163.6775 115.925 ;
      RECT  164.0925 115.51 164.3825 115.925 ;
      RECT  164.7975 115.51 165.0875 115.925 ;
      RECT  165.5025 115.51 165.7925 115.925 ;
      RECT  166.2075 115.51 166.4975 115.925 ;
      RECT  166.9125 115.51 167.2025 115.925 ;
      RECT  167.6175 115.51 167.9075 115.925 ;
      RECT  168.3225 115.51 168.6125 115.925 ;
      RECT  169.0275 115.51 169.3175 115.925 ;
      RECT  169.7325 115.51 170.0225 115.925 ;
      RECT  170.4375 115.51 170.7275 115.925 ;
      RECT  171.1425 115.51 171.4325 115.925 ;
      RECT  171.8475 115.51 172.1375 115.925 ;
      RECT  172.5525 115.51 172.8425 115.925 ;
      RECT  173.2575 115.51 173.5475 115.925 ;
      RECT  173.9625 115.51 174.2525 115.925 ;
      RECT  174.6675 115.51 174.9575 115.925 ;
      RECT  175.3725 115.51 175.6625 115.925 ;
      RECT  176.0775 115.51 176.3675 115.925 ;
      RECT  176.7825 115.51 177.0725 115.925 ;
      RECT  177.4875 115.51 177.7775 115.925 ;
      RECT  178.1925 115.51 178.4825 115.925 ;
      RECT  178.8975 115.51 179.1875 115.925 ;
      RECT  179.6025 115.51 179.8925 115.925 ;
      RECT  180.3075 115.51 180.5975 115.925 ;
      RECT  181.0125 115.51 181.3025 115.925 ;
      RECT  181.7175 115.51 182.0075 115.925 ;
      RECT  182.4225 115.51 182.7125 115.925 ;
      RECT  183.1275 115.51 183.4175 115.925 ;
      RECT  183.8325 115.51 184.1225 115.925 ;
      RECT  184.5375 115.51 184.8275 115.925 ;
      RECT  185.2425 115.51 185.5325 115.925 ;
      RECT  185.9475 115.51 186.2375 115.925 ;
      RECT  186.6525 115.51 186.9425 115.925 ;
      RECT  187.3575 115.51 187.6475 115.925 ;
      RECT  188.0625 115.51 188.3525 115.925 ;
      RECT  188.7675 115.51 189.0575 115.925 ;
      RECT  189.4725 115.51 189.7625 115.925 ;
      RECT  190.1775 115.51 190.4675 115.925 ;
      RECT  190.8825 115.51 191.1725 115.925 ;
      RECT  191.5875 115.51 191.8775 115.925 ;
      RECT  192.2925 115.51 192.5825 115.925 ;
      RECT  192.9975 115.51 193.2875 115.925 ;
      RECT  193.7025 115.51 193.9925 115.925 ;
      RECT  194.4075 115.51 194.6975 115.925 ;
      RECT  195.1125 115.51 195.4025 115.925 ;
      RECT  195.8175 115.51 196.1075 115.925 ;
      RECT  196.5225 115.51 196.8125 115.925 ;
      RECT  197.2275 115.51 197.5175 115.925 ;
      RECT  197.9325 115.51 198.2225 115.925 ;
      RECT  198.6375 115.51 198.9275 115.925 ;
      RECT  199.3425 115.51 199.6325 115.925 ;
      RECT  200.0475 115.51 200.3375 115.925 ;
      RECT  200.7525 115.51 201.0425 115.925 ;
      RECT  201.4575 115.51 201.7475 115.925 ;
      RECT  202.1625 115.51 202.4525 115.925 ;
      RECT  202.8675 115.51 203.1575 115.925 ;
      RECT  203.5725 115.51 203.8625 115.925 ;
      RECT  204.2775 115.51 204.5675 115.925 ;
      RECT  204.9825 115.51 205.2725 115.925 ;
      RECT  205.6875 115.51 205.9775 115.925 ;
      RECT  206.3925 115.51 206.6825 115.925 ;
      RECT  207.0975 115.51 207.3875 115.925 ;
      RECT  207.8025 115.51 208.0925 115.925 ;
      RECT  208.5075 115.51 208.7975 115.925 ;
      RECT  209.2125 115.51 209.5025 115.925 ;
      RECT  209.9175 115.51 210.2075 115.925 ;
      RECT  210.6225 115.51 210.9125 115.925 ;
      RECT  211.3275 115.51 211.6175 115.925 ;
      RECT  212.0325 115.51 212.3225 115.925 ;
      RECT  212.7375 115.51 213.0275 115.925 ;
      RECT  213.4425 115.51 213.7325 115.925 ;
      RECT  214.1475 115.51 214.4375 115.925 ;
      RECT  214.8525 115.51 215.1425 115.925 ;
      RECT  215.5575 115.51 215.8475 115.925 ;
      RECT  216.2625 115.51 216.5525 115.925 ;
      RECT  216.9675 115.51 217.2575 115.925 ;
      RECT  217.6725 115.51 217.9625 115.925 ;
      RECT  218.3775 115.51 218.6675 115.925 ;
      RECT  219.0825 115.51 219.3725 115.925 ;
      RECT  219.7875 115.51 220.0775 115.925 ;
      RECT  220.4925 115.51 220.7825 115.925 ;
      RECT  221.1975 115.51 221.4875 115.925 ;
      RECT  221.9025 115.51 222.1925 115.925 ;
      RECT  222.6075 115.51 222.8975 115.925 ;
      RECT  223.3125 115.51 223.6025 115.925 ;
      RECT  224.0175 115.51 224.3075 115.925 ;
      RECT  224.7225 115.51 225.0125 115.925 ;
      RECT  225.4275 115.51 225.7175 115.925 ;
      RECT  226.1325 115.51 226.4225 115.925 ;
      RECT  226.8375 115.51 227.1275 115.925 ;
      RECT  227.5425 115.51 227.8325 115.925 ;
      RECT  228.2475 115.51 228.5375 115.925 ;
      RECT  228.9525 115.51 229.2425 115.925 ;
      RECT  229.6575 115.51 229.9475 115.925 ;
      RECT  230.3625 115.51 230.6525 115.925 ;
      RECT  231.0675 115.51 231.3575 115.925 ;
      RECT  231.7725 115.51 232.0625 115.925 ;
      RECT  232.4775 115.51 232.7675 115.925 ;
      RECT  233.1825 115.51 233.4725 115.925 ;
      RECT  233.8875 115.51 234.1775 115.925 ;
      RECT  234.5925 115.51 234.8825 115.925 ;
      RECT  235.2975 115.51 235.5875 115.925 ;
      RECT  236.0025 115.51 236.2925 115.925 ;
      RECT  236.7075 115.51 236.9975 115.925 ;
      RECT  237.4125 115.51 237.7025 115.925 ;
      RECT  238.1175 115.51 238.4075 115.925 ;
      RECT  238.8225 115.51 239.1125 115.925 ;
      RECT  239.5275 115.51 239.8175 115.925 ;
      RECT  240.2325 115.51 240.5225 115.925 ;
      RECT  240.9375 115.51 241.2275 115.925 ;
      RECT  241.6425 115.51 241.9325 115.925 ;
      RECT  242.3475 115.51 242.6375 115.925 ;
      RECT  243.0525 115.51 243.3425 115.925 ;
      RECT  243.7575 115.51 244.0475 115.925 ;
      RECT  244.4625 115.51 244.7525 115.925 ;
      RECT  245.1675 115.51 245.4575 115.925 ;
      RECT  245.8725 115.51 246.1625 115.925 ;
      RECT  246.5775 115.51 246.8675 115.925 ;
      RECT  247.2825 115.51 247.5725 115.925 ;
      RECT  247.9875 115.51 248.2775 115.925 ;
      RECT  248.6925 115.51 248.9825 115.925 ;
      RECT  249.3975 115.51 249.6875 115.925 ;
      RECT  250.1025 115.51 250.3925 115.925 ;
      RECT  250.8075 115.51 251.0975 115.925 ;
      RECT  251.5125 115.51 251.8025 115.925 ;
      RECT  252.2175 115.51 252.5075 115.925 ;
      RECT  252.9225 115.51 253.2125 115.925 ;
      RECT  253.6275 115.51 253.9175 115.925 ;
      RECT  254.3325 115.51 254.6225 115.925 ;
      RECT  255.0375 115.51 255.3275 115.925 ;
      RECT  255.7425 115.51 256.0325 115.925 ;
      RECT  256.4475 115.51 256.7375 115.925 ;
      RECT  257.1525 115.51 257.4425 115.925 ;
      RECT  257.8575 115.51 258.1475 115.925 ;
      RECT  258.5625 115.51 258.8525 115.925 ;
      RECT  259.2675 115.51 259.5575 115.925 ;
      RECT  259.9725 115.51 260.2625 115.925 ;
      RECT  260.6775 115.51 260.9675 115.925 ;
      RECT  261.3825 115.51 261.6725 115.925 ;
      RECT  262.0875 115.51 262.3775 115.925 ;
      RECT  262.7925 115.51 263.0825 115.925 ;
      RECT  263.4975 115.51 263.7875 115.925 ;
      RECT  264.2025 115.51 264.4925 115.925 ;
      RECT  264.9075 115.51 265.1975 115.925 ;
      RECT  265.6125 115.51 265.9025 115.925 ;
      RECT  266.3175 115.51 266.6075 115.925 ;
      RECT  267.0225 115.51 267.3125 115.925 ;
      RECT  267.7275 115.51 268.0175 115.925 ;
      RECT  268.4325 115.51 268.7225 115.925 ;
      RECT  269.1375 115.51 269.4275 115.925 ;
      RECT  269.8425 115.51 270.1325 115.925 ;
      RECT  270.5475 115.51 270.8375 115.925 ;
      RECT  271.2525 115.51 271.5425 115.925 ;
      RECT  271.9575 115.51 272.2475 115.925 ;
      RECT  272.6625 115.51 272.9525 115.925 ;
      RECT  273.3675 115.51 273.6575 115.925 ;
      RECT  274.0725 115.51 274.3625 115.925 ;
      RECT  274.7775 115.51 275.0675 115.925 ;
      RECT  275.4825 115.51 275.7725 115.925 ;
      RECT  276.1875 115.51 276.4775 115.925 ;
      RECT  276.8925 115.51 277.1825 115.925 ;
      RECT  277.5975 115.51 277.8875 115.925 ;
      RECT  278.3025 115.51 278.5925 115.925 ;
      RECT  279.0075 115.51 279.2975 115.925 ;
      RECT  279.7125 115.51 280.0025 115.925 ;
      RECT  280.4175 115.51 280.7075 115.925 ;
      RECT  281.1225 115.51 281.4125 115.925 ;
      RECT  281.8275 115.51 282.1175 115.925 ;
      RECT  282.5325 115.51 282.8225 115.925 ;
      RECT  283.2375 115.51 283.5275 115.925 ;
      RECT  283.9425 115.51 284.2325 115.925 ;
      RECT  284.6475 115.51 284.9375 115.925 ;
      RECT  285.3525 115.51 285.6425 115.925 ;
      RECT  286.0575 115.51 286.3475 115.925 ;
      RECT  286.7625 115.51 287.0525 115.925 ;
      RECT  287.4675 115.51 287.7575 115.925 ;
      RECT  288.1725 115.51 288.4625 115.925 ;
      RECT  288.8775 115.51 289.1675 115.925 ;
      RECT  289.5825 115.51 289.8725 115.925 ;
      RECT  290.2875 115.51 290.5775 115.925 ;
      RECT  290.9925 115.51 291.2825 115.925 ;
      RECT  291.6975 115.51 291.9875 115.925 ;
      RECT  292.4025 115.51 292.6925 115.925 ;
      RECT  293.1075 115.51 293.3975 115.925 ;
      RECT  293.8125 115.51 294.1025 115.925 ;
      RECT  294.5175 115.51 294.8075 115.925 ;
      RECT  295.2225 115.51 295.5125 115.925 ;
      RECT  295.9275 115.51 296.2175 115.925 ;
      RECT  296.6325 115.51 296.9225 115.925 ;
      RECT  297.3375 115.51 297.6275 115.925 ;
      RECT  298.0425 115.51 298.3325 115.925 ;
      RECT  298.7475 115.51 299.0375 115.925 ;
      RECT  299.4525 115.51 299.7425 115.925 ;
      RECT  300.1575 115.51 300.4475 115.925 ;
      RECT  300.8625 115.51 301.1525 115.925 ;
      RECT  301.5675 115.51 301.8575 115.925 ;
      RECT  302.2725 115.51 302.5625 115.925 ;
      RECT  302.9775 115.51 303.2675 115.925 ;
      RECT  303.6825 115.51 303.9725 115.925 ;
      RECT  304.3875 115.51 304.6775 115.925 ;
      RECT  305.0925 115.51 305.3825 115.925 ;
      RECT  305.7975 115.51 306.0875 115.925 ;
      RECT  306.5025 115.51 306.7925 115.925 ;
      RECT  307.2075 115.51 307.4975 115.925 ;
      RECT  307.9125 115.51 308.2025 115.925 ;
      RECT  308.6175 115.51 308.9075 115.925 ;
      RECT  309.3225 115.51 309.6125 115.925 ;
      RECT  310.0275 115.51 310.3175 115.925 ;
      RECT  310.7325 115.51 311.0225 115.925 ;
      RECT  311.4375 115.51 311.7275 115.925 ;
      RECT  312.1425 115.51 312.4325 115.925 ;
      RECT  312.8475 115.51 313.1375 115.925 ;
      RECT  313.5525 115.51 313.8425 115.925 ;
      RECT  314.2575 115.51 314.5475 115.925 ;
      RECT  314.9625 115.51 315.2525 115.925 ;
      RECT  315.6675 115.51 315.9575 115.925 ;
      RECT  316.3725 115.51 316.6625 115.925 ;
      RECT  317.0775 115.51 317.3675 115.925 ;
      RECT  317.7825 115.51 318.0725 115.925 ;
      RECT  318.4875 115.51 318.7775 115.925 ;
      RECT  319.1925 115.51 319.4825 115.925 ;
      RECT  319.8975 115.51 320.1875 115.925 ;
      RECT  320.6025 115.51 320.8925 115.925 ;
      RECT  321.3075 115.51 321.5975 115.925 ;
      RECT  322.0125 115.51 322.3025 115.925 ;
      RECT  322.7175 115.51 323.0075 115.925 ;
      RECT  323.4225 115.51 323.7125 115.925 ;
      RECT  324.1275 115.51 324.4175 115.925 ;
      RECT  324.8325 115.51 325.1225 115.925 ;
      RECT  325.5375 115.51 325.8275 115.925 ;
      RECT  326.2425 115.51 326.5325 115.925 ;
      RECT  326.9475 115.51 327.2375 115.925 ;
      RECT  327.6525 115.51 327.9425 115.925 ;
      RECT  328.3575 115.51 328.6475 115.925 ;
      RECT  329.0625 115.51 329.3525 115.925 ;
      RECT  329.7675 115.51 330.0575 115.925 ;
      RECT  330.4725 115.51 330.7625 115.925 ;
      RECT  331.1775 115.51 331.4675 115.925 ;
      RECT  331.8825 115.51 332.1725 115.925 ;
      RECT  332.5875 115.51 332.8775 115.925 ;
      RECT  333.2925 115.51 333.5825 115.925 ;
      RECT  333.9975 115.51 334.2875 115.925 ;
      RECT  334.7025 115.51 334.9925 115.925 ;
      RECT  335.4075 115.51 335.6975 115.925 ;
      RECT  336.1125 115.51 336.4025 115.925 ;
      RECT  336.8175 115.51 337.1075 115.925 ;
      RECT  337.5225 115.51 337.8125 115.925 ;
      RECT  338.2275 115.51 338.5175 115.925 ;
      RECT  338.9325 115.51 339.2225 115.925 ;
      RECT  339.6375 115.51 339.9275 115.925 ;
      RECT  340.3425 115.51 340.6325 115.925 ;
      RECT  341.0475 115.51 341.3375 115.925 ;
      RECT  341.7525 115.51 342.0425 115.925 ;
      RECT  342.4575 115.51 342.7475 115.925 ;
      RECT  343.1625 115.51 343.4525 115.925 ;
      RECT  343.8675 115.51 344.1575 115.925 ;
      RECT  344.5725 115.51 344.8625 115.925 ;
      RECT  345.2775 115.51 345.5675 115.925 ;
      RECT  345.9825 115.51 346.2725 115.925 ;
      RECT  346.6875 115.51 346.9775 115.925 ;
      RECT  347.3925 115.51 347.6825 115.925 ;
      RECT  348.0975 115.51 348.3875 115.925 ;
      RECT  348.8025 115.51 349.0925 115.925 ;
      RECT  349.5075 115.51 349.7975 115.925 ;
      RECT  350.2125 115.51 350.5025 115.925 ;
      RECT  350.9175 115.51 351.2075 115.925 ;
      RECT  351.6225 115.51 351.9125 115.925 ;
      RECT  352.3275 115.51 352.6175 115.925 ;
      RECT  353.0325 115.51 353.3225 115.925 ;
      RECT  353.7375 115.51 354.0275 115.925 ;
      RECT  354.4425 115.51 354.7325 115.925 ;
      RECT  355.1475 115.51 355.4375 115.925 ;
      RECT  355.8525 115.51 356.1425 115.925 ;
      RECT  356.5575 115.51 356.8475 115.925 ;
      RECT  357.2625 115.51 357.5525 115.925 ;
      RECT  357.9675 115.51 358.2575 115.925 ;
      RECT  358.6725 115.51 358.9625 115.925 ;
      RECT  359.3775 115.51 359.6675 115.925 ;
      RECT  360.0825 115.51 360.3725 115.925 ;
      RECT  360.7875 115.51 361.0775 115.925 ;
      RECT  361.4925 115.51 361.7825 115.925 ;
      RECT  362.1975 115.51 362.4875 115.925 ;
      RECT  362.9025 115.51 363.1925 115.925 ;
      RECT  363.6075 115.51 363.8975 115.925 ;
      RECT  364.3125 115.51 364.6025 115.925 ;
      RECT  365.0175 115.51 365.3075 115.925 ;
      RECT  365.7225 115.51 366.0125 115.925 ;
      RECT  366.4275 115.51 366.7175 115.925 ;
      RECT  367.1325 115.51 367.4225 115.925 ;
      RECT  367.8375 115.51 368.1275 115.925 ;
      RECT  368.5425 115.51 368.8325 115.925 ;
      RECT  369.2475 115.51 369.5375 115.925 ;
      RECT  369.9525 115.51 370.2425 115.925 ;
      RECT  370.6575 115.51 370.9475 115.925 ;
      RECT  371.3625 115.51 371.6525 115.925 ;
      RECT  372.0675 115.51 372.3575 115.925 ;
      RECT  372.7725 115.51 373.0625 115.925 ;
      RECT  373.4775 115.51 373.7675 115.925 ;
      RECT  374.1825 115.51 374.4725 115.925 ;
      RECT  374.8875 115.51 375.1775 115.925 ;
      RECT  375.5925 115.51 375.8825 115.925 ;
      RECT  376.2975 115.51 376.5875 115.925 ;
      RECT  377.0025 115.51 377.2925 115.925 ;
      RECT  377.7075 115.51 377.9975 115.925 ;
      RECT  378.4125 115.51 378.7025 115.925 ;
      RECT  379.1175 115.51 379.4075 115.925 ;
      RECT  379.8225 115.51 380.1125 115.925 ;
      RECT  380.5275 115.51 380.8175 115.925 ;
      RECT  381.2325 115.51 381.5225 115.925 ;
      RECT  381.9375 115.51 382.2275 115.925 ;
      RECT  382.6425 115.51 382.9325 115.925 ;
      RECT  383.3475 115.51 383.6375 115.925 ;
      RECT  384.0525 115.51 384.3425 115.925 ;
      RECT  384.7575 115.51 385.0475 115.925 ;
      RECT  385.4625 115.51 385.7525 115.925 ;
      RECT  386.1675 115.51 386.4575 115.925 ;
      RECT  386.8725 115.51 387.1625 115.925 ;
      RECT  387.5775 115.51 387.8675 115.925 ;
      RECT  388.2825 115.51 388.5725 115.925 ;
      RECT  388.9875 115.51 389.2775 115.925 ;
      RECT  389.6925 115.51 389.9825 115.925 ;
      RECT  390.3975 115.51 390.6875 115.925 ;
      RECT  391.1025 115.51 391.3925 115.925 ;
      RECT  391.8075 115.51 392.0975 115.925 ;
      RECT  392.5125 115.51 392.8025 115.925 ;
      RECT  393.2175 115.51 393.5075 115.925 ;
      RECT  393.9225 115.51 394.2125 115.925 ;
      RECT  394.6275 115.51 394.9175 115.925 ;
      RECT  395.3325 115.51 395.6225 115.925 ;
      RECT  396.0375 115.51 396.3275 115.925 ;
      RECT  396.7425 115.51 397.0325 115.925 ;
      RECT  397.4475 115.51 397.7375 115.925 ;
      RECT  398.1525 115.51 398.4425 115.925 ;
      RECT  398.8575 115.51 399.1475 115.925 ;
      RECT  399.5625 115.51 399.8525 115.925 ;
      RECT  400.2675 115.51 400.5575 115.925 ;
      RECT  400.9725 115.51 401.2625 115.925 ;
      RECT  401.6775 115.51 401.9675 115.925 ;
      RECT  402.3825 115.51 402.6725 115.925 ;
      RECT  403.0875 115.51 403.3775 115.925 ;
      RECT  403.7925 115.51 404.0825 115.925 ;
      RECT  404.4975 115.51 404.7875 115.925 ;
      RECT  405.2025 115.51 405.4925 115.925 ;
      RECT  405.9075 115.51 406.1975 115.925 ;
      RECT  406.6125 115.51 406.9025 115.925 ;
      RECT  407.3175 115.51 407.6075 115.925 ;
      RECT  408.0225 115.51 408.3125 115.925 ;
      RECT  408.7275 115.51 409.0175 115.925 ;
      RECT  409.4325 115.51 409.7225 115.925 ;
      RECT  410.1375 115.51 410.4275 115.925 ;
      RECT  410.8425 115.51 411.1325 115.925 ;
      RECT  411.5475 115.51 411.8375 115.925 ;
      RECT  412.2525 115.51 412.5425 115.925 ;
      RECT  412.9575 115.51 413.2475 115.925 ;
      RECT  413.6625 115.51 413.9525 115.925 ;
      RECT  414.3675 115.51 414.6575 115.925 ;
      RECT  415.0725 115.51 415.3625 115.925 ;
      RECT  415.7775 115.51 416.0675 115.925 ;
      RECT  416.4825 115.51 416.7725 115.925 ;
      RECT  417.1875 115.51 417.4775 115.925 ;
      RECT  417.8925 115.51 418.1825 115.925 ;
      RECT  418.5975 115.51 418.8875 115.925 ;
      RECT  419.3025 115.51 419.5925 115.925 ;
      RECT  420.0075 115.51 420.2975 115.925 ;
      RECT  420.7125 115.51 421.0025 115.925 ;
      RECT  421.4175 115.51 421.7075 115.925 ;
      RECT  422.1225 115.51 422.4125 115.925 ;
      RECT  422.8275 115.51 423.1175 115.925 ;
      RECT  423.5325 115.51 423.8225 115.925 ;
      RECT  424.2375 115.51 424.5275 115.925 ;
      RECT  424.9425 115.51 425.2325 115.925 ;
      RECT  425.6475 115.51 425.9375 115.925 ;
      RECT  426.3525 115.51 426.6425 115.925 ;
      RECT  427.0575 115.51 427.3475 115.925 ;
      RECT  427.7625 115.51 428.0525 115.925 ;
      RECT  428.4675 115.51 428.7575 115.925 ;
      RECT  429.1725 115.51 429.4625 115.925 ;
      RECT  429.8775 115.51 430.1675 115.925 ;
      RECT  430.5825 115.51 430.8725 115.925 ;
      RECT  431.2875 115.51 431.5775 115.925 ;
      RECT  431.9925 115.51 432.2825 115.925 ;
      RECT  432.6975 115.51 432.9875 115.925 ;
      RECT  433.4025 115.51 433.6925 115.925 ;
      RECT  434.1075 115.51 434.3975 115.925 ;
      RECT  434.8125 115.51 435.1025 115.925 ;
      RECT  435.5175 115.51 435.8075 115.925 ;
      RECT  436.2225 115.51 436.5125 115.925 ;
      RECT  436.9275 115.51 437.2175 115.925 ;
      RECT  437.6325 115.51 437.9225 115.925 ;
      RECT  438.3375 115.51 438.6275 115.925 ;
      RECT  439.0425 115.51 439.3325 115.925 ;
      RECT  439.7475 115.51 440.0375 115.925 ;
      RECT  440.4525 115.51 440.7425 115.925 ;
      RECT  441.1575 115.51 441.4475 115.925 ;
      RECT  441.8625 115.51 442.1525 115.925 ;
      RECT  442.5675 115.51 442.8575 115.925 ;
      RECT  443.2725 115.51 443.5625 115.925 ;
      RECT  443.9775 115.51 444.2675 115.925 ;
      RECT  444.6825 115.51 444.9725 115.925 ;
      RECT  445.3875 115.51 445.6775 115.925 ;
      RECT  446.0925 115.51 446.3825 115.925 ;
      RECT  446.7975 115.51 447.0875 115.925 ;
      RECT  447.5025 115.51 447.7925 115.925 ;
      RECT  448.2075 115.51 448.4975 115.925 ;
      RECT  448.9125 115.51 449.2025 115.925 ;
      RECT  449.6175 115.51 449.9075 115.925 ;
      RECT  450.3225 115.51 450.6125 115.925 ;
      RECT  451.0275 115.51 451.3175 115.925 ;
      RECT  451.7325 115.51 452.0225 115.925 ;
      RECT  452.4375 115.51 452.7275 115.925 ;
      RECT  453.1425 115.51 453.4325 115.925 ;
      RECT  453.8475 115.51 454.1375 115.925 ;
      RECT  454.5525 115.51 454.8425 115.925 ;
      RECT  455.2575 115.51 455.5475 115.925 ;
      RECT  455.9625 115.51 456.2525 115.925 ;
      RECT  456.6675 115.51 456.9575 115.925 ;
      RECT  457.3725 115.51 457.6625 115.925 ;
      RECT  458.0775 115.51 458.3675 115.925 ;
      RECT  458.7825 115.51 459.0725 115.925 ;
      RECT  459.4875 115.51 459.7775 115.925 ;
      RECT  460.1925 115.51 460.4825 115.925 ;
      RECT  460.8975 115.51 461.1875 115.925 ;
      RECT  461.6025 115.51 461.8925 115.925 ;
      RECT  462.3075 115.51 462.5975 115.925 ;
      RECT  463.0125 115.51 463.3025 115.925 ;
      RECT  463.7175 115.51 464.0075 115.925 ;
      RECT  464.4225 115.51 464.7125 115.925 ;
      RECT  465.1275 115.51 465.4175 115.925 ;
      RECT  465.8325 115.51 466.1225 115.925 ;
      RECT  466.5375 115.51 466.8275 115.925 ;
      RECT  467.2425 115.51 467.5325 115.925 ;
      RECT  467.9475 115.51 468.2375 115.925 ;
      RECT  468.6525 115.51 468.9425 115.925 ;
      RECT  469.3575 115.51 469.6475 115.925 ;
      RECT  470.0625 115.51 470.3525 115.925 ;
      RECT  470.7675 115.51 471.0575 115.925 ;
      RECT  471.4725 115.51 471.7625 115.925 ;
      RECT  472.1775 115.51 472.4675 115.925 ;
      RECT  472.8825 115.51 473.1725 115.925 ;
      RECT  473.5875 115.51 473.8775 115.925 ;
      RECT  474.2925 115.51 474.5825 115.925 ;
      RECT  474.9975 115.51 475.2875 115.925 ;
      RECT  475.7025 115.51 475.9925 115.925 ;
      RECT  476.4075 115.51 476.6975 115.925 ;
      RECT  477.1125 115.51 477.4025 115.925 ;
      RECT  477.8175 115.51 478.1075 115.925 ;
      RECT  478.5225 115.51 478.8125 115.925 ;
      RECT  479.2275 115.51 479.5175 115.925 ;
      RECT  479.9325 115.51 480.2225 115.925 ;
      RECT  480.6375 115.51 480.9275 115.925 ;
      RECT  481.3425 115.51 481.6325 115.925 ;
      RECT  482.0475 115.51 482.3375 115.925 ;
      RECT  482.7525 115.51 483.0425 115.925 ;
      RECT  483.4575 115.51 483.7475 115.925 ;
      RECT  484.1625 115.51 484.4525 115.925 ;
      RECT  484.8675 115.51 485.1575 115.925 ;
      RECT  485.5725 115.51 485.8625 115.925 ;
      RECT  486.2775 115.51 486.5675 115.925 ;
      RECT  486.9825 115.51 487.2725 115.925 ;
      RECT  487.6875 115.51 487.9775 115.925 ;
      RECT  488.3925 115.51 488.6825 115.925 ;
      RECT  489.0975 115.51 489.3875 115.925 ;
      RECT  489.8025 115.51 490.0925 115.925 ;
      RECT  490.5075 115.51 490.7975 115.925 ;
      RECT  491.2125 115.51 491.5025 115.925 ;
      RECT  491.9175 115.51 492.2075 115.925 ;
      RECT  492.6225 115.51 492.9125 115.925 ;
      RECT  493.3275 115.51 493.6175 115.925 ;
      RECT  494.0325 115.51 494.3225 115.925 ;
      RECT  494.7375 115.51 495.0275 115.925 ;
      RECT  495.4425 115.51 495.7325 115.925 ;
      RECT  496.1475 115.51 496.4375 115.925 ;
      RECT  496.8525 115.51 497.1425 115.925 ;
      RECT  497.5575 115.51 497.8475 115.925 ;
      RECT  498.2625 115.51 498.5525 115.925 ;
      RECT  498.9675 115.51 499.2575 115.925 ;
      RECT  499.6725 115.51 499.9625 115.925 ;
      RECT  500.3775 115.51 500.6675 115.925 ;
      RECT  501.0825 115.51 501.3725 115.925 ;
      RECT  501.7875 115.51 502.0775 115.925 ;
      RECT  502.4925 115.51 502.7825 115.925 ;
      RECT  503.1975 115.51 503.4875 115.925 ;
      RECT  503.9025 115.51 504.1925 115.925 ;
      RECT  504.6075 115.51 504.8975 115.925 ;
      RECT  505.3125 115.51 505.6025 115.925 ;
      RECT  506.0175 115.51 506.3075 115.925 ;
      RECT  506.7225 115.51 507.0125 115.925 ;
      RECT  507.4275 115.51 507.7175 115.925 ;
      RECT  508.1325 115.51 508.4225 115.925 ;
      RECT  508.8375 115.51 509.1275 115.925 ;
      RECT  509.5425 115.51 509.8325 115.925 ;
      RECT  510.2475 115.51 510.5375 115.925 ;
      RECT  510.9525 115.51 511.2425 115.925 ;
      RECT  511.6575 115.51 511.9475 115.925 ;
      RECT  512.3625 115.51 512.6525 115.925 ;
      RECT  513.0675 115.51 513.3575 115.925 ;
      RECT  513.7725 115.51 514.0625 115.925 ;
      RECT  514.4775 115.51 514.7675 115.925 ;
      RECT  515.1825 115.51 515.4725 115.925 ;
      RECT  515.8875 115.51 516.1775 115.925 ;
      RECT  516.5925 115.51 516.8825 115.925 ;
      RECT  517.2975 115.51 517.5875 115.925 ;
      RECT  518.0025 115.51 518.2925 115.925 ;
      RECT  518.7075 115.51 518.9975 115.925 ;
      RECT  519.4125 115.51 519.7025 115.925 ;
      RECT  520.1175 115.51 520.4075 115.925 ;
      RECT  520.8225 115.51 521.1125 115.925 ;
      RECT  521.5275 115.51 521.8175 115.925 ;
      RECT  522.2325 115.51 522.5225 115.925 ;
      RECT  522.9375 115.51 523.2275 115.925 ;
      RECT  523.6425 115.51 1593.48 115.925 ;
      RECT  0.14 1.26 1.26 2.24 ;
      RECT  0.14 2.24 1.26 4.0975 ;
      RECT  1.26 2.24 126.205 4.0975 ;
      RECT  126.205 2.24 126.62 4.0975 ;
      RECT  126.62 2.24 1592.36 4.0975 ;
      RECT  1592.36 1.26 1593.48 2.24 ;
      RECT  1592.36 2.24 1593.48 4.0975 ;
      RECT  126.205 4.5125 126.62 216.58 ;
      RECT  0.14 148.9975 1.26 216.58 ;
      RECT  0.14 216.58 1.26 217.56 ;
      RECT  1.26 148.9975 120.485 216.58 ;
      RECT  120.9 148.9975 126.205 216.58 ;
      RECT  120.485 161.6075 120.9 216.58 ;
      RECT  126.62 115.925 162.9725 216.58 ;
      RECT  162.9725 115.925 163.3875 216.58 ;
      RECT  163.3875 115.925 1592.36 216.58 ;
      RECT  1592.36 115.925 1593.48 216.58 ;
      RECT  1592.36 216.58 1593.48 217.56 ;
      RECT  0.14 0.84 1.26 1.26 ;
      RECT  1.26 0.84 126.205 1.26 ;
      RECT  126.205 0.84 126.62 1.26 ;
      RECT  126.62 0.84 1592.36 1.26 ;
      RECT  1592.36 0.84 1593.48 1.26 ;
      RECT  126.205 217.56 126.62 217.98 ;
      RECT  0.14 217.56 1.26 217.98 ;
      RECT  1.26 217.56 120.485 217.98 ;
      RECT  120.9 217.56 126.205 217.98 ;
      RECT  120.485 217.56 120.9 217.98 ;
      RECT  126.62 217.56 162.9725 217.98 ;
      RECT  162.9725 217.56 163.3875 217.98 ;
      RECT  163.3875 217.56 1592.36 217.98 ;
      RECT  1592.36 217.56 1593.48 217.98 ;
   LAYER  metal4 ;
      RECT  1591.24 0.14 1592.5 1.12 ;
      RECT  1591.24 217.7 1592.5 218.68 ;
      RECT  2.38 1.12 1591.24 217.7 ;
      RECT  1592.5 0.14 1592.64 1.12 ;
      RECT  1592.5 1.12 1592.64 217.7 ;
      RECT  1592.5 217.7 1592.64 218.68 ;
      RECT  0.98 0.14 1591.24 1.12 ;
      RECT  0.98 217.7 1591.24 218.68 ;
      RECT  0.98 1.12 1.12 217.7 ;
   END
END    freepdk45_sram_1rw0r_45x512
END    LIBRARY
