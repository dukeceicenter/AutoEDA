../macros/freepdk45_sram_1w1r_32x72/freepdk45_sram_1w1r_32x72.lef