../macros/freepdk45_sram_1w1r_34x128_32/freepdk45_sram_1w1r_34x128_32.lef