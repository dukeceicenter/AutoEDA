VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_40x240
   CLASS BLOCK ;
   SIZE 752.775 BY 128.2725 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.59 1.105 66.725 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.45 1.105 69.585 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.31 1.105 72.445 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.17 1.105 75.305 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.03 1.105 78.165 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.89 1.105 81.025 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.75 1.105 83.885 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.61 1.105 86.745 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.47 1.105 89.605 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.33 1.105 92.465 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.19 1.105 95.325 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.05 1.105 98.185 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.91 1.105 101.045 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.77 1.105 103.905 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.63 1.105 106.765 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.49 1.105 109.625 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.35 1.105 112.485 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.21 1.105 115.345 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.07 1.105 118.205 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.93 1.105 121.065 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.79 1.105 123.925 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.65 1.105 126.785 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.51 1.105 129.645 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.37 1.105 132.505 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.23 1.105 135.365 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.09 1.105 138.225 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.95 1.105 141.085 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.81 1.105 143.945 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.67 1.105 146.805 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.53 1.105 149.665 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.39 1.105 152.525 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.25 1.105 155.385 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.11 1.105 158.245 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.97 1.105 161.105 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.83 1.105 163.965 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.69 1.105 166.825 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.55 1.105 169.685 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.41 1.105 172.545 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.27 1.105 175.405 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.13 1.105 178.265 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.99 1.105 181.125 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.85 1.105 183.985 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.71 1.105 186.845 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.57 1.105 189.705 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.43 1.105 192.565 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.29 1.105 195.425 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.15 1.105 198.285 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.01 1.105 201.145 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.87 1.105 204.005 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.73 1.105 206.865 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.59 1.105 209.725 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.45 1.105 212.585 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.31 1.105 215.445 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.17 1.105 218.305 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.03 1.105 221.165 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.89 1.105 224.025 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.75 1.105 226.885 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.61 1.105 229.745 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.47 1.105 232.605 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.33 1.105 235.465 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.19 1.105 238.325 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.05 1.105 241.185 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.91 1.105 244.045 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.77 1.105 246.905 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.63 1.105 249.765 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.49 1.105 252.625 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.35 1.105 255.485 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.21 1.105 258.345 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.07 1.105 261.205 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.93 1.105 264.065 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.79 1.105 266.925 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.65 1.105 269.785 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.51 1.105 272.645 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.37 1.105 275.505 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.23 1.105 278.365 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.09 1.105 281.225 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.95 1.105 284.085 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.81 1.105 286.945 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.67 1.105 289.805 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.53 1.105 292.665 1.24 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.39 1.105 295.525 1.24 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.25 1.105 298.385 1.24 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.11 1.105 301.245 1.24 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.97 1.105 304.105 1.24 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.83 1.105 306.965 1.24 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.69 1.105 309.825 1.24 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.55 1.105 312.685 1.24 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.41 1.105 315.545 1.24 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.27 1.105 318.405 1.24 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.13 1.105 321.265 1.24 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.99 1.105 324.125 1.24 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.85 1.105 326.985 1.24 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.71 1.105 329.845 1.24 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.57 1.105 332.705 1.24 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.43 1.105 335.565 1.24 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.29 1.105 338.425 1.24 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.15 1.105 341.285 1.24 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.01 1.105 344.145 1.24 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.87 1.105 347.005 1.24 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.73 1.105 349.865 1.24 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.59 1.105 352.725 1.24 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.45 1.105 355.585 1.24 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.31 1.105 358.445 1.24 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.17 1.105 361.305 1.24 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.03 1.105 364.165 1.24 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.89 1.105 367.025 1.24 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.75 1.105 369.885 1.24 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.61 1.105 372.745 1.24 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.47 1.105 375.605 1.24 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.33 1.105 378.465 1.24 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.19 1.105 381.325 1.24 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.05 1.105 384.185 1.24 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.91 1.105 387.045 1.24 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.77 1.105 389.905 1.24 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.63 1.105 392.765 1.24 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.49 1.105 395.625 1.24 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.35 1.105 398.485 1.24 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.21 1.105 401.345 1.24 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.07 1.105 404.205 1.24 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.93 1.105 407.065 1.24 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.79 1.105 409.925 1.24 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.65 1.105 412.785 1.24 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.51 1.105 415.645 1.24 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.37 1.105 418.505 1.24 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.23 1.105 421.365 1.24 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.09 1.105 424.225 1.24 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.95 1.105 427.085 1.24 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.81 1.105 429.945 1.24 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.67 1.105 432.805 1.24 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.53 1.105 435.665 1.24 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.39 1.105 438.525 1.24 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.25 1.105 441.385 1.24 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.11 1.105 444.245 1.24 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.97 1.105 447.105 1.24 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.83 1.105 449.965 1.24 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.69 1.105 452.825 1.24 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.55 1.105 455.685 1.24 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.41 1.105 458.545 1.24 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.27 1.105 461.405 1.24 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.13 1.105 464.265 1.24 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.99 1.105 467.125 1.24 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.85 1.105 469.985 1.24 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.71 1.105 472.845 1.24 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.57 1.105 475.705 1.24 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.43 1.105 478.565 1.24 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.29 1.105 481.425 1.24 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.15 1.105 484.285 1.24 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.01 1.105 487.145 1.24 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.87 1.105 490.005 1.24 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.73 1.105 492.865 1.24 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.59 1.105 495.725 1.24 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.45 1.105 498.585 1.24 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.31 1.105 501.445 1.24 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.17 1.105 504.305 1.24 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.03 1.105 507.165 1.24 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.89 1.105 510.025 1.24 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.75 1.105 512.885 1.24 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.61 1.105 515.745 1.24 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.47 1.105 518.605 1.24 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.33 1.105 521.465 1.24 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  524.19 1.105 524.325 1.24 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.05 1.105 527.185 1.24 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  529.91 1.105 530.045 1.24 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  532.77 1.105 532.905 1.24 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  535.63 1.105 535.765 1.24 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  538.49 1.105 538.625 1.24 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  541.35 1.105 541.485 1.24 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  544.21 1.105 544.345 1.24 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  547.07 1.105 547.205 1.24 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  549.93 1.105 550.065 1.24 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  552.79 1.105 552.925 1.24 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  555.65 1.105 555.785 1.24 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  558.51 1.105 558.645 1.24 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  561.37 1.105 561.505 1.24 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  564.23 1.105 564.365 1.24 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  567.09 1.105 567.225 1.24 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  569.95 1.105 570.085 1.24 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  572.81 1.105 572.945 1.24 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  575.67 1.105 575.805 1.24 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  578.53 1.105 578.665 1.24 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  581.39 1.105 581.525 1.24 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  584.25 1.105 584.385 1.24 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  587.11 1.105 587.245 1.24 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  589.97 1.105 590.105 1.24 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  592.83 1.105 592.965 1.24 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  595.69 1.105 595.825 1.24 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  598.55 1.105 598.685 1.24 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  601.41 1.105 601.545 1.24 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  604.27 1.105 604.405 1.24 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  607.13 1.105 607.265 1.24 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  609.99 1.105 610.125 1.24 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  612.85 1.105 612.985 1.24 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  615.71 1.105 615.845 1.24 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  618.57 1.105 618.705 1.24 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  621.43 1.105 621.565 1.24 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  624.29 1.105 624.425 1.24 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  627.15 1.105 627.285 1.24 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  630.01 1.105 630.145 1.24 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  632.87 1.105 633.005 1.24 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  635.73 1.105 635.865 1.24 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  638.59 1.105 638.725 1.24 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  641.45 1.105 641.585 1.24 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  644.31 1.105 644.445 1.24 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  647.17 1.105 647.305 1.24 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  650.03 1.105 650.165 1.24 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  652.89 1.105 653.025 1.24 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  655.75 1.105 655.885 1.24 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  658.61 1.105 658.745 1.24 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  661.47 1.105 661.605 1.24 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  664.33 1.105 664.465 1.24 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  667.19 1.105 667.325 1.24 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  670.05 1.105 670.185 1.24 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  672.91 1.105 673.045 1.24 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  675.77 1.105 675.905 1.24 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  678.63 1.105 678.765 1.24 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  681.49 1.105 681.625 1.24 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  684.35 1.105 684.485 1.24 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  687.21 1.105 687.345 1.24 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  690.07 1.105 690.205 1.24 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  692.93 1.105 693.065 1.24 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  695.79 1.105 695.925 1.24 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  698.65 1.105 698.785 1.24 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  701.51 1.105 701.645 1.24 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  704.37 1.105 704.505 1.24 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  707.23 1.105 707.365 1.24 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  710.09 1.105 710.225 1.24 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  712.95 1.105 713.085 1.24 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  715.81 1.105 715.945 1.24 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  718.67 1.105 718.805 1.24 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  721.53 1.105 721.665 1.24 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  724.39 1.105 724.525 1.24 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  727.25 1.105 727.385 1.24 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  730.11 1.105 730.245 1.24 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  732.97 1.105 733.105 1.24 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  735.83 1.105 735.965 1.24 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  738.69 1.105 738.825 1.24 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  741.55 1.105 741.685 1.24 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  744.41 1.105 744.545 1.24 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  747.27 1.105 747.405 1.24 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  750.13 1.105 750.265 1.24 ;
      END
   END din0[239]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 75.34 61.005 75.475 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 78.07 61.005 78.205 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 80.28 61.005 80.415 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 83.01 61.005 83.145 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 85.22 61.005 85.355 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 87.95 61.005 88.085 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.05 49.21 399.185 49.345 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.05 46.48 399.185 46.615 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.05 44.27 399.185 44.405 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.05 41.54 399.185 41.675 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.05 39.33 399.185 39.465 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.05 36.6 399.185 36.735 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 30.75 0.42 30.885 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  459.775 127.03 459.91 127.165 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 30.835 6.3825 30.97 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.6725 126.945 453.8075 127.08 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.8975 120.3225 89.0325 120.4575 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.0725 120.3225 90.2075 120.4575 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.2475 120.3225 91.3825 120.4575 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.4225 120.3225 92.5575 120.4575 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.5975 120.3225 93.7325 120.4575 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.7725 120.3225 94.9075 120.4575 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.9475 120.3225 96.0825 120.4575 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.1225 120.3225 97.2575 120.4575 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.2975 120.3225 98.4325 120.4575 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.4725 120.3225 99.6075 120.4575 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.6475 120.3225 100.7825 120.4575 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.8225 120.3225 101.9575 120.4575 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.9975 120.3225 103.1325 120.4575 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.1725 120.3225 104.3075 120.4575 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.3475 120.3225 105.4825 120.4575 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.5225 120.3225 106.6575 120.4575 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.6975 120.3225 107.8325 120.4575 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.8725 120.3225 109.0075 120.4575 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.0475 120.3225 110.1825 120.4575 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.2225 120.3225 111.3575 120.4575 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.3975 120.3225 112.5325 120.4575 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.5725 120.3225 113.7075 120.4575 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.7475 120.3225 114.8825 120.4575 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.9225 120.3225 116.0575 120.4575 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.0975 120.3225 117.2325 120.4575 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.2725 120.3225 118.4075 120.4575 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.4475 120.3225 119.5825 120.4575 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.6225 120.3225 120.7575 120.4575 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.7975 120.3225 121.9325 120.4575 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.9725 120.3225 123.1075 120.4575 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.1475 120.3225 124.2825 120.4575 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.3225 120.3225 125.4575 120.4575 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.4975 120.3225 126.6325 120.4575 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.6725 120.3225 127.8075 120.4575 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.8475 120.3225 128.9825 120.4575 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.0225 120.3225 130.1575 120.4575 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.1975 120.3225 131.3325 120.4575 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.3725 120.3225 132.5075 120.4575 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.5475 120.3225 133.6825 120.4575 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.7225 120.3225 134.8575 120.4575 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.8975 120.3225 136.0325 120.4575 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.0725 120.3225 137.2075 120.4575 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.2475 120.3225 138.3825 120.4575 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.4225 120.3225 139.5575 120.4575 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.5975 120.3225 140.7325 120.4575 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.7725 120.3225 141.9075 120.4575 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.9475 120.3225 143.0825 120.4575 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.1225 120.3225 144.2575 120.4575 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.2975 120.3225 145.4325 120.4575 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.4725 120.3225 146.6075 120.4575 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.6475 120.3225 147.7825 120.4575 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.8225 120.3225 148.9575 120.4575 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.9975 120.3225 150.1325 120.4575 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.1725 120.3225 151.3075 120.4575 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.3475 120.3225 152.4825 120.4575 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.5225 120.3225 153.6575 120.4575 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.6975 120.3225 154.8325 120.4575 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.8725 120.3225 156.0075 120.4575 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.0475 120.3225 157.1825 120.4575 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.2225 120.3225 158.3575 120.4575 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.3975 120.3225 159.5325 120.4575 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.5725 120.3225 160.7075 120.4575 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.7475 120.3225 161.8825 120.4575 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.9225 120.3225 163.0575 120.4575 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.0975 120.3225 164.2325 120.4575 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.2725 120.3225 165.4075 120.4575 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.4475 120.3225 166.5825 120.4575 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.6225 120.3225 167.7575 120.4575 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.7975 120.3225 168.9325 120.4575 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.9725 120.3225 170.1075 120.4575 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.1475 120.3225 171.2825 120.4575 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.3225 120.3225 172.4575 120.4575 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.4975 120.3225 173.6325 120.4575 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.6725 120.3225 174.8075 120.4575 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.8475 120.3225 175.9825 120.4575 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.0225 120.3225 177.1575 120.4575 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.1975 120.3225 178.3325 120.4575 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.3725 120.3225 179.5075 120.4575 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.5475 120.3225 180.6825 120.4575 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.7225 120.3225 181.8575 120.4575 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.8975 120.3225 183.0325 120.4575 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.0725 120.3225 184.2075 120.4575 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.2475 120.3225 185.3825 120.4575 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.4225 120.3225 186.5575 120.4575 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.5975 120.3225 187.7325 120.4575 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.7725 120.3225 188.9075 120.4575 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.9475 120.3225 190.0825 120.4575 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.1225 120.3225 191.2575 120.4575 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.2975 120.3225 192.4325 120.4575 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.4725 120.3225 193.6075 120.4575 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.6475 120.3225 194.7825 120.4575 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.8225 120.3225 195.9575 120.4575 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.9975 120.3225 197.1325 120.4575 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.1725 120.3225 198.3075 120.4575 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.3475 120.3225 199.4825 120.4575 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.5225 120.3225 200.6575 120.4575 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.6975 120.3225 201.8325 120.4575 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.8725 120.3225 203.0075 120.4575 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.0475 120.3225 204.1825 120.4575 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.2225 120.3225 205.3575 120.4575 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.3975 120.3225 206.5325 120.4575 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.5725 120.3225 207.7075 120.4575 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.7475 120.3225 208.8825 120.4575 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.9225 120.3225 210.0575 120.4575 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.0975 120.3225 211.2325 120.4575 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.2725 120.3225 212.4075 120.4575 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.4475 120.3225 213.5825 120.4575 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.6225 120.3225 214.7575 120.4575 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.7975 120.3225 215.9325 120.4575 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.9725 120.3225 217.1075 120.4575 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.1475 120.3225 218.2825 120.4575 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.3225 120.3225 219.4575 120.4575 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.4975 120.3225 220.6325 120.4575 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.6725 120.3225 221.8075 120.4575 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.8475 120.3225 222.9825 120.4575 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.0225 120.3225 224.1575 120.4575 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.1975 120.3225 225.3325 120.4575 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.3725 120.3225 226.5075 120.4575 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.5475 120.3225 227.6825 120.4575 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.7225 120.3225 228.8575 120.4575 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.8975 120.3225 230.0325 120.4575 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.0725 120.3225 231.2075 120.4575 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.2475 120.3225 232.3825 120.4575 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.4225 120.3225 233.5575 120.4575 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.5975 120.3225 234.7325 120.4575 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.7725 120.3225 235.9075 120.4575 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.9475 120.3225 237.0825 120.4575 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.1225 120.3225 238.2575 120.4575 ;
      END
   END dout1[127]
   PIN dout1[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.2975 120.3225 239.4325 120.4575 ;
      END
   END dout1[128]
   PIN dout1[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.4725 120.3225 240.6075 120.4575 ;
      END
   END dout1[129]
   PIN dout1[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.6475 120.3225 241.7825 120.4575 ;
      END
   END dout1[130]
   PIN dout1[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.8225 120.3225 242.9575 120.4575 ;
      END
   END dout1[131]
   PIN dout1[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.9975 120.3225 244.1325 120.4575 ;
      END
   END dout1[132]
   PIN dout1[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.1725 120.3225 245.3075 120.4575 ;
      END
   END dout1[133]
   PIN dout1[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.3475 120.3225 246.4825 120.4575 ;
      END
   END dout1[134]
   PIN dout1[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.5225 120.3225 247.6575 120.4575 ;
      END
   END dout1[135]
   PIN dout1[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.6975 120.3225 248.8325 120.4575 ;
      END
   END dout1[136]
   PIN dout1[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.8725 120.3225 250.0075 120.4575 ;
      END
   END dout1[137]
   PIN dout1[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.0475 120.3225 251.1825 120.4575 ;
      END
   END dout1[138]
   PIN dout1[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.2225 120.3225 252.3575 120.4575 ;
      END
   END dout1[139]
   PIN dout1[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.3975 120.3225 253.5325 120.4575 ;
      END
   END dout1[140]
   PIN dout1[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.5725 120.3225 254.7075 120.4575 ;
      END
   END dout1[141]
   PIN dout1[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.7475 120.3225 255.8825 120.4575 ;
      END
   END dout1[142]
   PIN dout1[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.9225 120.3225 257.0575 120.4575 ;
      END
   END dout1[143]
   PIN dout1[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.0975 120.3225 258.2325 120.4575 ;
      END
   END dout1[144]
   PIN dout1[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.2725 120.3225 259.4075 120.4575 ;
      END
   END dout1[145]
   PIN dout1[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.4475 120.3225 260.5825 120.4575 ;
      END
   END dout1[146]
   PIN dout1[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.6225 120.3225 261.7575 120.4575 ;
      END
   END dout1[147]
   PIN dout1[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.7975 120.3225 262.9325 120.4575 ;
      END
   END dout1[148]
   PIN dout1[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.9725 120.3225 264.1075 120.4575 ;
      END
   END dout1[149]
   PIN dout1[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.1475 120.3225 265.2825 120.4575 ;
      END
   END dout1[150]
   PIN dout1[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.3225 120.3225 266.4575 120.4575 ;
      END
   END dout1[151]
   PIN dout1[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.4975 120.3225 267.6325 120.4575 ;
      END
   END dout1[152]
   PIN dout1[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.6725 120.3225 268.8075 120.4575 ;
      END
   END dout1[153]
   PIN dout1[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.8475 120.3225 269.9825 120.4575 ;
      END
   END dout1[154]
   PIN dout1[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.0225 120.3225 271.1575 120.4575 ;
      END
   END dout1[155]
   PIN dout1[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.1975 120.3225 272.3325 120.4575 ;
      END
   END dout1[156]
   PIN dout1[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.3725 120.3225 273.5075 120.4575 ;
      END
   END dout1[157]
   PIN dout1[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.5475 120.3225 274.6825 120.4575 ;
      END
   END dout1[158]
   PIN dout1[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.7225 120.3225 275.8575 120.4575 ;
      END
   END dout1[159]
   PIN dout1[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.8975 120.3225 277.0325 120.4575 ;
      END
   END dout1[160]
   PIN dout1[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.0725 120.3225 278.2075 120.4575 ;
      END
   END dout1[161]
   PIN dout1[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.2475 120.3225 279.3825 120.4575 ;
      END
   END dout1[162]
   PIN dout1[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.4225 120.3225 280.5575 120.4575 ;
      END
   END dout1[163]
   PIN dout1[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.5975 120.3225 281.7325 120.4575 ;
      END
   END dout1[164]
   PIN dout1[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  282.7725 120.3225 282.9075 120.4575 ;
      END
   END dout1[165]
   PIN dout1[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.9475 120.3225 284.0825 120.4575 ;
      END
   END dout1[166]
   PIN dout1[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.1225 120.3225 285.2575 120.4575 ;
      END
   END dout1[167]
   PIN dout1[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.2975 120.3225 286.4325 120.4575 ;
      END
   END dout1[168]
   PIN dout1[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.4725 120.3225 287.6075 120.4575 ;
      END
   END dout1[169]
   PIN dout1[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.6475 120.3225 288.7825 120.4575 ;
      END
   END dout1[170]
   PIN dout1[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.8225 120.3225 289.9575 120.4575 ;
      END
   END dout1[171]
   PIN dout1[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.9975 120.3225 291.1325 120.4575 ;
      END
   END dout1[172]
   PIN dout1[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.1725 120.3225 292.3075 120.4575 ;
      END
   END dout1[173]
   PIN dout1[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.3475 120.3225 293.4825 120.4575 ;
      END
   END dout1[174]
   PIN dout1[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.5225 120.3225 294.6575 120.4575 ;
      END
   END dout1[175]
   PIN dout1[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.6975 120.3225 295.8325 120.4575 ;
      END
   END dout1[176]
   PIN dout1[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.8725 120.3225 297.0075 120.4575 ;
      END
   END dout1[177]
   PIN dout1[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.0475 120.3225 298.1825 120.4575 ;
      END
   END dout1[178]
   PIN dout1[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.2225 120.3225 299.3575 120.4575 ;
      END
   END dout1[179]
   PIN dout1[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.3975 120.3225 300.5325 120.4575 ;
      END
   END dout1[180]
   PIN dout1[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.5725 120.3225 301.7075 120.4575 ;
      END
   END dout1[181]
   PIN dout1[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  302.7475 120.3225 302.8825 120.4575 ;
      END
   END dout1[182]
   PIN dout1[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.9225 120.3225 304.0575 120.4575 ;
      END
   END dout1[183]
   PIN dout1[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.0975 120.3225 305.2325 120.4575 ;
      END
   END dout1[184]
   PIN dout1[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.2725 120.3225 306.4075 120.4575 ;
      END
   END dout1[185]
   PIN dout1[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.4475 120.3225 307.5825 120.4575 ;
      END
   END dout1[186]
   PIN dout1[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.6225 120.3225 308.7575 120.4575 ;
      END
   END dout1[187]
   PIN dout1[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.7975 120.3225 309.9325 120.4575 ;
      END
   END dout1[188]
   PIN dout1[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.9725 120.3225 311.1075 120.4575 ;
      END
   END dout1[189]
   PIN dout1[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.1475 120.3225 312.2825 120.4575 ;
      END
   END dout1[190]
   PIN dout1[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.3225 120.3225 313.4575 120.4575 ;
      END
   END dout1[191]
   PIN dout1[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.4975 120.3225 314.6325 120.4575 ;
      END
   END dout1[192]
   PIN dout1[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.6725 120.3225 315.8075 120.4575 ;
      END
   END dout1[193]
   PIN dout1[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.8475 120.3225 316.9825 120.4575 ;
      END
   END dout1[194]
   PIN dout1[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.0225 120.3225 318.1575 120.4575 ;
      END
   END dout1[195]
   PIN dout1[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.1975 120.3225 319.3325 120.4575 ;
      END
   END dout1[196]
   PIN dout1[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.3725 120.3225 320.5075 120.4575 ;
      END
   END dout1[197]
   PIN dout1[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.5475 120.3225 321.6825 120.4575 ;
      END
   END dout1[198]
   PIN dout1[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  322.7225 120.3225 322.8575 120.4575 ;
      END
   END dout1[199]
   PIN dout1[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.8975 120.3225 324.0325 120.4575 ;
      END
   END dout1[200]
   PIN dout1[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.0725 120.3225 325.2075 120.4575 ;
      END
   END dout1[201]
   PIN dout1[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.2475 120.3225 326.3825 120.4575 ;
      END
   END dout1[202]
   PIN dout1[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.4225 120.3225 327.5575 120.4575 ;
      END
   END dout1[203]
   PIN dout1[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.5975 120.3225 328.7325 120.4575 ;
      END
   END dout1[204]
   PIN dout1[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.7725 120.3225 329.9075 120.4575 ;
      END
   END dout1[205]
   PIN dout1[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.9475 120.3225 331.0825 120.4575 ;
      END
   END dout1[206]
   PIN dout1[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.1225 120.3225 332.2575 120.4575 ;
      END
   END dout1[207]
   PIN dout1[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.2975 120.3225 333.4325 120.4575 ;
      END
   END dout1[208]
   PIN dout1[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.4725 120.3225 334.6075 120.4575 ;
      END
   END dout1[209]
   PIN dout1[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.6475 120.3225 335.7825 120.4575 ;
      END
   END dout1[210]
   PIN dout1[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.8225 120.3225 336.9575 120.4575 ;
      END
   END dout1[211]
   PIN dout1[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.9975 120.3225 338.1325 120.4575 ;
      END
   END dout1[212]
   PIN dout1[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.1725 120.3225 339.3075 120.4575 ;
      END
   END dout1[213]
   PIN dout1[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.3475 120.3225 340.4825 120.4575 ;
      END
   END dout1[214]
   PIN dout1[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.5225 120.3225 341.6575 120.4575 ;
      END
   END dout1[215]
   PIN dout1[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.6975 120.3225 342.8325 120.4575 ;
      END
   END dout1[216]
   PIN dout1[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.8725 120.3225 344.0075 120.4575 ;
      END
   END dout1[217]
   PIN dout1[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.0475 120.3225 345.1825 120.4575 ;
      END
   END dout1[218]
   PIN dout1[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.2225 120.3225 346.3575 120.4575 ;
      END
   END dout1[219]
   PIN dout1[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.3975 120.3225 347.5325 120.4575 ;
      END
   END dout1[220]
   PIN dout1[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.5725 120.3225 348.7075 120.4575 ;
      END
   END dout1[221]
   PIN dout1[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.7475 120.3225 349.8825 120.4575 ;
      END
   END dout1[222]
   PIN dout1[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.9225 120.3225 351.0575 120.4575 ;
      END
   END dout1[223]
   PIN dout1[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.0975 120.3225 352.2325 120.4575 ;
      END
   END dout1[224]
   PIN dout1[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.2725 120.3225 353.4075 120.4575 ;
      END
   END dout1[225]
   PIN dout1[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.4475 120.3225 354.5825 120.4575 ;
      END
   END dout1[226]
   PIN dout1[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.6225 120.3225 355.7575 120.4575 ;
      END
   END dout1[227]
   PIN dout1[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.7975 120.3225 356.9325 120.4575 ;
      END
   END dout1[228]
   PIN dout1[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.9725 120.3225 358.1075 120.4575 ;
      END
   END dout1[229]
   PIN dout1[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.1475 120.3225 359.2825 120.4575 ;
      END
   END dout1[230]
   PIN dout1[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.3225 120.3225 360.4575 120.4575 ;
      END
   END dout1[231]
   PIN dout1[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.4975 120.3225 361.6325 120.4575 ;
      END
   END dout1[232]
   PIN dout1[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.6725 120.3225 362.8075 120.4575 ;
      END
   END dout1[233]
   PIN dout1[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.8475 120.3225 363.9825 120.4575 ;
      END
   END dout1[234]
   PIN dout1[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.0225 120.3225 365.1575 120.4575 ;
      END
   END dout1[235]
   PIN dout1[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.1975 120.3225 366.3325 120.4575 ;
      END
   END dout1[236]
   PIN dout1[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.3725 120.3225 367.5075 120.4575 ;
      END
   END dout1[237]
   PIN dout1[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.5475 120.3225 368.6825 120.4575 ;
      END
   END dout1[238]
   PIN dout1[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.7225 120.3225 369.8575 120.4575 ;
      END
   END dout1[239]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  374.075 47.1425 374.215 113.1725 ;
         LAYER metal4 ;
         RECT  459.3675 96.0225 459.5075 118.425 ;
         LAYER metal3 ;
         RECT  661.1875 2.47 661.3225 2.605 ;
         LAYER metal3 ;
         RECT  66.6875 69.75 66.8225 69.885 ;
         LAYER metal3 ;
         RECT  393.0375 63.77 393.1725 63.905 ;
         LAYER metal3 ;
         RECT  638.3075 2.47 638.4425 2.605 ;
         LAYER metal3 ;
         RECT  523.9075 2.47 524.0425 2.605 ;
         LAYER metal3 ;
         RECT  146.3875 2.47 146.5225 2.605 ;
         LAYER metal4 ;
         RECT  387.48 50.3125 387.62 110.3225 ;
         LAYER metal3 ;
         RECT  66.6875 54.8 66.8225 54.935 ;
         LAYER metal3 ;
         RECT  352.3075 2.47 352.4425 2.605 ;
         LAYER metal3 ;
         RECT  501.0275 2.47 501.1625 2.605 ;
         LAYER metal3 ;
         RECT  169.2675 2.47 169.4025 2.605 ;
         LAYER metal3 ;
         RECT  393.0375 60.78 393.1725 60.915 ;
         LAYER metal3 ;
         RECT  457.635 125.665 457.77 125.8 ;
         LAYER metal3 ;
         RECT  569.6675 2.47 569.8025 2.605 ;
         LAYER metal4 ;
         RECT  396.61 115.7825 396.75 125.8025 ;
         LAYER metal3 ;
         RECT  72.86 49.6075 72.995 49.7425 ;
         LAYER metal4 ;
         RECT  60.585 74.2325 60.725 89.1925 ;
         LAYER metal3 ;
         RECT  66.6875 60.78 66.8225 60.915 ;
         LAYER metal3 ;
         RECT  112.0675 2.47 112.2025 2.605 ;
         LAYER metal3 ;
         RECT  295.1075 2.47 295.2425 2.605 ;
         LAYER metal4 ;
         RECT  72.24 50.3125 72.38 110.3225 ;
         LAYER metal3 ;
         RECT  66.3075 2.47 66.4425 2.605 ;
         LAYER metal3 ;
         RECT  512.4675 2.47 512.6025 2.605 ;
         LAYER metal3 ;
         RECT  85.7125 46.4475 370.9975 46.5175 ;
         LAYER metal3 ;
         RECT  649.7475 2.47 649.8825 2.605 ;
         LAYER metal3 ;
         RECT  489.5875 2.47 489.7225 2.605 ;
         LAYER metal3 ;
         RECT  272.2275 2.47 272.3625 2.605 ;
         LAYER metal3 ;
         RECT  393.0375 72.74 393.1725 72.875 ;
         LAYER metal3 ;
         RECT  203.5875 2.47 203.7225 2.605 ;
         LAYER metal3 ;
         RECT  85.7125 117.765 370.5275 117.835 ;
         LAYER metal3 ;
         RECT  66.6875 51.81 66.8225 51.945 ;
         LAYER metal3 ;
         RECT  592.5475 2.47 592.6825 2.605 ;
         LAYER metal3 ;
         RECT  386.6275 2.47 386.7625 2.605 ;
         LAYER metal3 ;
         RECT  466.7075 2.47 466.8425 2.605 ;
         LAYER metal3 ;
         RECT  741.2675 2.47 741.4025 2.605 ;
         LAYER metal3 ;
         RECT  85.7125 41.0125 370.5275 41.0825 ;
         LAYER metal3 ;
         RECT  626.8675 2.47 627.0025 2.605 ;
         LAYER metal4 ;
         RECT  375.155 50.3125 375.295 110.2525 ;
         LAYER metal3 ;
         RECT  157.8275 2.47 157.9625 2.605 ;
         LAYER metal3 ;
         RECT  89.1875 2.47 89.3225 2.605 ;
         LAYER metal3 ;
         RECT  393.0375 69.75 393.1725 69.885 ;
         LAYER metal3 ;
         RECT  329.4275 2.47 329.5625 2.605 ;
         LAYER metal3 ;
         RECT  535.3475 2.47 535.4825 2.605 ;
         LAYER metal3 ;
         RECT  398.0675 2.47 398.2025 2.605 ;
         LAYER metal3 ;
         RECT  134.9475 2.47 135.0825 2.605 ;
         LAYER metal3 ;
         RECT  603.9875 2.47 604.1225 2.605 ;
         LAYER metal3 ;
         RECT  386.865 110.8225 387.0 110.9575 ;
         LAYER metal3 ;
         RECT  455.2675 2.47 455.4025 2.605 ;
         LAYER metal3 ;
         RECT  478.1475 2.47 478.2825 2.605 ;
         LAYER metal3 ;
         RECT  237.9075 2.47 238.0425 2.605 ;
         LAYER metal3 ;
         RECT  249.3475 2.47 249.4825 2.605 ;
         LAYER metal3 ;
         RECT  340.8675 2.47 341.0025 2.605 ;
         LAYER metal4 ;
         RECT  63.305 32.1125 63.445 47.0725 ;
         LAYER metal3 ;
         RECT  375.1875 2.47 375.3225 2.605 ;
         LAYER metal3 ;
         RECT  260.7875 2.47 260.9225 2.605 ;
         LAYER metal4 ;
         RECT  84.565 50.3125 84.705 110.2525 ;
         LAYER metal3 ;
         RECT  432.3875 2.47 432.5225 2.605 ;
         LAYER metal3 ;
         RECT  317.9875 2.47 318.1225 2.605 ;
         LAYER metal3 ;
         RECT  226.4675 2.47 226.6025 2.605 ;
         LAYER metal3 ;
         RECT  85.7125 113.8675 372.1725 113.9375 ;
         LAYER metal3 ;
         RECT  283.6675 2.47 283.8025 2.605 ;
         LAYER metal3 ;
         RECT  684.0675 2.47 684.2025 2.605 ;
         LAYER metal3 ;
         RECT  581.1075 2.47 581.2425 2.605 ;
         LAYER metal3 ;
         RECT  729.8275 2.47 729.9625 2.605 ;
         LAYER metal3 ;
         RECT  558.2275 2.47 558.3625 2.605 ;
         LAYER metal3 ;
         RECT  615.4275 2.47 615.5625 2.605 ;
         LAYER metal3 ;
         RECT  718.3875 2.47 718.5225 2.605 ;
         LAYER metal3 ;
         RECT  2.425 32.115 2.56 32.25 ;
         LAYER metal3 ;
         RECT  66.6875 72.74 66.8225 72.875 ;
         LAYER metal3 ;
         RECT  215.0275 2.47 215.1625 2.605 ;
         LAYER metal3 ;
         RECT  77.7475 2.47 77.8825 2.605 ;
         LAYER metal3 ;
         RECT  672.6275 2.47 672.7625 2.605 ;
         LAYER metal3 ;
         RECT  306.5475 2.47 306.6825 2.605 ;
         LAYER metal3 ;
         RECT  393.0375 54.8 393.1725 54.935 ;
         LAYER metal3 ;
         RECT  100.6275 2.47 100.7625 2.605 ;
         LAYER metal3 ;
         RECT  123.5075 2.47 123.6425 2.605 ;
         LAYER metal3 ;
         RECT  695.5075 2.47 695.6425 2.605 ;
         LAYER metal3 ;
         RECT  192.1475 2.47 192.2825 2.605 ;
         LAYER metal3 ;
         RECT  420.9475 2.47 421.0825 2.605 ;
         LAYER metal3 ;
         RECT  84.5675 48.82 84.7025 48.955 ;
         LAYER metal4 ;
         RECT  85.645 47.1425 85.785 113.1725 ;
         LAYER metal3 ;
         RECT  409.5075 2.47 409.6425 2.605 ;
         LAYER metal3 ;
         RECT  443.8275 2.47 443.9625 2.605 ;
         LAYER metal3 ;
         RECT  546.7875 2.47 546.9225 2.605 ;
         LAYER metal4 ;
         RECT  399.33 35.4925 399.47 50.4525 ;
         LAYER metal4 ;
         RECT  0.6875 39.49 0.8275 61.8925 ;
         LAYER metal3 ;
         RECT  66.6875 63.77 66.8225 63.905 ;
         LAYER metal3 ;
         RECT  706.9475 2.47 707.0825 2.605 ;
         LAYER metal3 ;
         RECT  363.7475 2.47 363.8825 2.605 ;
         LAYER metal3 ;
         RECT  180.7075 2.47 180.8425 2.605 ;
         LAYER metal3 ;
         RECT  393.0375 51.81 393.1725 51.945 ;
         LAYER metal3 ;
         RECT  375.1575 111.61 375.2925 111.745 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  320.8475 0.0 320.9825 0.135 ;
         LAYER metal3 ;
         RECT  309.4075 0.0 309.5425 0.135 ;
         LAYER metal3 ;
         RECT  412.3675 0.0 412.5025 0.135 ;
         LAYER metal3 ;
         RECT  65.16 53.305 65.295 53.44 ;
         LAYER metal4 ;
         RECT  453.81 113.3125 453.95 128.2725 ;
         LAYER metal3 ;
         RECT  85.7125 43.0625 370.5275 43.1325 ;
         LAYER metal3 ;
         RECT  394.565 74.235 394.7 74.37 ;
         LAYER metal4 ;
         RECT  63.445 74.1675 63.585 89.2575 ;
         LAYER metal3 ;
         RECT  394.565 56.295 394.7 56.43 ;
         LAYER metal3 ;
         RECT  538.2075 0.0 538.3425 0.135 ;
         LAYER metal3 ;
         RECT  80.6075 0.0 80.7425 0.135 ;
         LAYER metal3 ;
         RECT  492.4475 0.0 492.5825 0.135 ;
         LAYER metal3 ;
         RECT  572.5275 0.0 572.6625 0.135 ;
         LAYER metal3 ;
         RECT  721.2475 0.0 721.3825 0.135 ;
         LAYER metal3 ;
         RECT  65.16 74.235 65.295 74.37 ;
         LAYER metal3 ;
         RECT  172.1275 0.0 172.2625 0.135 ;
         LAYER metal3 ;
         RECT  458.1275 0.0 458.2625 0.135 ;
         LAYER metal3 ;
         RECT  732.6875 0.0 732.8225 0.135 ;
         LAYER metal4 ;
         RECT  6.105 29.6425 6.245 44.6025 ;
         LAYER metal3 ;
         RECT  446.6875 0.0 446.8225 0.135 ;
         LAYER metal4 ;
         RECT  70.305 50.28 70.445 110.3225 ;
         LAYER metal3 ;
         RECT  217.8875 0.0 218.0225 0.135 ;
         LAYER metal3 ;
         RECT  394.565 59.285 394.7 59.42 ;
         LAYER metal3 ;
         RECT  65.16 56.295 65.295 56.43 ;
         LAYER metal3 ;
         RECT  664.0475 0.0 664.1825 0.135 ;
         LAYER metal3 ;
         RECT  423.8075 0.0 423.9425 0.135 ;
         LAYER metal3 ;
         RECT  394.565 50.315 394.7 50.45 ;
         LAYER metal4 ;
         RECT  389.415 50.28 389.555 110.3225 ;
         LAYER metal3 ;
         RECT  709.8075 0.0 709.9425 0.135 ;
         LAYER metal3 ;
         RECT  126.3675 0.0 126.5025 0.135 ;
         LAYER metal3 ;
         RECT  229.3275 0.0 229.4625 0.135 ;
         LAYER metal3 ;
         RECT  394.565 53.305 394.7 53.44 ;
         LAYER metal3 ;
         RECT  92.0475 0.0 92.1825 0.135 ;
         LAYER metal3 ;
         RECT  515.3275 0.0 515.4625 0.135 ;
         LAYER metal3 ;
         RECT  2.425 29.645 2.56 29.78 ;
         LAYER metal3 ;
         RECT  457.635 128.135 457.77 128.27 ;
         LAYER metal3 ;
         RECT  606.8475 0.0 606.9825 0.135 ;
         LAYER metal3 ;
         RECT  675.4875 0.0 675.6225 0.135 ;
         LAYER metal4 ;
         RECT  396.47 35.4275 396.61 50.5175 ;
         LAYER metal3 ;
         RECT  65.16 50.315 65.295 50.45 ;
         LAYER metal3 ;
         RECT  149.2475 0.0 149.3825 0.135 ;
         LAYER metal3 ;
         RECT  332.2875 0.0 332.4225 0.135 ;
         LAYER metal3 ;
         RECT  183.5675 0.0 183.7025 0.135 ;
         LAYER metal3 ;
         RECT  206.4475 0.0 206.5825 0.135 ;
         LAYER metal4 ;
         RECT  457.305 95.99 457.445 118.3925 ;
         LAYER metal3 ;
         RECT  595.4075 0.0 595.5425 0.135 ;
         LAYER metal3 ;
         RECT  394.565 65.265 394.7 65.4 ;
         LAYER metal3 ;
         RECT  69.1675 0.0 69.3025 0.135 ;
         LAYER metal3 ;
         RECT  275.0875 0.0 275.2225 0.135 ;
         LAYER metal3 ;
         RECT  137.8075 0.0 137.9425 0.135 ;
         LAYER metal3 ;
         RECT  503.8875 0.0 504.0225 0.135 ;
         LAYER metal3 ;
         RECT  652.6075 0.0 652.7425 0.135 ;
         LAYER metal4 ;
         RECT  386.92 50.28 387.06 110.285 ;
         LAYER metal3 ;
         RECT  394.565 68.255 394.7 68.39 ;
         LAYER metal3 ;
         RECT  698.3675 0.0 698.5025 0.135 ;
         LAYER metal4 ;
         RECT  2.75 39.5225 2.89 61.925 ;
         LAYER metal3 ;
         RECT  469.5675 0.0 469.7025 0.135 ;
         LAYER metal4 ;
         RECT  72.8 50.28 72.94 110.285 ;
         LAYER metal3 ;
         RECT  583.9675 0.0 584.1025 0.135 ;
         LAYER metal3 ;
         RECT  561.0875 0.0 561.2225 0.135 ;
         LAYER metal3 ;
         RECT  435.2475 0.0 435.3825 0.135 ;
         LAYER metal3 ;
         RECT  744.1275 0.0 744.2625 0.135 ;
         LAYER metal3 ;
         RECT  195.0075 0.0 195.1425 0.135 ;
         LAYER metal3 ;
         RECT  65.16 62.275 65.295 62.41 ;
         LAYER metal3 ;
         RECT  252.2075 0.0 252.3425 0.135 ;
         LAYER metal4 ;
         RECT  373.615 47.1425 373.755 113.1725 ;
         LAYER metal3 ;
         RECT  114.9275 0.0 115.0625 0.135 ;
         LAYER metal3 ;
         RECT  160.6875 0.0 160.8225 0.135 ;
         LAYER metal3 ;
         RECT  686.9275 0.0 687.0625 0.135 ;
         LAYER metal3 ;
         RECT  85.7125 115.8725 370.5625 115.9425 ;
         LAYER metal3 ;
         RECT  629.7275 0.0 629.8625 0.135 ;
         LAYER metal3 ;
         RECT  65.16 65.265 65.295 65.4 ;
         LAYER metal3 ;
         RECT  240.7675 0.0 240.9025 0.135 ;
         LAYER metal3 ;
         RECT  641.1675 0.0 641.3025 0.135 ;
         LAYER metal3 ;
         RECT  286.5275 0.0 286.6625 0.135 ;
         LAYER metal3 ;
         RECT  355.1675 0.0 355.3025 0.135 ;
         LAYER metal3 ;
         RECT  65.16 59.285 65.295 59.42 ;
         LAYER metal3 ;
         RECT  389.4875 0.0 389.6225 0.135 ;
         LAYER metal3 ;
         RECT  103.4875 0.0 103.6225 0.135 ;
         LAYER metal3 ;
         RECT  394.565 62.275 394.7 62.41 ;
         LAYER metal3 ;
         RECT  481.0075 0.0 481.1425 0.135 ;
         LAYER metal3 ;
         RECT  65.16 68.255 65.295 68.39 ;
         LAYER metal3 ;
         RECT  526.7675 0.0 526.9025 0.135 ;
         LAYER metal3 ;
         RECT  400.9275 0.0 401.0625 0.135 ;
         LAYER metal3 ;
         RECT  366.6075 0.0 366.7425 0.135 ;
         LAYER metal3 ;
         RECT  618.2875 0.0 618.4225 0.135 ;
         LAYER metal3 ;
         RECT  343.7275 0.0 343.8625 0.135 ;
         LAYER metal3 ;
         RECT  263.6475 0.0 263.7825 0.135 ;
         LAYER metal3 ;
         RECT  378.0475 0.0 378.1825 0.135 ;
         LAYER metal4 ;
         RECT  86.105 47.1425 86.245 113.1725 ;
         LAYER metal3 ;
         RECT  297.9675 0.0 298.1025 0.135 ;
         LAYER metal3 ;
         RECT  549.6475 0.0 549.7825 0.135 ;
         LAYER metal3 ;
         RECT  65.16 71.245 65.295 71.38 ;
         LAYER metal3 ;
         RECT  394.565 71.245 394.7 71.38 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 752.635 128.1325 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 752.635 128.1325 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 66.45 0.965 ;
      RECT  0.14 0.965 66.45 1.38 ;
      RECT  66.45 0.14 66.865 0.965 ;
      RECT  66.865 0.965 69.31 1.38 ;
      RECT  69.725 0.965 72.17 1.38 ;
      RECT  72.585 0.965 75.03 1.38 ;
      RECT  75.445 0.965 77.89 1.38 ;
      RECT  78.305 0.965 80.75 1.38 ;
      RECT  81.165 0.965 83.61 1.38 ;
      RECT  84.025 0.965 86.47 1.38 ;
      RECT  86.885 0.965 89.33 1.38 ;
      RECT  89.745 0.965 92.19 1.38 ;
      RECT  92.605 0.965 95.05 1.38 ;
      RECT  95.465 0.965 97.91 1.38 ;
      RECT  98.325 0.965 100.77 1.38 ;
      RECT  101.185 0.965 103.63 1.38 ;
      RECT  104.045 0.965 106.49 1.38 ;
      RECT  106.905 0.965 109.35 1.38 ;
      RECT  109.765 0.965 112.21 1.38 ;
      RECT  112.625 0.965 115.07 1.38 ;
      RECT  115.485 0.965 117.93 1.38 ;
      RECT  118.345 0.965 120.79 1.38 ;
      RECT  121.205 0.965 123.65 1.38 ;
      RECT  124.065 0.965 126.51 1.38 ;
      RECT  126.925 0.965 129.37 1.38 ;
      RECT  129.785 0.965 132.23 1.38 ;
      RECT  132.645 0.965 135.09 1.38 ;
      RECT  135.505 0.965 137.95 1.38 ;
      RECT  138.365 0.965 140.81 1.38 ;
      RECT  141.225 0.965 143.67 1.38 ;
      RECT  144.085 0.965 146.53 1.38 ;
      RECT  146.945 0.965 149.39 1.38 ;
      RECT  149.805 0.965 152.25 1.38 ;
      RECT  152.665 0.965 155.11 1.38 ;
      RECT  155.525 0.965 157.97 1.38 ;
      RECT  158.385 0.965 160.83 1.38 ;
      RECT  161.245 0.965 163.69 1.38 ;
      RECT  164.105 0.965 166.55 1.38 ;
      RECT  166.965 0.965 169.41 1.38 ;
      RECT  169.825 0.965 172.27 1.38 ;
      RECT  172.685 0.965 175.13 1.38 ;
      RECT  175.545 0.965 177.99 1.38 ;
      RECT  178.405 0.965 180.85 1.38 ;
      RECT  181.265 0.965 183.71 1.38 ;
      RECT  184.125 0.965 186.57 1.38 ;
      RECT  186.985 0.965 189.43 1.38 ;
      RECT  189.845 0.965 192.29 1.38 ;
      RECT  192.705 0.965 195.15 1.38 ;
      RECT  195.565 0.965 198.01 1.38 ;
      RECT  198.425 0.965 200.87 1.38 ;
      RECT  201.285 0.965 203.73 1.38 ;
      RECT  204.145 0.965 206.59 1.38 ;
      RECT  207.005 0.965 209.45 1.38 ;
      RECT  209.865 0.965 212.31 1.38 ;
      RECT  212.725 0.965 215.17 1.38 ;
      RECT  215.585 0.965 218.03 1.38 ;
      RECT  218.445 0.965 220.89 1.38 ;
      RECT  221.305 0.965 223.75 1.38 ;
      RECT  224.165 0.965 226.61 1.38 ;
      RECT  227.025 0.965 229.47 1.38 ;
      RECT  229.885 0.965 232.33 1.38 ;
      RECT  232.745 0.965 235.19 1.38 ;
      RECT  235.605 0.965 238.05 1.38 ;
      RECT  238.465 0.965 240.91 1.38 ;
      RECT  241.325 0.965 243.77 1.38 ;
      RECT  244.185 0.965 246.63 1.38 ;
      RECT  247.045 0.965 249.49 1.38 ;
      RECT  249.905 0.965 252.35 1.38 ;
      RECT  252.765 0.965 255.21 1.38 ;
      RECT  255.625 0.965 258.07 1.38 ;
      RECT  258.485 0.965 260.93 1.38 ;
      RECT  261.345 0.965 263.79 1.38 ;
      RECT  264.205 0.965 266.65 1.38 ;
      RECT  267.065 0.965 269.51 1.38 ;
      RECT  269.925 0.965 272.37 1.38 ;
      RECT  272.785 0.965 275.23 1.38 ;
      RECT  275.645 0.965 278.09 1.38 ;
      RECT  278.505 0.965 280.95 1.38 ;
      RECT  281.365 0.965 283.81 1.38 ;
      RECT  284.225 0.965 286.67 1.38 ;
      RECT  287.085 0.965 289.53 1.38 ;
      RECT  289.945 0.965 292.39 1.38 ;
      RECT  292.805 0.965 295.25 1.38 ;
      RECT  295.665 0.965 298.11 1.38 ;
      RECT  298.525 0.965 300.97 1.38 ;
      RECT  301.385 0.965 303.83 1.38 ;
      RECT  304.245 0.965 306.69 1.38 ;
      RECT  307.105 0.965 309.55 1.38 ;
      RECT  309.965 0.965 312.41 1.38 ;
      RECT  312.825 0.965 315.27 1.38 ;
      RECT  315.685 0.965 318.13 1.38 ;
      RECT  318.545 0.965 320.99 1.38 ;
      RECT  321.405 0.965 323.85 1.38 ;
      RECT  324.265 0.965 326.71 1.38 ;
      RECT  327.125 0.965 329.57 1.38 ;
      RECT  329.985 0.965 332.43 1.38 ;
      RECT  332.845 0.965 335.29 1.38 ;
      RECT  335.705 0.965 338.15 1.38 ;
      RECT  338.565 0.965 341.01 1.38 ;
      RECT  341.425 0.965 343.87 1.38 ;
      RECT  344.285 0.965 346.73 1.38 ;
      RECT  347.145 0.965 349.59 1.38 ;
      RECT  350.005 0.965 352.45 1.38 ;
      RECT  352.865 0.965 355.31 1.38 ;
      RECT  355.725 0.965 358.17 1.38 ;
      RECT  358.585 0.965 361.03 1.38 ;
      RECT  361.445 0.965 363.89 1.38 ;
      RECT  364.305 0.965 366.75 1.38 ;
      RECT  367.165 0.965 369.61 1.38 ;
      RECT  370.025 0.965 372.47 1.38 ;
      RECT  372.885 0.965 375.33 1.38 ;
      RECT  375.745 0.965 378.19 1.38 ;
      RECT  378.605 0.965 381.05 1.38 ;
      RECT  381.465 0.965 383.91 1.38 ;
      RECT  384.325 0.965 386.77 1.38 ;
      RECT  387.185 0.965 389.63 1.38 ;
      RECT  390.045 0.965 392.49 1.38 ;
      RECT  392.905 0.965 395.35 1.38 ;
      RECT  395.765 0.965 398.21 1.38 ;
      RECT  398.625 0.965 401.07 1.38 ;
      RECT  401.485 0.965 403.93 1.38 ;
      RECT  404.345 0.965 406.79 1.38 ;
      RECT  407.205 0.965 409.65 1.38 ;
      RECT  410.065 0.965 412.51 1.38 ;
      RECT  412.925 0.965 415.37 1.38 ;
      RECT  415.785 0.965 418.23 1.38 ;
      RECT  418.645 0.965 421.09 1.38 ;
      RECT  421.505 0.965 423.95 1.38 ;
      RECT  424.365 0.965 426.81 1.38 ;
      RECT  427.225 0.965 429.67 1.38 ;
      RECT  430.085 0.965 432.53 1.38 ;
      RECT  432.945 0.965 435.39 1.38 ;
      RECT  435.805 0.965 438.25 1.38 ;
      RECT  438.665 0.965 441.11 1.38 ;
      RECT  441.525 0.965 443.97 1.38 ;
      RECT  444.385 0.965 446.83 1.38 ;
      RECT  447.245 0.965 449.69 1.38 ;
      RECT  450.105 0.965 452.55 1.38 ;
      RECT  452.965 0.965 455.41 1.38 ;
      RECT  455.825 0.965 458.27 1.38 ;
      RECT  458.685 0.965 461.13 1.38 ;
      RECT  461.545 0.965 463.99 1.38 ;
      RECT  464.405 0.965 466.85 1.38 ;
      RECT  467.265 0.965 469.71 1.38 ;
      RECT  470.125 0.965 472.57 1.38 ;
      RECT  472.985 0.965 475.43 1.38 ;
      RECT  475.845 0.965 478.29 1.38 ;
      RECT  478.705 0.965 481.15 1.38 ;
      RECT  481.565 0.965 484.01 1.38 ;
      RECT  484.425 0.965 486.87 1.38 ;
      RECT  487.285 0.965 489.73 1.38 ;
      RECT  490.145 0.965 492.59 1.38 ;
      RECT  493.005 0.965 495.45 1.38 ;
      RECT  495.865 0.965 498.31 1.38 ;
      RECT  498.725 0.965 501.17 1.38 ;
      RECT  501.585 0.965 504.03 1.38 ;
      RECT  504.445 0.965 506.89 1.38 ;
      RECT  507.305 0.965 509.75 1.38 ;
      RECT  510.165 0.965 512.61 1.38 ;
      RECT  513.025 0.965 515.47 1.38 ;
      RECT  515.885 0.965 518.33 1.38 ;
      RECT  518.745 0.965 521.19 1.38 ;
      RECT  521.605 0.965 524.05 1.38 ;
      RECT  524.465 0.965 526.91 1.38 ;
      RECT  527.325 0.965 529.77 1.38 ;
      RECT  530.185 0.965 532.63 1.38 ;
      RECT  533.045 0.965 535.49 1.38 ;
      RECT  535.905 0.965 538.35 1.38 ;
      RECT  538.765 0.965 541.21 1.38 ;
      RECT  541.625 0.965 544.07 1.38 ;
      RECT  544.485 0.965 546.93 1.38 ;
      RECT  547.345 0.965 549.79 1.38 ;
      RECT  550.205 0.965 552.65 1.38 ;
      RECT  553.065 0.965 555.51 1.38 ;
      RECT  555.925 0.965 558.37 1.38 ;
      RECT  558.785 0.965 561.23 1.38 ;
      RECT  561.645 0.965 564.09 1.38 ;
      RECT  564.505 0.965 566.95 1.38 ;
      RECT  567.365 0.965 569.81 1.38 ;
      RECT  570.225 0.965 572.67 1.38 ;
      RECT  573.085 0.965 575.53 1.38 ;
      RECT  575.945 0.965 578.39 1.38 ;
      RECT  578.805 0.965 581.25 1.38 ;
      RECT  581.665 0.965 584.11 1.38 ;
      RECT  584.525 0.965 586.97 1.38 ;
      RECT  587.385 0.965 589.83 1.38 ;
      RECT  590.245 0.965 592.69 1.38 ;
      RECT  593.105 0.965 595.55 1.38 ;
      RECT  595.965 0.965 598.41 1.38 ;
      RECT  598.825 0.965 601.27 1.38 ;
      RECT  601.685 0.965 604.13 1.38 ;
      RECT  604.545 0.965 606.99 1.38 ;
      RECT  607.405 0.965 609.85 1.38 ;
      RECT  610.265 0.965 612.71 1.38 ;
      RECT  613.125 0.965 615.57 1.38 ;
      RECT  615.985 0.965 618.43 1.38 ;
      RECT  618.845 0.965 621.29 1.38 ;
      RECT  621.705 0.965 624.15 1.38 ;
      RECT  624.565 0.965 627.01 1.38 ;
      RECT  627.425 0.965 629.87 1.38 ;
      RECT  630.285 0.965 632.73 1.38 ;
      RECT  633.145 0.965 635.59 1.38 ;
      RECT  636.005 0.965 638.45 1.38 ;
      RECT  638.865 0.965 641.31 1.38 ;
      RECT  641.725 0.965 644.17 1.38 ;
      RECT  644.585 0.965 647.03 1.38 ;
      RECT  647.445 0.965 649.89 1.38 ;
      RECT  650.305 0.965 652.75 1.38 ;
      RECT  653.165 0.965 655.61 1.38 ;
      RECT  656.025 0.965 658.47 1.38 ;
      RECT  658.885 0.965 661.33 1.38 ;
      RECT  661.745 0.965 664.19 1.38 ;
      RECT  664.605 0.965 667.05 1.38 ;
      RECT  667.465 0.965 669.91 1.38 ;
      RECT  670.325 0.965 672.77 1.38 ;
      RECT  673.185 0.965 675.63 1.38 ;
      RECT  676.045 0.965 678.49 1.38 ;
      RECT  678.905 0.965 681.35 1.38 ;
      RECT  681.765 0.965 684.21 1.38 ;
      RECT  684.625 0.965 687.07 1.38 ;
      RECT  687.485 0.965 689.93 1.38 ;
      RECT  690.345 0.965 692.79 1.38 ;
      RECT  693.205 0.965 695.65 1.38 ;
      RECT  696.065 0.965 698.51 1.38 ;
      RECT  698.925 0.965 701.37 1.38 ;
      RECT  701.785 0.965 704.23 1.38 ;
      RECT  704.645 0.965 707.09 1.38 ;
      RECT  707.505 0.965 709.95 1.38 ;
      RECT  710.365 0.965 712.81 1.38 ;
      RECT  713.225 0.965 715.67 1.38 ;
      RECT  716.085 0.965 718.53 1.38 ;
      RECT  718.945 0.965 721.39 1.38 ;
      RECT  721.805 0.965 724.25 1.38 ;
      RECT  724.665 0.965 727.11 1.38 ;
      RECT  727.525 0.965 729.97 1.38 ;
      RECT  730.385 0.965 732.83 1.38 ;
      RECT  733.245 0.965 735.69 1.38 ;
      RECT  736.105 0.965 738.55 1.38 ;
      RECT  738.965 0.965 741.41 1.38 ;
      RECT  741.825 0.965 744.27 1.38 ;
      RECT  744.685 0.965 747.13 1.38 ;
      RECT  747.545 0.965 749.99 1.38 ;
      RECT  750.405 0.965 752.635 1.38 ;
      RECT  0.14 75.2 60.73 75.615 ;
      RECT  0.14 75.615 60.73 128.1325 ;
      RECT  60.73 1.38 61.145 75.2 ;
      RECT  61.145 75.2 66.45 75.615 ;
      RECT  61.145 75.615 66.45 128.1325 ;
      RECT  60.73 75.615 61.145 77.93 ;
      RECT  60.73 78.345 61.145 80.14 ;
      RECT  60.73 80.555 61.145 82.87 ;
      RECT  60.73 83.285 61.145 85.08 ;
      RECT  60.73 85.495 61.145 87.81 ;
      RECT  60.73 88.225 61.145 128.1325 ;
      RECT  398.91 49.485 399.325 128.1325 ;
      RECT  399.325 49.07 752.635 49.485 ;
      RECT  398.91 46.755 399.325 49.07 ;
      RECT  398.91 44.545 399.325 46.34 ;
      RECT  398.91 41.815 399.325 44.13 ;
      RECT  398.91 39.605 399.325 41.4 ;
      RECT  398.91 1.38 399.325 36.46 ;
      RECT  398.91 36.875 399.325 39.19 ;
      RECT  0.14 1.38 0.145 30.61 ;
      RECT  0.14 30.61 0.145 31.025 ;
      RECT  0.14 31.025 0.145 75.2 ;
      RECT  0.145 1.38 0.56 30.61 ;
      RECT  0.145 31.025 0.56 75.2 ;
      RECT  459.635 49.485 460.05 126.89 ;
      RECT  459.635 127.305 460.05 128.1325 ;
      RECT  460.05 49.485 752.635 126.89 ;
      RECT  460.05 126.89 752.635 127.305 ;
      RECT  460.05 127.305 752.635 128.1325 ;
      RECT  0.56 30.61 6.1075 30.695 ;
      RECT  0.56 30.695 6.1075 31.025 ;
      RECT  6.1075 30.61 6.5225 30.695 ;
      RECT  6.5225 30.61 60.73 30.695 ;
      RECT  6.5225 30.695 60.73 31.025 ;
      RECT  0.56 31.025 6.1075 31.11 ;
      RECT  6.1075 31.11 6.5225 75.2 ;
      RECT  6.5225 31.025 60.73 31.11 ;
      RECT  6.5225 31.11 60.73 75.2 ;
      RECT  399.325 49.485 453.5325 126.805 ;
      RECT  399.325 126.805 453.5325 126.89 ;
      RECT  453.5325 49.485 453.9475 126.805 ;
      RECT  453.9475 126.805 459.635 126.89 ;
      RECT  399.325 126.89 453.5325 127.22 ;
      RECT  399.325 127.22 453.5325 127.305 ;
      RECT  453.5325 127.22 453.9475 127.305 ;
      RECT  453.9475 126.89 459.635 127.22 ;
      RECT  453.9475 127.22 459.635 127.305 ;
      RECT  66.865 120.1825 88.7575 120.5975 ;
      RECT  66.865 120.5975 88.7575 128.1325 ;
      RECT  88.7575 120.5975 89.1725 128.1325 ;
      RECT  89.1725 120.5975 398.91 128.1325 ;
      RECT  89.1725 120.1825 89.9325 120.5975 ;
      RECT  90.3475 120.1825 91.1075 120.5975 ;
      RECT  91.5225 120.1825 92.2825 120.5975 ;
      RECT  92.6975 120.1825 93.4575 120.5975 ;
      RECT  93.8725 120.1825 94.6325 120.5975 ;
      RECT  95.0475 120.1825 95.8075 120.5975 ;
      RECT  96.2225 120.1825 96.9825 120.5975 ;
      RECT  97.3975 120.1825 98.1575 120.5975 ;
      RECT  98.5725 120.1825 99.3325 120.5975 ;
      RECT  99.7475 120.1825 100.5075 120.5975 ;
      RECT  100.9225 120.1825 101.6825 120.5975 ;
      RECT  102.0975 120.1825 102.8575 120.5975 ;
      RECT  103.2725 120.1825 104.0325 120.5975 ;
      RECT  104.4475 120.1825 105.2075 120.5975 ;
      RECT  105.6225 120.1825 106.3825 120.5975 ;
      RECT  106.7975 120.1825 107.5575 120.5975 ;
      RECT  107.9725 120.1825 108.7325 120.5975 ;
      RECT  109.1475 120.1825 109.9075 120.5975 ;
      RECT  110.3225 120.1825 111.0825 120.5975 ;
      RECT  111.4975 120.1825 112.2575 120.5975 ;
      RECT  112.6725 120.1825 113.4325 120.5975 ;
      RECT  113.8475 120.1825 114.6075 120.5975 ;
      RECT  115.0225 120.1825 115.7825 120.5975 ;
      RECT  116.1975 120.1825 116.9575 120.5975 ;
      RECT  117.3725 120.1825 118.1325 120.5975 ;
      RECT  118.5475 120.1825 119.3075 120.5975 ;
      RECT  119.7225 120.1825 120.4825 120.5975 ;
      RECT  120.8975 120.1825 121.6575 120.5975 ;
      RECT  122.0725 120.1825 122.8325 120.5975 ;
      RECT  123.2475 120.1825 124.0075 120.5975 ;
      RECT  124.4225 120.1825 125.1825 120.5975 ;
      RECT  125.5975 120.1825 126.3575 120.5975 ;
      RECT  126.7725 120.1825 127.5325 120.5975 ;
      RECT  127.9475 120.1825 128.7075 120.5975 ;
      RECT  129.1225 120.1825 129.8825 120.5975 ;
      RECT  130.2975 120.1825 131.0575 120.5975 ;
      RECT  131.4725 120.1825 132.2325 120.5975 ;
      RECT  132.6475 120.1825 133.4075 120.5975 ;
      RECT  133.8225 120.1825 134.5825 120.5975 ;
      RECT  134.9975 120.1825 135.7575 120.5975 ;
      RECT  136.1725 120.1825 136.9325 120.5975 ;
      RECT  137.3475 120.1825 138.1075 120.5975 ;
      RECT  138.5225 120.1825 139.2825 120.5975 ;
      RECT  139.6975 120.1825 140.4575 120.5975 ;
      RECT  140.8725 120.1825 141.6325 120.5975 ;
      RECT  142.0475 120.1825 142.8075 120.5975 ;
      RECT  143.2225 120.1825 143.9825 120.5975 ;
      RECT  144.3975 120.1825 145.1575 120.5975 ;
      RECT  145.5725 120.1825 146.3325 120.5975 ;
      RECT  146.7475 120.1825 147.5075 120.5975 ;
      RECT  147.9225 120.1825 148.6825 120.5975 ;
      RECT  149.0975 120.1825 149.8575 120.5975 ;
      RECT  150.2725 120.1825 151.0325 120.5975 ;
      RECT  151.4475 120.1825 152.2075 120.5975 ;
      RECT  152.6225 120.1825 153.3825 120.5975 ;
      RECT  153.7975 120.1825 154.5575 120.5975 ;
      RECT  154.9725 120.1825 155.7325 120.5975 ;
      RECT  156.1475 120.1825 156.9075 120.5975 ;
      RECT  157.3225 120.1825 158.0825 120.5975 ;
      RECT  158.4975 120.1825 159.2575 120.5975 ;
      RECT  159.6725 120.1825 160.4325 120.5975 ;
      RECT  160.8475 120.1825 161.6075 120.5975 ;
      RECT  162.0225 120.1825 162.7825 120.5975 ;
      RECT  163.1975 120.1825 163.9575 120.5975 ;
      RECT  164.3725 120.1825 165.1325 120.5975 ;
      RECT  165.5475 120.1825 166.3075 120.5975 ;
      RECT  166.7225 120.1825 167.4825 120.5975 ;
      RECT  167.8975 120.1825 168.6575 120.5975 ;
      RECT  169.0725 120.1825 169.8325 120.5975 ;
      RECT  170.2475 120.1825 171.0075 120.5975 ;
      RECT  171.4225 120.1825 172.1825 120.5975 ;
      RECT  172.5975 120.1825 173.3575 120.5975 ;
      RECT  173.7725 120.1825 174.5325 120.5975 ;
      RECT  174.9475 120.1825 175.7075 120.5975 ;
      RECT  176.1225 120.1825 176.8825 120.5975 ;
      RECT  177.2975 120.1825 178.0575 120.5975 ;
      RECT  178.4725 120.1825 179.2325 120.5975 ;
      RECT  179.6475 120.1825 180.4075 120.5975 ;
      RECT  180.8225 120.1825 181.5825 120.5975 ;
      RECT  181.9975 120.1825 182.7575 120.5975 ;
      RECT  183.1725 120.1825 183.9325 120.5975 ;
      RECT  184.3475 120.1825 185.1075 120.5975 ;
      RECT  185.5225 120.1825 186.2825 120.5975 ;
      RECT  186.6975 120.1825 187.4575 120.5975 ;
      RECT  187.8725 120.1825 188.6325 120.5975 ;
      RECT  189.0475 120.1825 189.8075 120.5975 ;
      RECT  190.2225 120.1825 190.9825 120.5975 ;
      RECT  191.3975 120.1825 192.1575 120.5975 ;
      RECT  192.5725 120.1825 193.3325 120.5975 ;
      RECT  193.7475 120.1825 194.5075 120.5975 ;
      RECT  194.9225 120.1825 195.6825 120.5975 ;
      RECT  196.0975 120.1825 196.8575 120.5975 ;
      RECT  197.2725 120.1825 198.0325 120.5975 ;
      RECT  198.4475 120.1825 199.2075 120.5975 ;
      RECT  199.6225 120.1825 200.3825 120.5975 ;
      RECT  200.7975 120.1825 201.5575 120.5975 ;
      RECT  201.9725 120.1825 202.7325 120.5975 ;
      RECT  203.1475 120.1825 203.9075 120.5975 ;
      RECT  204.3225 120.1825 205.0825 120.5975 ;
      RECT  205.4975 120.1825 206.2575 120.5975 ;
      RECT  206.6725 120.1825 207.4325 120.5975 ;
      RECT  207.8475 120.1825 208.6075 120.5975 ;
      RECT  209.0225 120.1825 209.7825 120.5975 ;
      RECT  210.1975 120.1825 210.9575 120.5975 ;
      RECT  211.3725 120.1825 212.1325 120.5975 ;
      RECT  212.5475 120.1825 213.3075 120.5975 ;
      RECT  213.7225 120.1825 214.4825 120.5975 ;
      RECT  214.8975 120.1825 215.6575 120.5975 ;
      RECT  216.0725 120.1825 216.8325 120.5975 ;
      RECT  217.2475 120.1825 218.0075 120.5975 ;
      RECT  218.4225 120.1825 219.1825 120.5975 ;
      RECT  219.5975 120.1825 220.3575 120.5975 ;
      RECT  220.7725 120.1825 221.5325 120.5975 ;
      RECT  221.9475 120.1825 222.7075 120.5975 ;
      RECT  223.1225 120.1825 223.8825 120.5975 ;
      RECT  224.2975 120.1825 225.0575 120.5975 ;
      RECT  225.4725 120.1825 226.2325 120.5975 ;
      RECT  226.6475 120.1825 227.4075 120.5975 ;
      RECT  227.8225 120.1825 228.5825 120.5975 ;
      RECT  228.9975 120.1825 229.7575 120.5975 ;
      RECT  230.1725 120.1825 230.9325 120.5975 ;
      RECT  231.3475 120.1825 232.1075 120.5975 ;
      RECT  232.5225 120.1825 233.2825 120.5975 ;
      RECT  233.6975 120.1825 234.4575 120.5975 ;
      RECT  234.8725 120.1825 235.6325 120.5975 ;
      RECT  236.0475 120.1825 236.8075 120.5975 ;
      RECT  237.2225 120.1825 237.9825 120.5975 ;
      RECT  238.3975 120.1825 239.1575 120.5975 ;
      RECT  239.5725 120.1825 240.3325 120.5975 ;
      RECT  240.7475 120.1825 241.5075 120.5975 ;
      RECT  241.9225 120.1825 242.6825 120.5975 ;
      RECT  243.0975 120.1825 243.8575 120.5975 ;
      RECT  244.2725 120.1825 245.0325 120.5975 ;
      RECT  245.4475 120.1825 246.2075 120.5975 ;
      RECT  246.6225 120.1825 247.3825 120.5975 ;
      RECT  247.7975 120.1825 248.5575 120.5975 ;
      RECT  248.9725 120.1825 249.7325 120.5975 ;
      RECT  250.1475 120.1825 250.9075 120.5975 ;
      RECT  251.3225 120.1825 252.0825 120.5975 ;
      RECT  252.4975 120.1825 253.2575 120.5975 ;
      RECT  253.6725 120.1825 254.4325 120.5975 ;
      RECT  254.8475 120.1825 255.6075 120.5975 ;
      RECT  256.0225 120.1825 256.7825 120.5975 ;
      RECT  257.1975 120.1825 257.9575 120.5975 ;
      RECT  258.3725 120.1825 259.1325 120.5975 ;
      RECT  259.5475 120.1825 260.3075 120.5975 ;
      RECT  260.7225 120.1825 261.4825 120.5975 ;
      RECT  261.8975 120.1825 262.6575 120.5975 ;
      RECT  263.0725 120.1825 263.8325 120.5975 ;
      RECT  264.2475 120.1825 265.0075 120.5975 ;
      RECT  265.4225 120.1825 266.1825 120.5975 ;
      RECT  266.5975 120.1825 267.3575 120.5975 ;
      RECT  267.7725 120.1825 268.5325 120.5975 ;
      RECT  268.9475 120.1825 269.7075 120.5975 ;
      RECT  270.1225 120.1825 270.8825 120.5975 ;
      RECT  271.2975 120.1825 272.0575 120.5975 ;
      RECT  272.4725 120.1825 273.2325 120.5975 ;
      RECT  273.6475 120.1825 274.4075 120.5975 ;
      RECT  274.8225 120.1825 275.5825 120.5975 ;
      RECT  275.9975 120.1825 276.7575 120.5975 ;
      RECT  277.1725 120.1825 277.9325 120.5975 ;
      RECT  278.3475 120.1825 279.1075 120.5975 ;
      RECT  279.5225 120.1825 280.2825 120.5975 ;
      RECT  280.6975 120.1825 281.4575 120.5975 ;
      RECT  281.8725 120.1825 282.6325 120.5975 ;
      RECT  283.0475 120.1825 283.8075 120.5975 ;
      RECT  284.2225 120.1825 284.9825 120.5975 ;
      RECT  285.3975 120.1825 286.1575 120.5975 ;
      RECT  286.5725 120.1825 287.3325 120.5975 ;
      RECT  287.7475 120.1825 288.5075 120.5975 ;
      RECT  288.9225 120.1825 289.6825 120.5975 ;
      RECT  290.0975 120.1825 290.8575 120.5975 ;
      RECT  291.2725 120.1825 292.0325 120.5975 ;
      RECT  292.4475 120.1825 293.2075 120.5975 ;
      RECT  293.6225 120.1825 294.3825 120.5975 ;
      RECT  294.7975 120.1825 295.5575 120.5975 ;
      RECT  295.9725 120.1825 296.7325 120.5975 ;
      RECT  297.1475 120.1825 297.9075 120.5975 ;
      RECT  298.3225 120.1825 299.0825 120.5975 ;
      RECT  299.4975 120.1825 300.2575 120.5975 ;
      RECT  300.6725 120.1825 301.4325 120.5975 ;
      RECT  301.8475 120.1825 302.6075 120.5975 ;
      RECT  303.0225 120.1825 303.7825 120.5975 ;
      RECT  304.1975 120.1825 304.9575 120.5975 ;
      RECT  305.3725 120.1825 306.1325 120.5975 ;
      RECT  306.5475 120.1825 307.3075 120.5975 ;
      RECT  307.7225 120.1825 308.4825 120.5975 ;
      RECT  308.8975 120.1825 309.6575 120.5975 ;
      RECT  310.0725 120.1825 310.8325 120.5975 ;
      RECT  311.2475 120.1825 312.0075 120.5975 ;
      RECT  312.4225 120.1825 313.1825 120.5975 ;
      RECT  313.5975 120.1825 314.3575 120.5975 ;
      RECT  314.7725 120.1825 315.5325 120.5975 ;
      RECT  315.9475 120.1825 316.7075 120.5975 ;
      RECT  317.1225 120.1825 317.8825 120.5975 ;
      RECT  318.2975 120.1825 319.0575 120.5975 ;
      RECT  319.4725 120.1825 320.2325 120.5975 ;
      RECT  320.6475 120.1825 321.4075 120.5975 ;
      RECT  321.8225 120.1825 322.5825 120.5975 ;
      RECT  322.9975 120.1825 323.7575 120.5975 ;
      RECT  324.1725 120.1825 324.9325 120.5975 ;
      RECT  325.3475 120.1825 326.1075 120.5975 ;
      RECT  326.5225 120.1825 327.2825 120.5975 ;
      RECT  327.6975 120.1825 328.4575 120.5975 ;
      RECT  328.8725 120.1825 329.6325 120.5975 ;
      RECT  330.0475 120.1825 330.8075 120.5975 ;
      RECT  331.2225 120.1825 331.9825 120.5975 ;
      RECT  332.3975 120.1825 333.1575 120.5975 ;
      RECT  333.5725 120.1825 334.3325 120.5975 ;
      RECT  334.7475 120.1825 335.5075 120.5975 ;
      RECT  335.9225 120.1825 336.6825 120.5975 ;
      RECT  337.0975 120.1825 337.8575 120.5975 ;
      RECT  338.2725 120.1825 339.0325 120.5975 ;
      RECT  339.4475 120.1825 340.2075 120.5975 ;
      RECT  340.6225 120.1825 341.3825 120.5975 ;
      RECT  341.7975 120.1825 342.5575 120.5975 ;
      RECT  342.9725 120.1825 343.7325 120.5975 ;
      RECT  344.1475 120.1825 344.9075 120.5975 ;
      RECT  345.3225 120.1825 346.0825 120.5975 ;
      RECT  346.4975 120.1825 347.2575 120.5975 ;
      RECT  347.6725 120.1825 348.4325 120.5975 ;
      RECT  348.8475 120.1825 349.6075 120.5975 ;
      RECT  350.0225 120.1825 350.7825 120.5975 ;
      RECT  351.1975 120.1825 351.9575 120.5975 ;
      RECT  352.3725 120.1825 353.1325 120.5975 ;
      RECT  353.5475 120.1825 354.3075 120.5975 ;
      RECT  354.7225 120.1825 355.4825 120.5975 ;
      RECT  355.8975 120.1825 356.6575 120.5975 ;
      RECT  357.0725 120.1825 357.8325 120.5975 ;
      RECT  358.2475 120.1825 359.0075 120.5975 ;
      RECT  359.4225 120.1825 360.1825 120.5975 ;
      RECT  360.5975 120.1825 361.3575 120.5975 ;
      RECT  361.7725 120.1825 362.5325 120.5975 ;
      RECT  362.9475 120.1825 363.7075 120.5975 ;
      RECT  364.1225 120.1825 364.8825 120.5975 ;
      RECT  365.2975 120.1825 366.0575 120.5975 ;
      RECT  366.4725 120.1825 367.2325 120.5975 ;
      RECT  367.6475 120.1825 368.4075 120.5975 ;
      RECT  368.8225 120.1825 369.5825 120.5975 ;
      RECT  369.9975 120.1825 398.91 120.5975 ;
      RECT  399.325 1.38 661.0475 2.33 ;
      RECT  399.325 2.745 661.0475 49.07 ;
      RECT  661.0475 1.38 661.4625 2.33 ;
      RECT  661.0475 2.745 661.4625 49.07 ;
      RECT  661.4625 1.38 752.635 2.33 ;
      RECT  661.4625 2.745 752.635 49.07 ;
      RECT  66.45 69.61 66.5475 70.025 ;
      RECT  66.45 70.025 66.5475 128.1325 ;
      RECT  66.9625 69.61 88.7575 70.025 ;
      RECT  89.1725 49.485 392.8975 63.63 ;
      RECT  89.1725 63.63 392.8975 64.045 ;
      RECT  393.3125 63.63 398.91 64.045 ;
      RECT  66.865 1.38 146.2475 2.33 ;
      RECT  146.2475 1.38 146.6625 2.33 ;
      RECT  146.6625 1.38 398.91 2.33 ;
      RECT  392.8975 61.055 393.3125 63.63 ;
      RECT  453.9475 49.485 457.495 125.525 ;
      RECT  453.9475 125.525 457.495 125.94 ;
      RECT  453.9475 125.94 457.495 126.805 ;
      RECT  457.495 49.485 457.91 125.525 ;
      RECT  457.495 125.94 457.91 126.805 ;
      RECT  457.91 49.485 459.635 125.525 ;
      RECT  457.91 125.525 459.635 125.94 ;
      RECT  457.91 125.94 459.635 126.805 ;
      RECT  66.865 49.07 72.72 49.4675 ;
      RECT  66.865 49.4675 72.72 49.485 ;
      RECT  72.72 49.07 73.135 49.4675 ;
      RECT  73.135 49.4675 398.91 49.485 ;
      RECT  66.9625 49.485 72.72 49.8825 ;
      RECT  66.9625 49.8825 72.72 69.61 ;
      RECT  72.72 49.8825 73.135 69.61 ;
      RECT  73.135 49.485 88.7575 49.8825 ;
      RECT  73.135 49.8825 88.7575 69.61 ;
      RECT  66.5475 55.075 66.865 60.64 ;
      RECT  66.865 55.075 66.9625 60.64 ;
      RECT  61.145 1.38 66.1675 2.33 ;
      RECT  61.145 2.33 66.1675 2.745 ;
      RECT  66.1675 1.38 66.45 2.33 ;
      RECT  66.1675 2.745 66.45 75.2 ;
      RECT  66.45 1.38 66.5475 2.33 ;
      RECT  66.45 2.745 66.5475 69.61 ;
      RECT  66.5475 1.38 66.5825 2.33 ;
      RECT  66.5825 1.38 66.865 2.33 ;
      RECT  66.5825 2.33 66.865 2.745 ;
      RECT  501.3025 2.33 512.3275 2.745 ;
      RECT  512.7425 2.33 523.7675 2.745 ;
      RECT  66.865 2.745 85.5725 46.3075 ;
      RECT  66.865 46.3075 85.5725 46.6575 ;
      RECT  85.5725 46.6575 146.2475 49.07 ;
      RECT  146.2475 46.6575 146.6625 49.07 ;
      RECT  146.6625 46.6575 371.1375 49.07 ;
      RECT  371.1375 2.745 398.91 46.3075 ;
      RECT  371.1375 46.3075 398.91 46.6575 ;
      RECT  371.1375 46.6575 398.91 49.07 ;
      RECT  638.5825 2.33 649.6075 2.745 ;
      RECT  650.0225 2.33 661.0475 2.745 ;
      RECT  489.8625 2.33 500.8875 2.745 ;
      RECT  392.8975 73.015 393.3125 120.1825 ;
      RECT  88.7575 117.975 89.1725 120.1825 ;
      RECT  66.9625 70.025 85.5725 117.625 ;
      RECT  66.9625 117.625 85.5725 117.975 ;
      RECT  66.9625 117.975 85.5725 120.1825 ;
      RECT  85.5725 117.975 88.7575 120.1825 ;
      RECT  89.1725 117.975 370.6675 120.1825 ;
      RECT  370.6675 117.625 392.8975 117.975 ;
      RECT  370.6675 117.975 392.8975 120.1825 ;
      RECT  66.865 49.485 66.9625 51.67 ;
      RECT  66.865 52.085 66.9625 54.66 ;
      RECT  66.5475 2.745 66.5825 51.67 ;
      RECT  66.5475 52.085 66.5825 54.66 ;
      RECT  66.5825 2.745 66.865 51.67 ;
      RECT  66.5825 52.085 66.865 54.66 ;
      RECT  741.5425 2.33 752.635 2.745 ;
      RECT  85.5725 2.745 146.2475 40.8725 ;
      RECT  146.2475 2.745 146.6625 40.8725 ;
      RECT  146.6625 2.745 370.6675 40.8725 ;
      RECT  370.6675 2.745 371.1375 40.8725 ;
      RECT  370.6675 40.8725 371.1375 41.2225 ;
      RECT  370.6675 41.2225 371.1375 46.3075 ;
      RECT  627.1425 2.33 638.1675 2.745 ;
      RECT  146.6625 2.33 157.6875 2.745 ;
      RECT  158.1025 2.33 169.1275 2.745 ;
      RECT  392.8975 64.045 393.3125 69.61 ;
      RECT  392.8975 70.025 393.3125 72.6 ;
      RECT  524.1825 2.33 535.2075 2.745 ;
      RECT  386.9025 2.33 397.9275 2.745 ;
      RECT  398.3425 2.33 398.91 2.745 ;
      RECT  135.2225 2.33 146.2475 2.745 ;
      RECT  592.8225 2.33 603.8475 2.745 ;
      RECT  370.6675 64.045 386.725 110.6825 ;
      RECT  370.6675 110.6825 386.725 111.0975 ;
      RECT  386.725 64.045 387.14 110.6825 ;
      RECT  386.725 111.0975 387.14 117.625 ;
      RECT  387.14 64.045 392.8975 110.6825 ;
      RECT  387.14 110.6825 392.8975 111.0975 ;
      RECT  387.14 111.0975 392.8975 117.625 ;
      RECT  455.5425 2.33 466.5675 2.745 ;
      RECT  466.9825 2.33 478.0075 2.745 ;
      RECT  478.4225 2.33 489.4475 2.745 ;
      RECT  238.1825 2.33 249.2075 2.745 ;
      RECT  329.7025 2.33 340.7275 2.745 ;
      RECT  341.1425 2.33 352.1675 2.745 ;
      RECT  375.4625 2.33 386.4875 2.745 ;
      RECT  249.6225 2.33 260.6475 2.745 ;
      RECT  261.0625 2.33 272.0875 2.745 ;
      RECT  318.2625 2.33 329.2875 2.745 ;
      RECT  226.7425 2.33 237.7675 2.745 ;
      RECT  88.7575 49.485 89.1725 113.7275 ;
      RECT  85.5725 70.025 88.7575 113.7275 ;
      RECT  89.1725 64.045 370.6675 113.7275 ;
      RECT  370.6675 111.0975 372.3125 113.7275 ;
      RECT  372.3125 113.7275 386.725 114.0775 ;
      RECT  372.3125 114.0775 386.725 117.625 ;
      RECT  272.5025 2.33 283.5275 2.745 ;
      RECT  283.9425 2.33 294.9675 2.745 ;
      RECT  569.9425 2.33 580.9675 2.745 ;
      RECT  581.3825 2.33 592.4075 2.745 ;
      RECT  730.1025 2.33 741.1275 2.745 ;
      RECT  558.5025 2.33 569.5275 2.745 ;
      RECT  604.2625 2.33 615.2875 2.745 ;
      RECT  615.7025 2.33 626.7275 2.745 ;
      RECT  718.6625 2.33 729.6875 2.745 ;
      RECT  0.56 31.11 2.285 31.975 ;
      RECT  0.56 31.975 2.285 32.39 ;
      RECT  0.56 32.39 2.285 75.2 ;
      RECT  2.285 31.11 2.7 31.975 ;
      RECT  2.285 32.39 2.7 75.2 ;
      RECT  2.7 31.11 6.1075 31.975 ;
      RECT  2.7 31.975 6.1075 32.39 ;
      RECT  2.7 32.39 6.1075 75.2 ;
      RECT  66.5475 70.025 66.865 72.6 ;
      RECT  66.5475 73.015 66.865 128.1325 ;
      RECT  66.865 70.025 66.9625 72.6 ;
      RECT  66.865 73.015 66.9625 120.1825 ;
      RECT  203.8625 2.33 214.8875 2.745 ;
      RECT  215.3025 2.33 226.3275 2.745 ;
      RECT  66.865 2.33 77.6075 2.745 ;
      RECT  78.0225 2.33 89.0475 2.745 ;
      RECT  661.4625 2.33 672.4875 2.745 ;
      RECT  672.9025 2.33 683.9275 2.745 ;
      RECT  295.3825 2.33 306.4075 2.745 ;
      RECT  306.8225 2.33 317.8475 2.745 ;
      RECT  392.8975 55.075 393.3125 60.64 ;
      RECT  89.4625 2.33 100.4875 2.745 ;
      RECT  100.9025 2.33 111.9275 2.745 ;
      RECT  112.3425 2.33 123.3675 2.745 ;
      RECT  123.7825 2.33 134.8075 2.745 ;
      RECT  684.3425 2.33 695.3675 2.745 ;
      RECT  192.4225 2.33 203.4475 2.745 ;
      RECT  421.2225 2.33 432.2475 2.745 ;
      RECT  73.135 49.07 84.4275 49.095 ;
      RECT  73.135 49.095 84.4275 49.4675 ;
      RECT  84.4275 49.095 84.8425 49.4675 ;
      RECT  84.8425 49.07 398.91 49.095 ;
      RECT  84.8425 49.095 398.91 49.4675 ;
      RECT  66.865 46.6575 84.4275 48.68 ;
      RECT  66.865 48.68 84.4275 49.07 ;
      RECT  84.4275 46.6575 84.8425 48.68 ;
      RECT  84.8425 46.6575 85.5725 48.68 ;
      RECT  84.8425 48.68 85.5725 49.07 ;
      RECT  399.325 2.33 409.3675 2.745 ;
      RECT  409.7825 2.33 420.8075 2.745 ;
      RECT  432.6625 2.33 443.6875 2.745 ;
      RECT  444.1025 2.33 455.1275 2.745 ;
      RECT  535.6225 2.33 546.6475 2.745 ;
      RECT  547.0625 2.33 558.0875 2.745 ;
      RECT  66.5475 61.055 66.865 63.63 ;
      RECT  66.5475 64.045 66.865 69.61 ;
      RECT  66.865 61.055 66.9625 63.63 ;
      RECT  66.865 64.045 66.9625 69.61 ;
      RECT  695.7825 2.33 706.8075 2.745 ;
      RECT  707.2225 2.33 718.2475 2.745 ;
      RECT  352.5825 2.33 363.6075 2.745 ;
      RECT  364.0225 2.33 375.0475 2.745 ;
      RECT  169.5425 2.33 180.5675 2.745 ;
      RECT  180.9825 2.33 192.0075 2.745 ;
      RECT  392.8975 49.485 393.3125 51.67 ;
      RECT  392.8975 52.085 393.3125 54.66 ;
      RECT  372.3125 111.0975 375.0175 111.47 ;
      RECT  372.3125 111.47 375.0175 111.885 ;
      RECT  372.3125 111.885 375.0175 113.7275 ;
      RECT  375.0175 111.0975 375.4325 111.47 ;
      RECT  375.0175 111.885 375.4325 113.7275 ;
      RECT  375.4325 111.0975 386.725 111.47 ;
      RECT  375.4325 111.47 386.725 111.885 ;
      RECT  375.4325 111.885 386.725 113.7275 ;
      RECT  66.865 0.275 320.7075 0.965 ;
      RECT  320.7075 0.275 321.1225 0.965 ;
      RECT  321.1225 0.275 752.635 0.965 ;
      RECT  309.6825 0.14 320.7075 0.275 ;
      RECT  61.145 2.745 65.02 53.165 ;
      RECT  61.145 53.165 65.02 53.58 ;
      RECT  61.145 53.58 65.02 75.2 ;
      RECT  65.435 2.745 66.1675 53.165 ;
      RECT  65.435 53.165 66.1675 53.58 ;
      RECT  65.435 53.58 66.1675 75.2 ;
      RECT  85.5725 41.2225 146.2475 42.9225 ;
      RECT  85.5725 43.2725 146.2475 46.3075 ;
      RECT  146.2475 41.2225 146.6625 42.9225 ;
      RECT  146.2475 43.2725 146.6625 46.3075 ;
      RECT  146.6625 41.2225 370.6675 42.9225 ;
      RECT  146.6625 43.2725 370.6675 46.3075 ;
      RECT  393.3125 64.045 394.425 74.095 ;
      RECT  393.3125 74.095 394.425 74.51 ;
      RECT  393.3125 74.51 394.425 120.1825 ;
      RECT  394.425 74.51 394.84 120.1825 ;
      RECT  394.84 64.045 398.91 74.095 ;
      RECT  394.84 74.095 398.91 74.51 ;
      RECT  394.84 74.51 398.91 120.1825 ;
      RECT  393.3125 49.485 394.425 56.155 ;
      RECT  393.3125 56.155 394.425 56.57 ;
      RECT  393.3125 56.57 394.425 63.63 ;
      RECT  394.84 49.485 398.91 56.155 ;
      RECT  394.84 56.155 398.91 56.57 ;
      RECT  394.84 56.57 398.91 63.63 ;
      RECT  65.02 74.51 65.435 75.2 ;
      RECT  721.5225 0.14 732.5475 0.275 ;
      RECT  446.9625 0.14 457.9875 0.275 ;
      RECT  394.425 56.57 394.84 59.145 ;
      RECT  65.02 53.58 65.435 56.155 ;
      RECT  412.6425 0.14 423.6675 0.275 ;
      RECT  394.425 49.485 394.84 50.175 ;
      RECT  710.0825 0.14 721.1075 0.275 ;
      RECT  218.1625 0.14 229.1875 0.275 ;
      RECT  394.425 50.59 394.84 53.165 ;
      RECT  394.425 53.58 394.84 56.155 ;
      RECT  80.8825 0.14 91.9075 0.275 ;
      RECT  0.56 1.38 2.285 29.505 ;
      RECT  0.56 29.505 2.285 29.92 ;
      RECT  0.56 29.92 2.285 30.61 ;
      RECT  2.285 1.38 2.7 29.505 ;
      RECT  2.285 29.92 2.7 30.61 ;
      RECT  2.7 1.38 60.73 29.505 ;
      RECT  2.7 29.505 60.73 29.92 ;
      RECT  2.7 29.92 60.73 30.61 ;
      RECT  399.325 127.305 457.495 127.995 ;
      RECT  399.325 127.995 457.495 128.1325 ;
      RECT  457.495 127.305 457.91 127.995 ;
      RECT  457.91 127.305 459.635 127.995 ;
      RECT  457.91 127.995 459.635 128.1325 ;
      RECT  664.3225 0.14 675.3475 0.275 ;
      RECT  65.02 2.745 65.435 50.175 ;
      RECT  65.02 50.59 65.435 53.165 ;
      RECT  321.1225 0.14 332.1475 0.275 ;
      RECT  172.4025 0.14 183.4275 0.275 ;
      RECT  206.7225 0.14 217.7475 0.275 ;
      RECT  595.6825 0.14 606.7075 0.275 ;
      RECT  394.425 64.045 394.84 65.125 ;
      RECT  66.865 0.14 69.0275 0.275 ;
      RECT  69.4425 0.14 80.4675 0.275 ;
      RECT  126.6425 0.14 137.6675 0.275 ;
      RECT  138.0825 0.14 149.1075 0.275 ;
      RECT  492.7225 0.14 503.7475 0.275 ;
      RECT  504.1625 0.14 515.1875 0.275 ;
      RECT  652.8825 0.14 663.9075 0.275 ;
      RECT  394.425 65.54 394.84 68.115 ;
      RECT  698.6425 0.14 709.6675 0.275 ;
      RECT  458.4025 0.14 469.4275 0.275 ;
      RECT  572.8025 0.14 583.8275 0.275 ;
      RECT  584.2425 0.14 595.2675 0.275 ;
      RECT  561.3625 0.14 572.3875 0.275 ;
      RECT  424.0825 0.14 435.1075 0.275 ;
      RECT  435.5225 0.14 446.5475 0.275 ;
      RECT  732.9625 0.14 743.9875 0.275 ;
      RECT  744.4025 0.14 752.635 0.275 ;
      RECT  183.8425 0.14 194.8675 0.275 ;
      RECT  195.2825 0.14 206.3075 0.275 ;
      RECT  115.2025 0.14 126.2275 0.275 ;
      RECT  149.5225 0.14 160.5475 0.275 ;
      RECT  160.9625 0.14 171.9875 0.275 ;
      RECT  675.7625 0.14 686.7875 0.275 ;
      RECT  687.2025 0.14 698.2275 0.275 ;
      RECT  88.7575 114.0775 89.1725 115.7325 ;
      RECT  88.7575 116.0825 89.1725 117.625 ;
      RECT  85.5725 114.0775 88.7575 115.7325 ;
      RECT  85.5725 116.0825 88.7575 117.625 ;
      RECT  89.1725 114.0775 370.6675 115.7325 ;
      RECT  89.1725 116.0825 370.6675 117.625 ;
      RECT  370.6675 114.0775 370.7025 115.7325 ;
      RECT  370.6675 116.0825 370.7025 117.625 ;
      RECT  370.7025 114.0775 372.3125 115.7325 ;
      RECT  370.7025 115.7325 372.3125 116.0825 ;
      RECT  370.7025 116.0825 372.3125 117.625 ;
      RECT  65.02 62.55 65.435 65.125 ;
      RECT  229.6025 0.14 240.6275 0.275 ;
      RECT  241.0425 0.14 252.0675 0.275 ;
      RECT  630.0025 0.14 641.0275 0.275 ;
      RECT  641.4425 0.14 652.4675 0.275 ;
      RECT  275.3625 0.14 286.3875 0.275 ;
      RECT  65.02 56.57 65.435 59.145 ;
      RECT  65.02 59.56 65.435 62.135 ;
      RECT  92.3225 0.14 103.3475 0.275 ;
      RECT  103.7625 0.14 114.7875 0.275 ;
      RECT  394.425 59.56 394.84 62.135 ;
      RECT  394.425 62.55 394.84 63.63 ;
      RECT  469.8425 0.14 480.8675 0.275 ;
      RECT  481.2825 0.14 492.3075 0.275 ;
      RECT  65.02 65.54 65.435 68.115 ;
      RECT  515.6025 0.14 526.6275 0.275 ;
      RECT  527.0425 0.14 538.0675 0.275 ;
      RECT  389.7625 0.14 400.7875 0.275 ;
      RECT  401.2025 0.14 412.2275 0.275 ;
      RECT  355.4425 0.14 366.4675 0.275 ;
      RECT  607.1225 0.14 618.1475 0.275 ;
      RECT  618.5625 0.14 629.5875 0.275 ;
      RECT  332.5625 0.14 343.5875 0.275 ;
      RECT  344.0025 0.14 355.0275 0.275 ;
      RECT  252.4825 0.14 263.5075 0.275 ;
      RECT  263.9225 0.14 274.9475 0.275 ;
      RECT  366.8825 0.14 377.9075 0.275 ;
      RECT  378.3225 0.14 389.3475 0.275 ;
      RECT  286.8025 0.14 297.8275 0.275 ;
      RECT  298.2425 0.14 309.2675 0.275 ;
      RECT  538.4825 0.14 549.5075 0.275 ;
      RECT  549.9225 0.14 560.9475 0.275 ;
      RECT  65.02 68.53 65.435 71.105 ;
      RECT  65.02 71.52 65.435 74.095 ;
      RECT  394.425 68.53 394.84 71.105 ;
      RECT  394.425 71.52 394.84 74.095 ;
   LAYER  metal4 ;
      RECT  0.14 113.4525 373.795 128.1325 ;
      RECT  373.795 0.14 374.495 46.8625 ;
      RECT  373.795 113.4525 374.495 128.1325 ;
      RECT  459.0875 46.8625 459.7875 95.7425 ;
      RECT  459.7875 46.8625 752.635 95.7425 ;
      RECT  459.7875 95.7425 752.635 113.4525 ;
      RECT  459.0875 118.705 459.7875 128.1325 ;
      RECT  459.7875 113.4525 752.635 118.705 ;
      RECT  459.7875 118.705 752.635 128.1325 ;
      RECT  374.495 110.6025 387.2 113.4525 ;
      RECT  387.2 110.6025 387.9 113.4525 ;
      RECT  374.495 113.4525 396.33 115.5025 ;
      RECT  374.495 115.5025 396.33 118.705 ;
      RECT  396.33 113.4525 397.03 115.5025 ;
      RECT  374.495 118.705 396.33 126.0825 ;
      RECT  374.495 126.0825 396.33 128.1325 ;
      RECT  396.33 126.0825 397.03 128.1325 ;
      RECT  0.14 73.9525 60.305 89.4725 ;
      RECT  0.14 89.4725 60.305 113.4525 ;
      RECT  60.305 46.8625 61.005 73.9525 ;
      RECT  60.305 89.4725 61.005 113.4525 ;
      RECT  61.005 110.6025 71.96 113.4525 ;
      RECT  71.96 110.6025 72.66 113.4525 ;
      RECT  374.495 50.0325 374.875 95.7425 ;
      RECT  374.495 95.7425 374.875 110.5325 ;
      RECT  374.495 110.5325 374.875 110.6025 ;
      RECT  374.875 110.5325 375.575 110.6025 ;
      RECT  63.025 0.14 63.725 31.8325 ;
      RECT  63.725 0.14 373.795 31.8325 ;
      RECT  63.725 31.8325 373.795 46.8625 ;
      RECT  61.005 46.8625 63.025 47.3525 ;
      RECT  61.005 47.3525 63.025 50.0325 ;
      RECT  63.025 47.3525 63.725 50.0325 ;
      RECT  63.725 46.8625 71.96 47.3525 ;
      RECT  84.285 110.5325 84.985 110.6025 ;
      RECT  72.66 110.6025 85.365 113.4525 ;
      RECT  84.985 50.0325 85.365 73.9525 ;
      RECT  84.985 73.9525 85.365 89.4725 ;
      RECT  84.985 89.4725 85.365 110.5325 ;
      RECT  84.985 110.5325 85.365 110.6025 ;
      RECT  399.05 0.14 399.75 35.2125 ;
      RECT  399.75 0.14 752.635 35.2125 ;
      RECT  399.75 35.2125 752.635 46.8625 ;
      RECT  399.75 46.8625 459.0875 50.0325 ;
      RECT  399.05 50.7325 399.75 95.7425 ;
      RECT  399.75 50.0325 459.0875 50.7325 ;
      RECT  0.14 46.8625 0.4075 62.1725 ;
      RECT  0.14 62.1725 0.4075 73.9525 ;
      RECT  0.4075 62.1725 1.1075 73.9525 ;
      RECT  0.14 31.8325 0.4075 39.21 ;
      RECT  0.14 39.21 0.4075 46.8625 ;
      RECT  0.4075 31.8325 1.1075 39.21 ;
      RECT  387.9 110.6025 453.53 113.0325 ;
      RECT  387.9 113.0325 453.53 113.4525 ;
      RECT  453.53 110.6025 454.23 113.0325 ;
      RECT  397.03 113.4525 453.53 115.5025 ;
      RECT  397.03 115.5025 453.53 118.705 ;
      RECT  397.03 118.705 453.53 126.0825 ;
      RECT  454.23 118.705 459.0875 126.0825 ;
      RECT  397.03 126.0825 453.53 128.1325 ;
      RECT  454.23 126.0825 459.0875 128.1325 ;
      RECT  61.005 50.0325 63.165 73.8875 ;
      RECT  61.005 73.8875 63.165 73.9525 ;
      RECT  63.165 50.0325 63.865 73.8875 ;
      RECT  61.005 73.9525 63.165 89.4725 ;
      RECT  61.005 89.4725 63.165 89.5375 ;
      RECT  61.005 89.5375 63.165 110.6025 ;
      RECT  63.165 89.5375 63.865 110.6025 ;
      RECT  0.14 0.14 5.825 29.3625 ;
      RECT  0.14 29.3625 5.825 31.8325 ;
      RECT  5.825 0.14 6.525 29.3625 ;
      RECT  6.525 0.14 63.025 29.3625 ;
      RECT  6.525 29.3625 63.025 31.8325 ;
      RECT  1.1075 31.8325 5.825 39.21 ;
      RECT  6.525 31.8325 63.025 39.21 ;
      RECT  5.825 44.8825 6.525 46.8625 ;
      RECT  6.525 39.21 63.025 44.8825 ;
      RECT  6.525 44.8825 63.025 46.8625 ;
      RECT  63.725 47.3525 70.025 50.0 ;
      RECT  63.725 50.0 70.025 50.0325 ;
      RECT  70.025 47.3525 70.725 50.0 ;
      RECT  70.725 47.3525 71.96 50.0 ;
      RECT  70.725 50.0 71.96 50.0325 ;
      RECT  63.865 50.0325 70.025 73.8875 ;
      RECT  70.725 50.0325 71.96 73.8875 ;
      RECT  63.865 73.8875 70.025 73.9525 ;
      RECT  70.725 73.8875 71.96 73.9525 ;
      RECT  63.865 73.9525 70.025 89.4725 ;
      RECT  70.725 73.9525 71.96 89.4725 ;
      RECT  63.865 89.4725 70.025 89.5375 ;
      RECT  70.725 89.4725 71.96 89.5375 ;
      RECT  63.865 89.5375 70.025 110.6025 ;
      RECT  70.725 89.5375 71.96 110.6025 ;
      RECT  387.9 95.7425 389.135 110.6025 ;
      RECT  387.9 46.8625 389.135 50.0 ;
      RECT  387.9 50.0 389.135 50.0325 ;
      RECT  389.135 46.8625 389.835 50.0 ;
      RECT  387.9 50.0325 389.135 50.7325 ;
      RECT  387.9 50.7325 389.135 95.7425 ;
      RECT  374.495 0.14 396.19 35.1475 ;
      RECT  374.495 35.1475 396.19 35.2125 ;
      RECT  396.19 0.14 396.89 35.1475 ;
      RECT  396.89 0.14 399.05 35.1475 ;
      RECT  396.89 35.1475 399.05 35.2125 ;
      RECT  374.495 35.2125 396.19 46.8625 ;
      RECT  396.89 35.2125 399.05 46.8625 ;
      RECT  389.835 46.8625 396.19 50.0 ;
      RECT  396.89 46.8625 399.05 50.0 ;
      RECT  389.835 50.0 396.19 50.0325 ;
      RECT  396.89 50.0 399.05 50.0325 ;
      RECT  389.835 50.0325 396.19 50.7325 ;
      RECT  396.89 50.0325 399.05 50.7325 ;
      RECT  389.835 50.7325 396.19 50.7975 ;
      RECT  389.835 50.7975 396.19 95.7425 ;
      RECT  396.19 50.7975 396.89 95.7425 ;
      RECT  396.89 50.7325 399.05 50.7975 ;
      RECT  396.89 50.7975 399.05 95.7425 ;
      RECT  399.75 50.7325 457.025 95.71 ;
      RECT  399.75 95.71 457.025 95.7425 ;
      RECT  457.025 50.7325 457.725 95.71 ;
      RECT  457.725 50.7325 459.0875 95.71 ;
      RECT  457.725 95.71 459.0875 95.7425 ;
      RECT  454.23 110.6025 457.025 113.0325 ;
      RECT  457.725 110.6025 459.0875 113.0325 ;
      RECT  454.23 113.0325 457.025 113.4525 ;
      RECT  457.725 113.0325 459.0875 113.4525 ;
      RECT  454.23 113.4525 457.025 115.5025 ;
      RECT  457.725 113.4525 459.0875 115.5025 ;
      RECT  454.23 115.5025 457.025 118.6725 ;
      RECT  454.23 118.6725 457.025 118.705 ;
      RECT  457.025 118.6725 457.725 118.705 ;
      RECT  457.725 115.5025 459.0875 118.6725 ;
      RECT  457.725 118.6725 459.0875 118.705 ;
      RECT  389.835 95.7425 457.025 110.6025 ;
      RECT  457.725 95.7425 459.0875 110.6025 ;
      RECT  374.495 46.8625 386.64 50.0 ;
      RECT  374.495 50.0 386.64 50.0325 ;
      RECT  386.64 46.8625 387.2 50.0 ;
      RECT  387.2 46.8625 387.34 50.0 ;
      RECT  387.34 46.8625 387.9 50.0 ;
      RECT  387.34 50.0 387.9 50.0325 ;
      RECT  375.575 50.0325 386.64 95.7425 ;
      RECT  375.575 95.7425 386.64 110.5325 ;
      RECT  375.575 110.5325 386.64 110.565 ;
      RECT  375.575 110.565 386.64 110.6025 ;
      RECT  386.64 110.565 387.2 110.6025 ;
      RECT  1.1075 46.8625 2.47 62.1725 ;
      RECT  3.17 46.8625 60.305 62.1725 ;
      RECT  1.1075 62.1725 2.47 62.205 ;
      RECT  1.1075 62.205 2.47 73.9525 ;
      RECT  2.47 62.205 3.17 73.9525 ;
      RECT  3.17 62.1725 60.305 62.205 ;
      RECT  3.17 62.205 60.305 73.9525 ;
      RECT  1.1075 39.21 2.47 39.2425 ;
      RECT  1.1075 39.2425 2.47 44.8825 ;
      RECT  2.47 39.21 3.17 39.2425 ;
      RECT  3.17 39.21 5.825 39.2425 ;
      RECT  3.17 39.2425 5.825 44.8825 ;
      RECT  1.1075 44.8825 2.47 46.8625 ;
      RECT  3.17 44.8825 5.825 46.8625 ;
      RECT  71.96 46.8625 72.52 50.0 ;
      RECT  71.96 50.0 72.52 50.0325 ;
      RECT  72.52 46.8625 72.66 50.0 ;
      RECT  73.22 50.0325 84.285 73.9525 ;
      RECT  73.22 73.9525 84.285 89.4725 ;
      RECT  73.22 89.4725 84.285 110.5325 ;
      RECT  72.66 110.565 73.22 110.6025 ;
      RECT  73.22 110.5325 84.285 110.565 ;
      RECT  73.22 110.565 84.285 110.6025 ;
      RECT  72.66 46.8625 73.22 50.0 ;
      RECT  73.22 46.8625 85.365 50.0 ;
      RECT  73.22 50.0 85.365 50.0325 ;
      RECT  86.525 46.8625 373.335 50.0325 ;
      RECT  86.525 110.6025 373.335 113.4525 ;
      RECT  86.525 50.0325 373.335 73.9525 ;
      RECT  86.525 73.9525 373.335 89.4725 ;
      RECT  86.525 89.4725 373.335 110.5325 ;
      RECT  86.525 110.5325 373.335 110.6025 ;
   END
END    freepdk45_sram_1w1r_40x240
END    LIBRARY
