VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1rw0r_64x80_20
   CLASS BLOCK ;
   SIZE 272.245 BY 126.1075 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.66 1.105 43.795 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.52 1.105 46.655 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.38 1.105 49.515 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.24 1.105 52.375 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.1 1.105 55.235 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.96 1.105 58.095 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.82 1.105 60.955 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.68 1.105 63.815 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.54 1.105 66.675 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.4 1.105 69.535 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.26 1.105 72.395 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.12 1.105 75.255 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.98 1.105 78.115 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.84 1.105 80.975 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.7 1.105 83.835 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.56 1.105 86.695 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.42 1.105 89.555 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.28 1.105 92.415 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.14 1.105 95.275 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.0 1.105 98.135 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.86 1.105 100.995 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.72 1.105 103.855 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.58 1.105 106.715 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.44 1.105 109.575 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.3 1.105 112.435 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.16 1.105 115.295 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.02 1.105 118.155 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.88 1.105 121.015 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.74 1.105 123.875 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.6 1.105 126.735 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.46 1.105 129.595 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.32 1.105 132.455 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.18 1.105 135.315 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.04 1.105 138.175 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.9 1.105 141.035 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.76 1.105 143.895 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.62 1.105 146.755 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.48 1.105 149.615 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.34 1.105 152.475 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.2 1.105 155.335 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.06 1.105 158.195 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.92 1.105 161.055 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.78 1.105 163.915 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.64 1.105 166.775 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.5 1.105 169.635 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.36 1.105 172.495 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.22 1.105 175.355 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.08 1.105 178.215 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.94 1.105 181.075 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.8 1.105 183.935 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.66 1.105 186.795 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.52 1.105 189.655 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.38 1.105 192.515 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.24 1.105 195.375 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.1 1.105 198.235 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.96 1.105 201.095 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.82 1.105 203.955 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.68 1.105 206.815 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.54 1.105 209.675 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.4 1.105 212.535 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.26 1.105 215.395 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.12 1.105 218.255 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.98 1.105 221.115 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.84 1.105 223.975 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.7 1.105 226.835 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.56 1.105 229.695 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.42 1.105 232.555 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.28 1.105 235.415 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.14 1.105 238.275 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.0 1.105 241.135 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.86 1.105 243.995 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.72 1.105 246.855 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.58 1.105 249.715 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.44 1.105 252.575 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.3 1.105 255.435 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.16 1.105 258.295 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.02 1.105 261.155 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.88 1.105 264.015 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.74 1.105 266.875 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.6 1.105 269.735 1.24 ;
      END
   END din0[79]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.5 60.0625 26.635 60.1975 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.5 62.7925 26.635 62.9275 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.5 65.0025 26.635 65.1375 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.5 67.7325 26.635 67.8675 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.5 69.9425 26.635 70.0775 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.5 72.6725 26.635 72.8075 ;
      END
   END addr0[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 15.3425 0.42 15.4775 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 18.0725 0.42 18.2075 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 15.4275 6.6625 15.5625 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.22 1.105 32.355 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.08 1.105 35.215 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.94 1.105 38.075 1.24 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.8 1.105 40.935 1.24 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.2625 26.9925 47.3975 27.1275 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.9675 26.9925 48.1025 27.1275 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.6725 26.9925 48.8075 27.1275 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.3775 26.9925 49.5125 27.1275 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.0825 26.9925 50.2175 27.1275 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.7875 26.9925 50.9225 27.1275 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.4925 26.9925 51.6275 27.1275 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.1975 26.9925 52.3325 27.1275 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.9025 26.9925 53.0375 27.1275 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.6075 26.9925 53.7425 27.1275 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.3125 26.9925 54.4475 27.1275 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.0175 26.9925 55.1525 27.1275 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.7225 26.9925 55.8575 27.1275 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.4275 26.9925 56.5625 27.1275 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.1325 26.9925 57.2675 27.1275 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.8375 26.9925 57.9725 27.1275 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.5425 26.9925 58.6775 27.1275 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.2475 26.9925 59.3825 27.1275 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.9525 26.9925 60.0875 27.1275 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.6575 26.9925 60.7925 27.1275 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.3625 26.9925 61.4975 27.1275 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.0675 26.9925 62.2025 27.1275 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.7725 26.9925 62.9075 27.1275 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.4775 26.9925 63.6125 27.1275 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.1825 26.9925 64.3175 27.1275 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.8875 26.9925 65.0225 27.1275 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.5925 26.9925 65.7275 27.1275 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.2975 26.9925 66.4325 27.1275 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.0025 26.9925 67.1375 27.1275 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.7075 26.9925 67.8425 27.1275 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.4125 26.9925 68.5475 27.1275 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.1175 26.9925 69.2525 27.1275 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.8225 26.9925 69.9575 27.1275 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.5275 26.9925 70.6625 27.1275 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.2325 26.9925 71.3675 27.1275 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.9375 26.9925 72.0725 27.1275 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.6425 26.9925 72.7775 27.1275 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.3475 26.9925 73.4825 27.1275 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.0525 26.9925 74.1875 27.1275 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.7575 26.9925 74.8925 27.1275 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.4625 26.9925 75.5975 27.1275 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.1675 26.9925 76.3025 27.1275 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.8725 26.9925 77.0075 27.1275 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.5775 26.9925 77.7125 27.1275 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.2825 26.9925 78.4175 27.1275 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.9875 26.9925 79.1225 27.1275 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.6925 26.9925 79.8275 27.1275 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.3975 26.9925 80.5325 27.1275 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.1025 26.9925 81.2375 27.1275 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.8075 26.9925 81.9425 27.1275 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.5125 26.9925 82.6475 27.1275 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.2175 26.9925 83.3525 27.1275 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.9225 26.9925 84.0575 27.1275 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.6275 26.9925 84.7625 27.1275 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.3325 26.9925 85.4675 27.1275 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.0375 26.9925 86.1725 27.1275 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.7425 26.9925 86.8775 27.1275 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.4475 26.9925 87.5825 27.1275 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.1525 26.9925 88.2875 27.1275 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.8575 26.9925 88.9925 27.1275 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.5625 26.9925 89.6975 27.1275 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.2675 26.9925 90.4025 27.1275 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.9725 26.9925 91.1075 27.1275 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.6775 26.9925 91.8125 27.1275 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.3825 26.9925 92.5175 27.1275 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.0875 26.9925 93.2225 27.1275 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.7925 26.9925 93.9275 27.1275 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.4975 26.9925 94.6325 27.1275 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.2025 26.9925 95.3375 27.1275 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.9075 26.9925 96.0425 27.1275 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.6125 26.9925 96.7475 27.1275 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.3175 26.9925 97.4525 27.1275 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.0225 26.9925 98.1575 27.1275 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.7275 26.9925 98.8625 27.1275 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.4325 26.9925 99.5675 27.1275 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.1375 26.9925 100.2725 27.1275 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.8425 26.9925 100.9775 27.1275 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.5475 26.9925 101.6825 27.1275 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.2525 26.9925 102.3875 27.1275 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.9575 26.9925 103.0925 27.1275 ;
      END
   END dout0[79]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  0.0 14.235 0.14 19.315 ;
         LAYER metal3 ;
         RECT  249.2975 2.47 249.4325 2.605 ;
         LAYER metal3 ;
         RECT  169.2175 2.47 169.3525 2.605 ;
         LAYER metal3 ;
         RECT  134.8975 2.47 135.0325 2.605 ;
         LAYER metal3 ;
         RECT  32.3175 57.5925 32.4525 57.7275 ;
         LAYER metal4 ;
         RECT  43.87 37.115 44.01 124.615 ;
         LAYER metal3 ;
         RECT  192.0975 2.47 192.2325 2.605 ;
         LAYER metal3 ;
         RECT  32.3175 41.2125 32.4525 41.3475 ;
         LAYER metal4 ;
         RECT  0.6875 24.0825 0.8275 46.485 ;
         LAYER metal3 ;
         RECT  237.8575 2.47 237.9925 2.605 ;
         LAYER metal4 ;
         RECT  105.195 34.205 105.335 125.91 ;
         LAYER metal3 ;
         RECT  260.7375 2.47 260.8725 2.605 ;
         LAYER metal3 ;
         RECT  146.3375 2.47 146.4725 2.605 ;
         LAYER metal3 ;
         RECT  44.8825 21.7175 45.0175 21.8525 ;
         LAYER metal3 ;
         RECT  77.6975 2.47 77.8325 2.605 ;
         LAYER metal3 ;
         RECT  54.8175 2.47 54.9525 2.605 ;
         LAYER metal4 ;
         RECT  44.95 34.205 45.09 125.91 ;
         LAYER metal4 ;
         RECT  37.87 37.115 38.01 124.685 ;
         LAYER metal3 ;
         RECT  43.3775 2.47 43.5125 2.605 ;
         LAYER metal3 ;
         RECT  214.9775 2.47 215.1125 2.605 ;
         LAYER metal4 ;
         RECT  26.215 58.955 26.355 73.915 ;
         LAYER metal3 ;
         RECT  45.0175 29.6125 103.7625 29.6825 ;
         LAYER metal3 ;
         RECT  89.1375 2.47 89.2725 2.605 ;
         LAYER metal3 ;
         RECT  100.5775 2.47 100.7125 2.605 ;
         LAYER metal3 ;
         RECT  45.0175 33.51 103.7625 33.58 ;
         LAYER metal3 ;
         RECT  32.3175 49.4025 32.4525 49.5375 ;
         LAYER metal3 ;
         RECT  31.9375 2.47 32.0725 2.605 ;
         LAYER metal3 ;
         RECT  32.3175 46.6725 32.4525 46.8075 ;
         LAYER metal3 ;
         RECT  66.2575 2.47 66.3925 2.605 ;
         LAYER metal3 ;
         RECT  180.6575 2.47 180.7925 2.605 ;
         LAYER metal4 ;
         RECT  28.935 16.705 29.075 31.665 ;
         LAYER metal3 ;
         RECT  226.4175 2.47 226.5525 2.605 ;
         LAYER metal3 ;
         RECT  123.4575 2.47 123.5925 2.605 ;
         LAYER metal3 ;
         RECT  157.7775 2.47 157.9125 2.605 ;
         LAYER metal3 ;
         RECT  203.5375 2.47 203.6725 2.605 ;
         LAYER metal3 ;
         RECT  43.8725 35.7525 44.0075 35.8875 ;
         LAYER metal3 ;
         RECT  32.3175 38.4825 32.4525 38.6175 ;
         LAYER metal3 ;
         RECT  103.6275 21.7175 103.7625 21.8525 ;
         LAYER metal3 ;
         RECT  38.49 36.41 38.625 36.545 ;
         LAYER metal3 ;
         RECT  32.3175 54.8625 32.4525 54.9975 ;
         LAYER metal3 ;
         RECT  45.0175 22.685 103.7625 22.755 ;
         LAYER metal3 ;
         RECT  112.0175 2.47 112.1525 2.605 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  252.1575 0.0 252.2925 0.135 ;
         LAYER metal4 ;
         RECT  29.075 58.89 29.215 73.98 ;
         LAYER metal3 ;
         RECT  229.2775 0.0 229.4125 0.135 ;
         LAYER metal3 ;
         RECT  30.79 56.2275 30.925 56.3625 ;
         LAYER metal3 ;
         RECT  30.79 48.0375 30.925 48.1725 ;
         LAYER metal3 ;
         RECT  263.5975 0.0 263.7325 0.135 ;
         LAYER metal3 ;
         RECT  217.8375 0.0 217.9725 0.135 ;
         LAYER metal3 ;
         RECT  103.4375 0.0 103.5725 0.135 ;
         LAYER metal4 ;
         RECT  2.75 24.115 2.89 46.5175 ;
         LAYER metal3 ;
         RECT  240.7175 0.0 240.8525 0.135 ;
         LAYER metal4 ;
         RECT  4.845 14.17 4.985 19.38 ;
         LAYER metal3 ;
         RECT  160.6375 0.0 160.7725 0.135 ;
         LAYER metal3 ;
         RECT  194.9575 0.0 195.0925 0.135 ;
         LAYER metal3 ;
         RECT  30.79 50.7675 30.925 50.9025 ;
         LAYER metal3 ;
         RECT  172.0775 0.0 172.2125 0.135 ;
         LAYER metal4 ;
         RECT  38.43 37.0825 38.57 124.6475 ;
         LAYER metal4 ;
         RECT  104.735 34.205 104.875 125.91 ;
         LAYER metal3 ;
         RECT  46.2375 0.0 46.3725 0.135 ;
         LAYER metal3 ;
         RECT  30.79 39.8475 30.925 39.9825 ;
         LAYER metal3 ;
         RECT  44.8825 19.8975 45.0175 20.0325 ;
         LAYER metal3 ;
         RECT  34.7975 0.0 34.9325 0.135 ;
         LAYER metal3 ;
         RECT  57.6775 0.0 57.8125 0.135 ;
         LAYER metal3 ;
         RECT  30.79 45.3075 30.925 45.4425 ;
         LAYER metal3 ;
         RECT  149.1975 0.0 149.3325 0.135 ;
         LAYER metal4 ;
         RECT  6.385 14.235 6.525 34.135 ;
         LAYER metal3 ;
         RECT  183.5175 0.0 183.6525 0.135 ;
         LAYER metal3 ;
         RECT  45.0175 24.735 103.7625 24.805 ;
         LAYER metal4 ;
         RECT  45.41 34.205 45.55 125.91 ;
         LAYER metal3 ;
         RECT  103.6275 19.8975 103.7625 20.0325 ;
         LAYER metal3 ;
         RECT  126.3175 0.0 126.4525 0.135 ;
         LAYER metal3 ;
         RECT  30.79 58.9575 30.925 59.0925 ;
         LAYER metal3 ;
         RECT  45.0175 31.505 103.7975 31.575 ;
         LAYER metal3 ;
         RECT  137.7575 0.0 137.8925 0.135 ;
         LAYER metal3 ;
         RECT  30.79 37.1175 30.925 37.2525 ;
         LAYER metal3 ;
         RECT  30.79 42.5775 30.925 42.7125 ;
         LAYER metal3 ;
         RECT  206.3975 0.0 206.5325 0.135 ;
         LAYER metal3 ;
         RECT  69.1175 0.0 69.2525 0.135 ;
         LAYER metal3 ;
         RECT  91.9975 0.0 92.1325 0.135 ;
         LAYER metal3 ;
         RECT  80.5575 0.0 80.6925 0.135 ;
         LAYER metal3 ;
         RECT  30.79 53.4975 30.925 53.6325 ;
         LAYER metal4 ;
         RECT  35.935 37.0825 36.075 124.685 ;
         LAYER metal3 ;
         RECT  114.8775 0.0 115.0125 0.135 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 272.105 125.9675 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 272.105 125.9675 ;
   LAYER  metal3 ;
      RECT  43.52 0.14 43.935 0.965 ;
      RECT  43.935 0.965 46.38 1.38 ;
      RECT  46.795 0.965 49.24 1.38 ;
      RECT  49.655 0.965 52.1 1.38 ;
      RECT  52.515 0.965 54.96 1.38 ;
      RECT  55.375 0.965 57.82 1.38 ;
      RECT  58.235 0.965 60.68 1.38 ;
      RECT  61.095 0.965 63.54 1.38 ;
      RECT  63.955 0.965 66.4 1.38 ;
      RECT  66.815 0.965 69.26 1.38 ;
      RECT  69.675 0.965 72.12 1.38 ;
      RECT  72.535 0.965 74.98 1.38 ;
      RECT  75.395 0.965 77.84 1.38 ;
      RECT  78.255 0.965 80.7 1.38 ;
      RECT  81.115 0.965 83.56 1.38 ;
      RECT  83.975 0.965 86.42 1.38 ;
      RECT  86.835 0.965 89.28 1.38 ;
      RECT  89.695 0.965 92.14 1.38 ;
      RECT  92.555 0.965 95.0 1.38 ;
      RECT  95.415 0.965 97.86 1.38 ;
      RECT  98.275 0.965 100.72 1.38 ;
      RECT  101.135 0.965 103.58 1.38 ;
      RECT  103.995 0.965 106.44 1.38 ;
      RECT  106.855 0.965 109.3 1.38 ;
      RECT  109.715 0.965 112.16 1.38 ;
      RECT  112.575 0.965 115.02 1.38 ;
      RECT  115.435 0.965 117.88 1.38 ;
      RECT  118.295 0.965 120.74 1.38 ;
      RECT  121.155 0.965 123.6 1.38 ;
      RECT  124.015 0.965 126.46 1.38 ;
      RECT  126.875 0.965 129.32 1.38 ;
      RECT  129.735 0.965 132.18 1.38 ;
      RECT  132.595 0.965 135.04 1.38 ;
      RECT  135.455 0.965 137.9 1.38 ;
      RECT  138.315 0.965 140.76 1.38 ;
      RECT  141.175 0.965 143.62 1.38 ;
      RECT  144.035 0.965 146.48 1.38 ;
      RECT  146.895 0.965 149.34 1.38 ;
      RECT  149.755 0.965 152.2 1.38 ;
      RECT  152.615 0.965 155.06 1.38 ;
      RECT  155.475 0.965 157.92 1.38 ;
      RECT  158.335 0.965 160.78 1.38 ;
      RECT  161.195 0.965 163.64 1.38 ;
      RECT  164.055 0.965 166.5 1.38 ;
      RECT  166.915 0.965 169.36 1.38 ;
      RECT  169.775 0.965 172.22 1.38 ;
      RECT  172.635 0.965 175.08 1.38 ;
      RECT  175.495 0.965 177.94 1.38 ;
      RECT  178.355 0.965 180.8 1.38 ;
      RECT  181.215 0.965 183.66 1.38 ;
      RECT  184.075 0.965 186.52 1.38 ;
      RECT  186.935 0.965 189.38 1.38 ;
      RECT  189.795 0.965 192.24 1.38 ;
      RECT  192.655 0.965 195.1 1.38 ;
      RECT  195.515 0.965 197.96 1.38 ;
      RECT  198.375 0.965 200.82 1.38 ;
      RECT  201.235 0.965 203.68 1.38 ;
      RECT  204.095 0.965 206.54 1.38 ;
      RECT  206.955 0.965 209.4 1.38 ;
      RECT  209.815 0.965 212.26 1.38 ;
      RECT  212.675 0.965 215.12 1.38 ;
      RECT  215.535 0.965 217.98 1.38 ;
      RECT  218.395 0.965 220.84 1.38 ;
      RECT  221.255 0.965 223.7 1.38 ;
      RECT  224.115 0.965 226.56 1.38 ;
      RECT  226.975 0.965 229.42 1.38 ;
      RECT  229.835 0.965 232.28 1.38 ;
      RECT  232.695 0.965 235.14 1.38 ;
      RECT  235.555 0.965 238.0 1.38 ;
      RECT  238.415 0.965 240.86 1.38 ;
      RECT  241.275 0.965 243.72 1.38 ;
      RECT  244.135 0.965 246.58 1.38 ;
      RECT  246.995 0.965 249.44 1.38 ;
      RECT  249.855 0.965 252.3 1.38 ;
      RECT  252.715 0.965 255.16 1.38 ;
      RECT  255.575 0.965 258.02 1.38 ;
      RECT  258.435 0.965 260.88 1.38 ;
      RECT  261.295 0.965 263.74 1.38 ;
      RECT  264.155 0.965 266.6 1.38 ;
      RECT  267.015 0.965 269.46 1.38 ;
      RECT  269.875 0.965 272.105 1.38 ;
      RECT  0.14 59.9225 26.36 60.3375 ;
      RECT  0.14 60.3375 26.36 125.9675 ;
      RECT  26.36 1.38 26.775 59.9225 ;
      RECT  26.775 59.9225 43.52 60.3375 ;
      RECT  26.775 60.3375 43.52 125.9675 ;
      RECT  26.36 60.3375 26.775 62.6525 ;
      RECT  26.36 63.0675 26.775 64.8625 ;
      RECT  26.36 65.2775 26.775 67.5925 ;
      RECT  26.36 68.0075 26.775 69.8025 ;
      RECT  26.36 70.2175 26.775 72.5325 ;
      RECT  26.36 72.9475 26.775 125.9675 ;
      RECT  0.14 1.38 0.145 15.2025 ;
      RECT  0.14 15.2025 0.145 15.6175 ;
      RECT  0.14 15.6175 0.145 59.9225 ;
      RECT  0.145 1.38 0.56 15.2025 ;
      RECT  0.56 1.38 26.36 15.2025 ;
      RECT  0.145 15.6175 0.56 17.9325 ;
      RECT  0.145 18.3475 0.56 59.9225 ;
      RECT  0.56 15.2025 6.3875 15.2875 ;
      RECT  0.56 15.2875 6.3875 15.6175 ;
      RECT  6.3875 15.2025 6.8025 15.2875 ;
      RECT  6.8025 15.2025 26.36 15.2875 ;
      RECT  6.8025 15.2875 26.36 15.6175 ;
      RECT  0.56 15.6175 6.3875 15.7025 ;
      RECT  0.56 15.7025 6.3875 59.9225 ;
      RECT  6.3875 15.7025 6.8025 59.9225 ;
      RECT  6.8025 15.6175 26.36 15.7025 ;
      RECT  6.8025 15.7025 26.36 59.9225 ;
      RECT  0.14 0.965 32.08 1.38 ;
      RECT  32.495 0.965 34.94 1.38 ;
      RECT  35.355 0.965 37.8 1.38 ;
      RECT  38.215 0.965 40.66 1.38 ;
      RECT  41.075 0.965 43.52 1.38 ;
      RECT  43.935 26.8525 47.1225 27.2675 ;
      RECT  47.5375 26.8525 47.8275 27.2675 ;
      RECT  48.2425 26.8525 48.5325 27.2675 ;
      RECT  48.9475 26.8525 49.2375 27.2675 ;
      RECT  49.6525 26.8525 49.9425 27.2675 ;
      RECT  50.3575 26.8525 50.6475 27.2675 ;
      RECT  51.0625 26.8525 51.3525 27.2675 ;
      RECT  51.7675 26.8525 52.0575 27.2675 ;
      RECT  52.4725 26.8525 52.7625 27.2675 ;
      RECT  53.1775 26.8525 53.4675 27.2675 ;
      RECT  53.8825 26.8525 54.1725 27.2675 ;
      RECT  54.5875 26.8525 54.8775 27.2675 ;
      RECT  55.2925 26.8525 55.5825 27.2675 ;
      RECT  55.9975 26.8525 56.2875 27.2675 ;
      RECT  56.7025 26.8525 56.9925 27.2675 ;
      RECT  57.4075 26.8525 57.6975 27.2675 ;
      RECT  58.1125 26.8525 58.4025 27.2675 ;
      RECT  58.8175 26.8525 59.1075 27.2675 ;
      RECT  59.5225 26.8525 59.8125 27.2675 ;
      RECT  60.2275 26.8525 60.5175 27.2675 ;
      RECT  60.9325 26.8525 61.2225 27.2675 ;
      RECT  61.6375 26.8525 61.9275 27.2675 ;
      RECT  62.3425 26.8525 62.6325 27.2675 ;
      RECT  63.0475 26.8525 63.3375 27.2675 ;
      RECT  63.7525 26.8525 64.0425 27.2675 ;
      RECT  64.4575 26.8525 64.7475 27.2675 ;
      RECT  65.1625 26.8525 65.4525 27.2675 ;
      RECT  65.8675 26.8525 66.1575 27.2675 ;
      RECT  66.5725 26.8525 66.8625 27.2675 ;
      RECT  67.2775 26.8525 67.5675 27.2675 ;
      RECT  67.9825 26.8525 68.2725 27.2675 ;
      RECT  68.6875 26.8525 68.9775 27.2675 ;
      RECT  69.3925 26.8525 69.6825 27.2675 ;
      RECT  70.0975 26.8525 70.3875 27.2675 ;
      RECT  70.8025 26.8525 71.0925 27.2675 ;
      RECT  71.5075 26.8525 71.7975 27.2675 ;
      RECT  72.2125 26.8525 72.5025 27.2675 ;
      RECT  72.9175 26.8525 73.2075 27.2675 ;
      RECT  73.6225 26.8525 73.9125 27.2675 ;
      RECT  74.3275 26.8525 74.6175 27.2675 ;
      RECT  75.0325 26.8525 75.3225 27.2675 ;
      RECT  75.7375 26.8525 76.0275 27.2675 ;
      RECT  76.4425 26.8525 76.7325 27.2675 ;
      RECT  77.1475 26.8525 77.4375 27.2675 ;
      RECT  77.8525 26.8525 78.1425 27.2675 ;
      RECT  78.5575 26.8525 78.8475 27.2675 ;
      RECT  79.2625 26.8525 79.5525 27.2675 ;
      RECT  79.9675 26.8525 80.2575 27.2675 ;
      RECT  80.6725 26.8525 80.9625 27.2675 ;
      RECT  81.3775 26.8525 81.6675 27.2675 ;
      RECT  82.0825 26.8525 82.3725 27.2675 ;
      RECT  82.7875 26.8525 83.0775 27.2675 ;
      RECT  83.4925 26.8525 83.7825 27.2675 ;
      RECT  84.1975 26.8525 84.4875 27.2675 ;
      RECT  84.9025 26.8525 85.1925 27.2675 ;
      RECT  85.6075 26.8525 85.8975 27.2675 ;
      RECT  86.3125 26.8525 86.6025 27.2675 ;
      RECT  87.0175 26.8525 87.3075 27.2675 ;
      RECT  87.7225 26.8525 88.0125 27.2675 ;
      RECT  88.4275 26.8525 88.7175 27.2675 ;
      RECT  89.1325 26.8525 89.4225 27.2675 ;
      RECT  89.8375 26.8525 90.1275 27.2675 ;
      RECT  90.5425 26.8525 90.8325 27.2675 ;
      RECT  91.2475 26.8525 91.5375 27.2675 ;
      RECT  91.9525 26.8525 92.2425 27.2675 ;
      RECT  92.6575 26.8525 92.9475 27.2675 ;
      RECT  93.3625 26.8525 93.6525 27.2675 ;
      RECT  94.0675 26.8525 94.3575 27.2675 ;
      RECT  94.7725 26.8525 95.0625 27.2675 ;
      RECT  95.4775 26.8525 95.7675 27.2675 ;
      RECT  96.1825 26.8525 96.4725 27.2675 ;
      RECT  96.8875 26.8525 97.1775 27.2675 ;
      RECT  97.5925 26.8525 97.8825 27.2675 ;
      RECT  98.2975 26.8525 98.5875 27.2675 ;
      RECT  99.0025 26.8525 99.2925 27.2675 ;
      RECT  99.7075 26.8525 99.9975 27.2675 ;
      RECT  100.4125 26.8525 100.7025 27.2675 ;
      RECT  101.1175 26.8525 101.4075 27.2675 ;
      RECT  101.8225 26.8525 102.1125 27.2675 ;
      RECT  102.5275 26.8525 102.8175 27.2675 ;
      RECT  103.2325 26.8525 272.105 27.2675 ;
      RECT  47.5375 1.38 249.1575 2.33 ;
      RECT  249.1575 1.38 249.5725 2.33 ;
      RECT  249.1575 2.745 249.5725 26.8525 ;
      RECT  249.5725 1.38 272.105 2.33 ;
      RECT  249.5725 2.745 272.105 26.8525 ;
      RECT  26.775 57.4525 32.1775 57.8675 ;
      RECT  32.1775 57.8675 32.5925 59.9225 ;
      RECT  32.5925 57.4525 43.52 57.8675 ;
      RECT  32.5925 57.8675 43.52 59.9225 ;
      RECT  238.1325 2.33 249.1575 2.745 ;
      RECT  249.5725 2.33 260.5975 2.745 ;
      RECT  261.0125 2.33 272.105 2.745 ;
      RECT  135.1725 2.33 146.1975 2.745 ;
      RECT  43.935 1.38 44.7425 21.5775 ;
      RECT  43.935 21.5775 44.7425 21.9925 ;
      RECT  43.935 21.9925 44.7425 26.8525 ;
      RECT  45.1575 1.38 47.1225 21.5775 ;
      RECT  45.1575 21.5775 47.1225 21.9925 ;
      RECT  47.5375 2.33 54.6775 2.745 ;
      RECT  43.52 1.38 43.6525 2.33 ;
      RECT  43.52 2.745 43.6525 125.9675 ;
      RECT  43.6525 1.38 43.935 2.33 ;
      RECT  43.6525 2.33 43.935 2.745 ;
      RECT  32.5925 1.38 43.2375 2.33 ;
      RECT  32.5925 2.33 43.2375 2.745 ;
      RECT  43.2375 1.38 43.52 2.33 ;
      RECT  43.2375 2.745 43.52 57.4525 ;
      RECT  43.935 27.2675 44.8775 29.4725 ;
      RECT  43.935 29.4725 44.8775 29.8225 ;
      RECT  44.8775 27.2675 47.1225 29.4725 ;
      RECT  47.1225 27.2675 47.5375 29.4725 ;
      RECT  47.5375 27.2675 103.9025 29.4725 ;
      RECT  103.9025 27.2675 272.105 29.4725 ;
      RECT  103.9025 29.4725 272.105 29.8225 ;
      RECT  77.9725 2.33 88.9975 2.745 ;
      RECT  89.4125 2.33 100.4375 2.745 ;
      RECT  44.8775 33.72 47.1225 125.9675 ;
      RECT  47.1225 33.72 47.5375 125.9675 ;
      RECT  47.5375 33.72 103.9025 125.9675 ;
      RECT  26.775 1.38 31.7975 2.33 ;
      RECT  26.775 2.33 31.7975 2.745 ;
      RECT  31.7975 1.38 32.1775 2.33 ;
      RECT  31.7975 2.745 32.1775 57.4525 ;
      RECT  32.1775 1.38 32.2125 2.33 ;
      RECT  32.2125 1.38 32.5925 2.33 ;
      RECT  32.2125 2.33 32.5925 2.745 ;
      RECT  32.1775 41.4875 32.5925 46.5325 ;
      RECT  32.1775 46.9475 32.5925 49.2625 ;
      RECT  55.0925 2.33 66.1175 2.745 ;
      RECT  66.5325 2.33 77.5575 2.745 ;
      RECT  169.4925 2.33 180.5175 2.745 ;
      RECT  180.9325 2.33 191.9575 2.745 ;
      RECT  215.2525 2.33 226.2775 2.745 ;
      RECT  226.6925 2.33 237.7175 2.745 ;
      RECT  123.7325 2.33 134.7575 2.745 ;
      RECT  146.6125 2.33 157.6375 2.745 ;
      RECT  158.0525 2.33 169.0775 2.745 ;
      RECT  192.3725 2.33 203.3975 2.745 ;
      RECT  203.8125 2.33 214.8375 2.745 ;
      RECT  43.6525 2.745 43.7325 35.6125 ;
      RECT  43.6525 35.6125 43.7325 36.0275 ;
      RECT  43.6525 36.0275 43.7325 125.9675 ;
      RECT  43.7325 2.745 43.935 35.6125 ;
      RECT  43.7325 36.0275 43.935 125.9675 ;
      RECT  43.935 29.8225 44.1475 35.6125 ;
      RECT  43.935 36.0275 44.1475 125.9675 ;
      RECT  44.1475 29.8225 44.8775 35.6125 ;
      RECT  44.1475 35.6125 44.8775 36.0275 ;
      RECT  44.1475 36.0275 44.8775 125.9675 ;
      RECT  32.1775 2.745 32.2125 38.3425 ;
      RECT  32.1775 38.7575 32.2125 41.0725 ;
      RECT  32.2125 2.745 32.5925 38.3425 ;
      RECT  32.2125 38.7575 32.5925 41.0725 ;
      RECT  47.5375 2.745 103.4875 21.5775 ;
      RECT  47.5375 21.5775 103.4875 21.9925 ;
      RECT  103.9025 2.745 249.1575 21.5775 ;
      RECT  103.9025 21.5775 249.1575 21.9925 ;
      RECT  103.9025 21.9925 249.1575 26.8525 ;
      RECT  32.5925 2.745 38.35 36.27 ;
      RECT  32.5925 36.27 38.35 36.685 ;
      RECT  32.5925 36.685 38.35 57.4525 ;
      RECT  38.35 2.745 38.765 36.27 ;
      RECT  38.35 36.685 38.765 57.4525 ;
      RECT  38.765 2.745 43.2375 36.27 ;
      RECT  38.765 36.27 43.2375 36.685 ;
      RECT  38.765 36.685 43.2375 57.4525 ;
      RECT  32.1775 49.6775 32.5925 54.7225 ;
      RECT  32.1775 55.1375 32.5925 57.4525 ;
      RECT  47.1225 1.38 47.5375 22.545 ;
      RECT  44.7425 21.9925 44.8775 22.545 ;
      RECT  44.7425 22.545 44.8775 22.895 ;
      RECT  44.7425 22.895 44.8775 26.8525 ;
      RECT  44.8775 21.9925 45.1575 22.545 ;
      RECT  45.1575 21.9925 47.1225 22.545 ;
      RECT  47.5375 21.9925 103.4875 22.545 ;
      RECT  103.4875 21.9925 103.9025 22.545 ;
      RECT  100.8525 2.33 111.8775 2.745 ;
      RECT  112.2925 2.33 123.3175 2.745 ;
      RECT  43.935 0.275 252.0175 0.965 ;
      RECT  252.0175 0.275 252.4325 0.965 ;
      RECT  252.4325 0.275 272.105 0.965 ;
      RECT  26.775 2.745 30.65 56.0875 ;
      RECT  26.775 56.0875 30.65 56.5025 ;
      RECT  26.775 56.5025 30.65 57.4525 ;
      RECT  30.65 56.5025 31.065 57.4525 ;
      RECT  31.065 2.745 31.7975 56.0875 ;
      RECT  31.065 56.0875 31.7975 56.5025 ;
      RECT  31.065 56.5025 31.7975 57.4525 ;
      RECT  252.4325 0.14 263.4575 0.275 ;
      RECT  263.8725 0.14 272.105 0.275 ;
      RECT  218.1125 0.14 229.1375 0.275 ;
      RECT  229.5525 0.14 240.5775 0.275 ;
      RECT  240.9925 0.14 252.0175 0.275 ;
      RECT  30.65 48.3125 31.065 50.6275 ;
      RECT  160.9125 0.14 171.9375 0.275 ;
      RECT  43.935 0.14 46.0975 0.275 ;
      RECT  44.7425 1.38 45.1575 19.7575 ;
      RECT  44.7425 20.1725 45.1575 21.5775 ;
      RECT  0.14 0.14 34.6575 0.275 ;
      RECT  0.14 0.275 34.6575 0.965 ;
      RECT  34.6575 0.275 35.0725 0.965 ;
      RECT  35.0725 0.14 43.52 0.275 ;
      RECT  35.0725 0.275 43.52 0.965 ;
      RECT  46.5125 0.14 57.5375 0.275 ;
      RECT  30.65 45.5825 31.065 47.8975 ;
      RECT  149.4725 0.14 160.4975 0.275 ;
      RECT  172.3525 0.14 183.3775 0.275 ;
      RECT  183.7925 0.14 194.8175 0.275 ;
      RECT  47.1225 22.895 47.5375 24.595 ;
      RECT  47.1225 24.945 47.5375 26.8525 ;
      RECT  44.8775 22.895 45.1575 24.595 ;
      RECT  44.8775 24.945 45.1575 26.8525 ;
      RECT  45.1575 22.895 47.1225 24.595 ;
      RECT  45.1575 24.945 47.1225 26.8525 ;
      RECT  47.5375 22.895 103.4875 24.595 ;
      RECT  47.5375 24.945 103.4875 26.8525 ;
      RECT  103.4875 22.895 103.9025 24.595 ;
      RECT  103.4875 24.945 103.9025 26.8525 ;
      RECT  103.4875 2.745 103.9025 19.7575 ;
      RECT  103.4875 20.1725 103.9025 21.5775 ;
      RECT  26.775 57.8675 30.65 58.8175 ;
      RECT  26.775 58.8175 30.65 59.2325 ;
      RECT  26.775 59.2325 30.65 59.9225 ;
      RECT  30.65 57.8675 31.065 58.8175 ;
      RECT  30.65 59.2325 31.065 59.9225 ;
      RECT  31.065 57.8675 32.1775 58.8175 ;
      RECT  31.065 58.8175 32.1775 59.2325 ;
      RECT  31.065 59.2325 32.1775 59.9225 ;
      RECT  103.9025 29.8225 103.9375 31.365 ;
      RECT  103.9025 31.715 103.9375 125.9675 ;
      RECT  103.9375 29.8225 272.105 31.365 ;
      RECT  103.9375 31.365 272.105 31.715 ;
      RECT  103.9375 31.715 272.105 125.9675 ;
      RECT  44.8775 29.8225 47.1225 31.365 ;
      RECT  44.8775 31.715 47.1225 33.37 ;
      RECT  47.1225 29.8225 47.5375 31.365 ;
      RECT  47.1225 31.715 47.5375 33.37 ;
      RECT  47.5375 29.8225 103.9025 31.365 ;
      RECT  47.5375 31.715 103.9025 33.37 ;
      RECT  126.5925 0.14 137.6175 0.275 ;
      RECT  138.0325 0.14 149.0575 0.275 ;
      RECT  30.65 2.745 31.065 36.9775 ;
      RECT  30.65 37.3925 31.065 39.7075 ;
      RECT  30.65 40.1225 31.065 42.4375 ;
      RECT  30.65 42.8525 31.065 45.1675 ;
      RECT  195.2325 0.14 206.2575 0.275 ;
      RECT  206.6725 0.14 217.6975 0.275 ;
      RECT  57.9525 0.14 68.9775 0.275 ;
      RECT  92.2725 0.14 103.2975 0.275 ;
      RECT  69.3925 0.14 80.4175 0.275 ;
      RECT  80.8325 0.14 91.8575 0.275 ;
      RECT  30.65 51.0425 31.065 53.3575 ;
      RECT  30.65 53.7725 31.065 56.0875 ;
      RECT  103.7125 0.14 114.7375 0.275 ;
      RECT  115.1525 0.14 126.1775 0.275 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 0.42 13.955 ;
      RECT  43.59 19.595 44.29 36.835 ;
      RECT  43.59 124.895 44.29 125.9675 ;
      RECT  0.14 19.595 0.4075 23.8025 ;
      RECT  0.14 23.8025 0.4075 46.765 ;
      RECT  0.14 46.765 0.4075 125.9675 ;
      RECT  0.4075 19.595 0.42 23.8025 ;
      RECT  0.4075 46.765 0.42 125.9675 ;
      RECT  0.42 19.595 1.1075 23.8025 ;
      RECT  0.42 46.765 1.1075 124.895 ;
      RECT  44.29 19.595 104.915 33.925 ;
      RECT  104.915 19.595 105.615 33.925 ;
      RECT  105.615 19.595 272.105 33.925 ;
      RECT  105.615 33.925 272.105 36.835 ;
      RECT  105.615 36.835 272.105 124.895 ;
      RECT  105.615 124.895 272.105 125.9675 ;
      RECT  44.29 33.925 44.67 36.835 ;
      RECT  44.29 36.835 44.67 124.895 ;
      RECT  44.29 124.895 44.67 125.9675 ;
      RECT  0.42 124.965 37.59 125.9675 ;
      RECT  37.59 124.965 38.29 125.9675 ;
      RECT  38.29 124.965 43.59 125.9675 ;
      RECT  1.1075 58.675 25.935 74.195 ;
      RECT  1.1075 74.195 25.935 124.895 ;
      RECT  25.935 46.765 26.635 58.675 ;
      RECT  25.935 74.195 26.635 124.895 ;
      RECT  28.655 13.955 29.355 16.425 ;
      RECT  29.355 13.955 272.105 16.425 ;
      RECT  29.355 16.425 272.105 19.595 ;
      RECT  29.355 19.595 43.59 23.8025 ;
      RECT  28.655 31.945 29.355 36.835 ;
      RECT  29.355 23.8025 43.59 31.945 ;
      RECT  26.635 46.765 28.795 58.61 ;
      RECT  26.635 58.61 28.795 58.675 ;
      RECT  28.795 46.765 29.495 58.61 ;
      RECT  26.635 58.675 28.795 74.195 ;
      RECT  26.635 74.195 28.795 74.26 ;
      RECT  26.635 74.26 28.795 124.895 ;
      RECT  28.795 74.26 29.495 124.895 ;
      RECT  1.1075 36.835 2.47 46.765 ;
      RECT  1.1075 46.765 2.47 46.7975 ;
      RECT  1.1075 46.7975 2.47 58.675 ;
      RECT  2.47 46.7975 3.17 58.675 ;
      RECT  3.17 46.765 25.935 46.7975 ;
      RECT  3.17 46.7975 25.935 58.675 ;
      RECT  1.1075 23.8025 2.47 23.835 ;
      RECT  1.1075 23.835 2.47 31.945 ;
      RECT  2.47 23.8025 3.17 23.835 ;
      RECT  1.1075 31.945 2.47 36.835 ;
      RECT  0.42 0.14 4.565 13.89 ;
      RECT  0.42 13.89 4.565 13.955 ;
      RECT  4.565 0.14 5.265 13.89 ;
      RECT  5.265 0.14 272.105 13.89 ;
      RECT  5.265 13.89 272.105 13.955 ;
      RECT  0.42 13.955 4.565 16.425 ;
      RECT  0.42 16.425 4.565 19.595 ;
      RECT  1.1075 19.595 4.565 19.66 ;
      RECT  1.1075 19.66 4.565 23.8025 ;
      RECT  4.565 19.66 5.265 23.8025 ;
      RECT  38.29 124.9275 38.85 124.965 ;
      RECT  38.85 124.895 43.59 124.9275 ;
      RECT  38.85 124.9275 43.59 124.965 ;
      RECT  38.85 36.835 43.59 46.765 ;
      RECT  38.85 46.765 43.59 124.895 ;
      RECT  29.355 31.945 38.15 36.8025 ;
      RECT  38.15 31.945 38.85 36.8025 ;
      RECT  38.85 31.945 43.59 36.8025 ;
      RECT  38.85 36.8025 43.59 36.835 ;
      RECT  3.17 23.8025 6.105 23.835 ;
      RECT  6.805 23.8025 28.655 23.835 ;
      RECT  3.17 23.835 6.105 31.945 ;
      RECT  6.805 23.835 28.655 31.945 ;
      RECT  3.17 31.945 6.105 34.415 ;
      RECT  3.17 34.415 6.105 36.835 ;
      RECT  6.105 34.415 6.805 36.835 ;
      RECT  6.805 31.945 28.655 34.415 ;
      RECT  6.805 34.415 28.655 36.835 ;
      RECT  5.265 13.955 6.105 16.425 ;
      RECT  6.805 13.955 28.655 16.425 ;
      RECT  5.265 16.425 6.105 19.595 ;
      RECT  6.805 16.425 28.655 19.595 ;
      RECT  5.265 19.595 6.105 19.66 ;
      RECT  6.805 19.595 28.655 19.66 ;
      RECT  5.265 19.66 6.105 23.8025 ;
      RECT  6.805 19.66 28.655 23.8025 ;
      RECT  45.83 33.925 104.455 36.835 ;
      RECT  45.83 36.835 104.455 124.895 ;
      RECT  45.83 124.895 104.455 125.9675 ;
      RECT  0.42 124.895 35.655 124.965 ;
      RECT  36.355 124.895 37.59 124.965 ;
      RECT  29.495 46.765 35.655 58.61 ;
      RECT  36.355 46.765 37.59 58.61 ;
      RECT  29.495 58.61 35.655 58.675 ;
      RECT  36.355 58.61 37.59 58.675 ;
      RECT  29.495 58.675 35.655 74.195 ;
      RECT  36.355 58.675 37.59 74.195 ;
      RECT  29.495 74.195 35.655 74.26 ;
      RECT  36.355 74.195 37.59 74.26 ;
      RECT  29.495 74.26 35.655 124.895 ;
      RECT  36.355 74.26 37.59 124.895 ;
      RECT  3.17 36.835 35.655 46.765 ;
      RECT  36.355 36.835 37.59 46.765 ;
      RECT  29.355 36.8025 35.655 36.835 ;
      RECT  36.355 36.8025 38.15 36.835 ;
   END
END    freepdk45_sram_1rw0r_64x80_20
END    LIBRARY
