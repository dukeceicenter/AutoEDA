../macros/freepdk45_sram_1w1r_40x128/freepdk45_sram_1w1r_40x128.lef