VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_16x32_32
   CLASS BLOCK ;
   SIZE 111.97 BY 62.75 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.665 1.1075 20.8 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.525 1.1075 23.66 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.385 1.1075 26.52 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.245 1.1075 29.38 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.105 1.1075 32.24 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.965 1.1075 35.1 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.825 1.1075 37.96 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.685 1.1075 40.82 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.545 1.1075 43.68 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.405 1.1075 46.54 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.265 1.1075 49.4 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.125 1.1075 52.26 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.985 1.1075 55.12 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.845 1.1075 57.98 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.705 1.1075 60.84 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.565 1.1075 63.7 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.425 1.1075 66.56 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.285 1.1075 69.42 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.145 1.1075 72.28 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.005 1.1075 75.14 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.865 1.1075 78.0 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.725 1.1075 80.86 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.585 1.1075 83.72 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.445 1.1075 86.58 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.305 1.1075 89.44 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.165 1.1075 92.3 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.025 1.1075 95.16 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.885 1.1075 98.02 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.745 1.1075 100.88 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.605 1.1075 103.74 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.465 1.1075 106.6 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.325 1.1075 109.46 1.2425 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14.945 36.7275 15.08 36.8625 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14.945 39.4575 15.08 39.5925 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14.945 41.6675 15.08 41.8025 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14.945 44.3975 15.08 44.5325 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.205 19.5675 88.34 19.7025 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.205 16.8375 88.34 16.9725 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.205 14.6275 88.34 14.7625 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.205 11.8975 88.34 12.0325 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.005 61.5075 103.14 61.6425 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.9025 61.4225 97.0375 61.5575 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.7125 54.8 32.8475 54.935 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.8875 54.8 34.0225 54.935 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.0625 54.8 35.1975 54.935 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.2375 54.8 36.3725 54.935 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.4125 54.8 37.5475 54.935 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.5875 54.8 38.7225 54.935 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.7625 54.8 39.8975 54.935 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.9375 54.8 41.0725 54.935 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.1125 54.8 42.2475 54.935 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.2875 54.8 43.4225 54.935 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.4625 54.8 44.5975 54.935 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.6375 54.8 45.7725 54.935 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.8125 54.8 46.9475 54.935 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.9875 54.8 48.1225 54.935 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.1625 54.8 49.2975 54.935 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.3375 54.8 50.4725 54.935 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.5125 54.8 51.6475 54.935 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.6875 54.8 52.8225 54.935 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.8625 54.8 53.9975 54.935 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.0375 54.8 55.1725 54.935 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.2125 54.8 56.3475 54.935 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.3875 54.8 57.5225 54.935 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.5625 54.8 58.6975 54.935 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.7375 54.8 59.8725 54.935 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.9125 54.8 61.0475 54.935 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.0875 54.8 62.2225 54.935 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.2625 54.8 63.3975 54.935 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.4375 54.8 64.5725 54.935 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.6125 54.8 65.7475 54.935 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.7875 54.8 66.9225 54.935 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.9625 54.8 68.0975 54.935 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.1375 54.8 69.2725 54.935 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  82.4725 25.1575 82.6075 25.2925 ;
         LAYER metal3 ;
         RECT  77.205 45.3 77.34 45.435 ;
         LAYER metal3 ;
         RECT  29.5275 48.345 71.5875 48.415 ;
         LAYER metal3 ;
         RECT  43.2625 2.4725 43.3975 2.6075 ;
         LAYER metal3 ;
         RECT  66.1425 2.4725 66.2775 2.6075 ;
         LAYER metal4 ;
         RECT  74.57 20.67 74.71 44.73 ;
         LAYER metal3 ;
         RECT  82.4725 22.1675 82.6075 22.3025 ;
         LAYER metal3 ;
         RECT  20.4825 22.1675 20.6175 22.3025 ;
         LAYER metal4 ;
         RECT  17.38 2.47 17.52 17.43 ;
         LAYER metal4 ;
         RECT  25.13 20.67 25.27 44.8 ;
         LAYER metal3 ;
         RECT  54.7025 2.4725 54.8375 2.6075 ;
         LAYER metal3 ;
         RECT  82.4725 34.1275 82.6075 34.2625 ;
         LAYER metal3 ;
         RECT  74.5725 46.0875 74.7075 46.2225 ;
         LAYER metal3 ;
         RECT  20.4825 34.1275 20.6175 34.2625 ;
         LAYER metal3 ;
         RECT  100.4625 2.4725 100.5975 2.6075 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
         LAYER metal3 ;
         RECT  20.4825 31.1375 20.6175 31.2725 ;
         LAYER metal3 ;
         RECT  25.75 19.965 25.885 20.1 ;
         LAYER metal3 ;
         RECT  20.4825 25.1575 20.6175 25.2925 ;
         LAYER metal3 ;
         RECT  29.5275 52.2425 69.9425 52.3125 ;
         LAYER metal3 ;
         RECT  29.5275 16.805 70.4125 16.875 ;
         LAYER metal4 ;
         RECT  77.82 20.67 77.96 44.8 ;
         LAYER metal3 ;
         RECT  89.0225 2.4725 89.1575 2.6075 ;
         LAYER metal4 ;
         RECT  85.765 50.26 85.905 60.28 ;
         LAYER metal3 ;
         RECT  20.3825 2.4725 20.5175 2.6075 ;
         LAYER metal3 ;
         RECT  77.5825 2.4725 77.7175 2.6075 ;
         LAYER metal3 ;
         RECT  29.5275 11.37 69.9425 11.44 ;
         LAYER metal4 ;
         RECT  28.38 20.67 28.52 44.73 ;
         LAYER metal4 ;
         RECT  29.46 17.5 29.6 47.65 ;
         LAYER metal3 ;
         RECT  82.4725 31.1375 82.6075 31.2725 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal3 ;
         RECT  100.865 60.1425 101.0 60.2775 ;
         LAYER metal4 ;
         RECT  102.5975 30.5 102.7375 52.9025 ;
         LAYER metal4 ;
         RECT  14.66 35.62 14.8 45.64 ;
         LAYER metal4 ;
         RECT  88.485 10.79 88.625 20.81 ;
         LAYER metal3 ;
         RECT  28.3825 19.1775 28.5175 19.3125 ;
         LAYER metal4 ;
         RECT  73.49 17.5 73.63 47.65 ;
         LAYER metal3 ;
         RECT  31.8225 2.4725 31.9575 2.6075 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  91.8825 0.0025 92.0175 0.1375 ;
         LAYER metal3 ;
         RECT  69.0025 0.0025 69.1375 0.1375 ;
         LAYER metal4 ;
         RECT  100.535 30.4675 100.675 52.87 ;
         LAYER metal3 ;
         RECT  23.2425 0.0025 23.3775 0.1375 ;
         LAYER metal4 ;
         RECT  23.54 20.6375 23.68 44.8 ;
         LAYER metal3 ;
         RECT  84.0 23.6625 84.135 23.7975 ;
         LAYER metal4 ;
         RECT  77.26 20.6375 77.4 44.7625 ;
         LAYER metal4 ;
         RECT  73.03 17.5 73.17 47.65 ;
         LAYER metal3 ;
         RECT  84.0 35.6225 84.135 35.7575 ;
         LAYER metal3 ;
         RECT  18.955 23.6625 19.09 23.7975 ;
         LAYER metal3 ;
         RECT  100.865 62.6125 101.0 62.7475 ;
         LAYER metal3 ;
         RECT  84.0 26.6525 84.135 26.7875 ;
         LAYER metal3 ;
         RECT  18.955 26.6525 19.09 26.7875 ;
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal3 ;
         RECT  18.955 29.6425 19.09 29.7775 ;
         LAYER metal3 ;
         RECT  29.5275 50.35 69.9775 50.42 ;
         LAYER metal3 ;
         RECT  84.0 29.6425 84.135 29.7775 ;
         LAYER metal4 ;
         RECT  85.625 10.725 85.765 20.875 ;
         LAYER metal4 ;
         RECT  97.04 47.79 97.18 62.75 ;
         LAYER metal4 ;
         RECT  17.52 35.555 17.66 45.705 ;
         LAYER metal3 ;
         RECT  57.5625 0.0025 57.6975 0.1375 ;
         LAYER metal3 ;
         RECT  46.1225 0.0025 46.2575 0.1375 ;
         LAYER metal3 ;
         RECT  84.0 20.6725 84.135 20.8075 ;
         LAYER metal3 ;
         RECT  18.955 32.6325 19.09 32.7675 ;
         LAYER metal3 ;
         RECT  84.0 32.6325 84.135 32.7675 ;
         LAYER metal4 ;
         RECT  25.69 20.6375 25.83 44.7625 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal3 ;
         RECT  103.3225 0.0025 103.4575 0.1375 ;
         LAYER metal3 ;
         RECT  80.4425 0.0025 80.5775 0.1375 ;
         LAYER metal3 ;
         RECT  18.955 20.6725 19.09 20.8075 ;
         LAYER metal4 ;
         RECT  79.41 20.6375 79.55 44.8 ;
         LAYER metal4 ;
         RECT  29.92 17.5 30.06 47.65 ;
         LAYER metal3 ;
         RECT  18.955 35.6225 19.09 35.7575 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal3 ;
         RECT  34.6825 0.0025 34.8175 0.1375 ;
         LAYER metal3 ;
         RECT  29.5275 13.42 69.9425 13.49 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 111.83 62.61 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 111.83 62.61 ;
   LAYER  metal3 ;
      RECT  20.525 0.14 20.94 0.9675 ;
      RECT  20.94 0.9675 23.385 1.3825 ;
      RECT  23.8 0.9675 26.245 1.3825 ;
      RECT  26.66 0.9675 29.105 1.3825 ;
      RECT  29.52 0.9675 31.965 1.3825 ;
      RECT  32.38 0.9675 34.825 1.3825 ;
      RECT  35.24 0.9675 37.685 1.3825 ;
      RECT  38.1 0.9675 40.545 1.3825 ;
      RECT  40.96 0.9675 43.405 1.3825 ;
      RECT  43.82 0.9675 46.265 1.3825 ;
      RECT  46.68 0.9675 49.125 1.3825 ;
      RECT  49.54 0.9675 51.985 1.3825 ;
      RECT  52.4 0.9675 54.845 1.3825 ;
      RECT  55.26 0.9675 57.705 1.3825 ;
      RECT  58.12 0.9675 60.565 1.3825 ;
      RECT  60.98 0.9675 63.425 1.3825 ;
      RECT  63.84 0.9675 66.285 1.3825 ;
      RECT  66.7 0.9675 69.145 1.3825 ;
      RECT  69.56 0.9675 72.005 1.3825 ;
      RECT  72.42 0.9675 74.865 1.3825 ;
      RECT  75.28 0.9675 77.725 1.3825 ;
      RECT  78.14 0.9675 80.585 1.3825 ;
      RECT  81.0 0.9675 83.445 1.3825 ;
      RECT  83.86 0.9675 86.305 1.3825 ;
      RECT  86.72 0.9675 89.165 1.3825 ;
      RECT  89.58 0.9675 92.025 1.3825 ;
      RECT  92.44 0.9675 94.885 1.3825 ;
      RECT  95.3 0.9675 97.745 1.3825 ;
      RECT  98.16 0.9675 100.605 1.3825 ;
      RECT  101.02 0.9675 103.465 1.3825 ;
      RECT  103.88 0.9675 106.325 1.3825 ;
      RECT  106.74 0.9675 109.185 1.3825 ;
      RECT  109.6 0.9675 111.83 1.3825 ;
      RECT  0.14 36.5875 14.805 37.0025 ;
      RECT  0.14 37.0025 14.805 62.61 ;
      RECT  14.805 1.3825 15.22 36.5875 ;
      RECT  15.22 36.5875 20.525 37.0025 ;
      RECT  15.22 37.0025 20.525 62.61 ;
      RECT  14.805 37.0025 15.22 39.3175 ;
      RECT  14.805 39.7325 15.22 41.5275 ;
      RECT  14.805 41.9425 15.22 44.2575 ;
      RECT  14.805 44.6725 15.22 62.61 ;
      RECT  88.065 19.8425 88.48 62.61 ;
      RECT  88.48 19.4275 111.83 19.8425 ;
      RECT  88.065 17.1125 88.48 19.4275 ;
      RECT  88.065 14.9025 88.48 16.6975 ;
      RECT  88.065 1.3825 88.48 11.7575 ;
      RECT  88.065 12.1725 88.48 14.4875 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  102.865 19.8425 103.28 61.3675 ;
      RECT  102.865 61.7825 103.28 62.61 ;
      RECT  103.28 19.8425 111.83 61.3675 ;
      RECT  103.28 61.3675 111.83 61.7825 ;
      RECT  103.28 61.7825 111.83 62.61 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 36.5875 ;
      RECT  6.5225 1.3825 14.805 1.4675 ;
      RECT  6.5225 1.4675 14.805 36.5875 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 20.525 1.0525 ;
      RECT  6.5225 1.0525 20.525 1.3825 ;
      RECT  88.48 19.8425 96.7625 61.2825 ;
      RECT  88.48 61.2825 96.7625 61.3675 ;
      RECT  96.7625 19.8425 97.1775 61.2825 ;
      RECT  97.1775 61.2825 102.865 61.3675 ;
      RECT  88.48 61.3675 96.7625 61.6975 ;
      RECT  88.48 61.6975 96.7625 61.7825 ;
      RECT  96.7625 61.6975 97.1775 61.7825 ;
      RECT  97.1775 61.3675 102.865 61.6975 ;
      RECT  97.1775 61.6975 102.865 61.7825 ;
      RECT  20.94 54.66 32.5725 55.075 ;
      RECT  20.94 55.075 32.5725 62.61 ;
      RECT  32.5725 55.075 32.9875 62.61 ;
      RECT  32.9875 55.075 88.065 62.61 ;
      RECT  32.9875 54.66 33.7475 55.075 ;
      RECT  34.1625 54.66 34.9225 55.075 ;
      RECT  35.3375 54.66 36.0975 55.075 ;
      RECT  36.5125 54.66 37.2725 55.075 ;
      RECT  37.6875 54.66 38.4475 55.075 ;
      RECT  38.8625 54.66 39.6225 55.075 ;
      RECT  40.0375 54.66 40.7975 55.075 ;
      RECT  41.2125 54.66 41.9725 55.075 ;
      RECT  42.3875 54.66 43.1475 55.075 ;
      RECT  43.5625 54.66 44.3225 55.075 ;
      RECT  44.7375 54.66 45.4975 55.075 ;
      RECT  45.9125 54.66 46.6725 55.075 ;
      RECT  47.0875 54.66 47.8475 55.075 ;
      RECT  48.2625 54.66 49.0225 55.075 ;
      RECT  49.4375 54.66 50.1975 55.075 ;
      RECT  50.6125 54.66 51.3725 55.075 ;
      RECT  51.7875 54.66 52.5475 55.075 ;
      RECT  52.9625 54.66 53.7225 55.075 ;
      RECT  54.1375 54.66 54.8975 55.075 ;
      RECT  55.3125 54.66 56.0725 55.075 ;
      RECT  56.4875 54.66 57.2475 55.075 ;
      RECT  57.6625 54.66 58.4225 55.075 ;
      RECT  58.8375 54.66 59.5975 55.075 ;
      RECT  60.0125 54.66 60.7725 55.075 ;
      RECT  61.1875 54.66 61.9475 55.075 ;
      RECT  62.3625 54.66 63.1225 55.075 ;
      RECT  63.5375 54.66 64.2975 55.075 ;
      RECT  64.7125 54.66 65.4725 55.075 ;
      RECT  65.8875 54.66 66.6475 55.075 ;
      RECT  67.0625 54.66 67.8225 55.075 ;
      RECT  68.2375 54.66 68.9975 55.075 ;
      RECT  69.4125 54.66 88.065 55.075 ;
      RECT  32.9875 19.8425 82.3325 25.0175 ;
      RECT  32.9875 25.0175 82.3325 25.4325 ;
      RECT  82.7475 25.0175 88.065 25.4325 ;
      RECT  32.9875 25.4325 77.065 45.16 ;
      RECT  32.9875 45.16 77.065 45.575 ;
      RECT  77.065 25.4325 77.48 45.16 ;
      RECT  77.065 45.575 77.48 54.66 ;
      RECT  77.48 25.4325 82.3325 45.16 ;
      RECT  77.48 45.16 82.3325 45.575 ;
      RECT  77.48 45.575 82.3325 54.66 ;
      RECT  20.94 48.205 29.3875 48.555 ;
      RECT  20.94 48.555 29.3875 54.66 ;
      RECT  29.3875 19.8425 32.5725 48.205 ;
      RECT  32.5725 19.8425 32.9875 48.205 ;
      RECT  32.9875 45.575 71.7275 48.205 ;
      RECT  71.7275 48.205 77.065 48.555 ;
      RECT  71.7275 48.555 77.065 54.66 ;
      RECT  20.94 1.3825 43.1225 2.3325 ;
      RECT  43.1225 1.3825 43.5375 2.3325 ;
      RECT  43.5375 1.3825 88.065 2.3325 ;
      RECT  82.3325 19.8425 82.7475 22.0275 ;
      RECT  82.3325 22.4425 82.7475 25.0175 ;
      RECT  20.7575 1.3825 20.94 22.0275 ;
      RECT  20.7575 22.0275 20.94 22.4425 ;
      RECT  20.7575 22.4425 20.94 62.61 ;
      RECT  15.22 22.0275 20.3425 22.4425 ;
      RECT  43.5375 2.3325 54.5625 2.7475 ;
      RECT  54.9775 2.3325 66.0025 2.7475 ;
      RECT  82.3325 34.4025 82.7475 54.66 ;
      RECT  71.7275 45.575 74.4325 45.9475 ;
      RECT  71.7275 45.9475 74.4325 46.3625 ;
      RECT  71.7275 46.3625 74.4325 48.205 ;
      RECT  74.4325 45.575 74.8475 45.9475 ;
      RECT  74.4325 46.3625 74.8475 48.205 ;
      RECT  74.8475 45.575 77.065 45.9475 ;
      RECT  74.8475 45.9475 77.065 46.3625 ;
      RECT  74.8475 46.3625 77.065 48.205 ;
      RECT  20.525 34.4025 20.7575 62.61 ;
      RECT  20.3425 34.4025 20.525 36.5875 ;
      RECT  88.48 1.3825 100.3225 2.3325 ;
      RECT  88.48 2.7475 100.3225 19.4275 ;
      RECT  100.3225 1.3825 100.7375 2.3325 ;
      RECT  100.3225 2.7475 100.7375 19.4275 ;
      RECT  100.7375 1.3825 111.83 2.3325 ;
      RECT  100.7375 2.3325 111.83 2.7475 ;
      RECT  100.7375 2.7475 111.83 19.4275 ;
      RECT  20.525 31.4125 20.7575 33.9875 ;
      RECT  20.3425 31.4125 20.525 33.9875 ;
      RECT  20.94 19.4275 25.61 19.825 ;
      RECT  20.94 19.825 25.61 19.8425 ;
      RECT  25.61 19.4275 26.025 19.825 ;
      RECT  26.025 19.825 88.065 19.8425 ;
      RECT  20.94 19.8425 25.61 20.24 ;
      RECT  20.94 20.24 25.61 48.205 ;
      RECT  25.61 20.24 26.025 48.205 ;
      RECT  26.025 19.8425 29.3875 20.24 ;
      RECT  26.025 20.24 29.3875 48.205 ;
      RECT  20.525 22.4425 20.7575 25.0175 ;
      RECT  20.525 25.4325 20.7575 30.9975 ;
      RECT  20.3425 22.4425 20.525 25.0175 ;
      RECT  20.3425 25.4325 20.525 30.9975 ;
      RECT  29.3875 52.4525 32.5725 54.66 ;
      RECT  32.5725 52.4525 32.9875 54.66 ;
      RECT  32.9875 52.4525 70.0825 54.66 ;
      RECT  70.0825 52.1025 71.7275 52.4525 ;
      RECT  70.0825 52.4525 71.7275 54.66 ;
      RECT  20.94 2.7475 29.3875 16.665 ;
      RECT  20.94 16.665 29.3875 17.015 ;
      RECT  29.3875 17.015 43.1225 19.4275 ;
      RECT  43.1225 17.015 43.5375 19.4275 ;
      RECT  43.5375 17.015 70.5525 19.4275 ;
      RECT  70.5525 2.7475 88.065 16.665 ;
      RECT  70.5525 16.665 88.065 17.015 ;
      RECT  70.5525 17.015 88.065 19.4275 ;
      RECT  88.48 2.3325 88.8825 2.7475 ;
      RECT  89.2975 2.3325 100.3225 2.7475 ;
      RECT  20.525 1.3825 20.6575 2.3325 ;
      RECT  20.525 2.7475 20.6575 22.0275 ;
      RECT  20.6575 1.3825 20.7575 2.3325 ;
      RECT  20.6575 2.3325 20.7575 2.7475 ;
      RECT  20.6575 2.7475 20.7575 22.0275 ;
      RECT  15.22 1.3825 20.2425 2.3325 ;
      RECT  15.22 2.3325 20.2425 2.7475 ;
      RECT  20.2425 1.3825 20.3425 2.3325 ;
      RECT  20.2425 2.7475 20.3425 22.0275 ;
      RECT  20.3425 1.3825 20.525 2.3325 ;
      RECT  20.3425 2.7475 20.525 22.0275 ;
      RECT  66.4175 2.3325 77.4425 2.7475 ;
      RECT  77.8575 2.3325 88.065 2.7475 ;
      RECT  29.3875 2.7475 43.1225 11.23 ;
      RECT  43.1225 2.7475 43.5375 11.23 ;
      RECT  43.5375 2.7475 70.0825 11.23 ;
      RECT  70.0825 2.7475 70.5525 11.23 ;
      RECT  70.0825 11.23 70.5525 11.58 ;
      RECT  70.0825 11.58 70.5525 16.665 ;
      RECT  82.3325 25.4325 82.7475 30.9975 ;
      RECT  82.3325 31.4125 82.7475 33.9875 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 36.5875 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 36.5875 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 36.5875 ;
      RECT  97.1775 19.8425 100.725 60.0025 ;
      RECT  97.1775 60.0025 100.725 60.4175 ;
      RECT  97.1775 60.4175 100.725 61.2825 ;
      RECT  100.725 19.8425 101.14 60.0025 ;
      RECT  100.725 60.4175 101.14 61.2825 ;
      RECT  101.14 19.8425 102.865 60.0025 ;
      RECT  101.14 60.0025 102.865 60.4175 ;
      RECT  101.14 60.4175 102.865 61.2825 ;
      RECT  26.025 19.4275 28.2425 19.4525 ;
      RECT  26.025 19.4525 28.2425 19.825 ;
      RECT  28.2425 19.4525 28.6575 19.825 ;
      RECT  28.6575 19.4275 88.065 19.4525 ;
      RECT  28.6575 19.4525 88.065 19.825 ;
      RECT  20.94 17.015 28.2425 19.0375 ;
      RECT  20.94 19.0375 28.2425 19.4275 ;
      RECT  28.2425 17.015 28.6575 19.0375 ;
      RECT  28.6575 17.015 29.3875 19.0375 ;
      RECT  28.6575 19.0375 29.3875 19.4275 ;
      RECT  20.94 2.3325 31.6825 2.7475 ;
      RECT  32.0975 2.3325 43.1225 2.7475 ;
      RECT  20.94 0.2775 91.7425 0.9675 ;
      RECT  91.7425 0.2775 92.1575 0.9675 ;
      RECT  92.1575 0.2775 111.83 0.9675 ;
      RECT  20.94 0.14 23.1025 0.2775 ;
      RECT  82.7475 19.8425 83.86 23.5225 ;
      RECT  82.7475 23.5225 83.86 23.9375 ;
      RECT  82.7475 23.9375 83.86 25.0175 ;
      RECT  83.86 23.9375 84.275 25.0175 ;
      RECT  84.275 19.8425 88.065 23.5225 ;
      RECT  84.275 23.5225 88.065 23.9375 ;
      RECT  84.275 23.9375 88.065 25.0175 ;
      RECT  82.7475 25.4325 83.86 35.4825 ;
      RECT  82.7475 35.4825 83.86 35.8975 ;
      RECT  82.7475 35.8975 83.86 54.66 ;
      RECT  83.86 35.8975 84.275 54.66 ;
      RECT  84.275 25.4325 88.065 35.4825 ;
      RECT  84.275 35.4825 88.065 35.8975 ;
      RECT  84.275 35.8975 88.065 54.66 ;
      RECT  15.22 22.4425 18.815 23.5225 ;
      RECT  15.22 23.5225 18.815 23.9375 ;
      RECT  15.22 23.9375 18.815 36.5875 ;
      RECT  18.815 22.4425 19.23 23.5225 ;
      RECT  19.23 22.4425 20.3425 23.5225 ;
      RECT  19.23 23.5225 20.3425 23.9375 ;
      RECT  19.23 23.9375 20.3425 36.5875 ;
      RECT  88.48 61.7825 100.725 62.4725 ;
      RECT  88.48 62.4725 100.725 62.61 ;
      RECT  100.725 61.7825 101.14 62.4725 ;
      RECT  101.14 61.7825 102.865 62.4725 ;
      RECT  101.14 62.4725 102.865 62.61 ;
      RECT  83.86 25.4325 84.275 26.5125 ;
      RECT  18.815 23.9375 19.23 26.5125 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  0.14 0.2775 2.285 0.9675 ;
      RECT  2.285 0.2775 2.7 0.9675 ;
      RECT  2.7 0.14 20.525 0.2775 ;
      RECT  2.7 0.2775 20.525 0.9675 ;
      RECT  18.815 26.9275 19.23 29.5025 ;
      RECT  29.3875 48.555 32.5725 50.21 ;
      RECT  29.3875 50.56 32.5725 52.1025 ;
      RECT  32.5725 48.555 32.9875 50.21 ;
      RECT  32.5725 50.56 32.9875 52.1025 ;
      RECT  32.9875 48.555 70.0825 50.21 ;
      RECT  32.9875 50.56 70.0825 52.1025 ;
      RECT  70.0825 48.555 70.1175 50.21 ;
      RECT  70.0825 50.56 70.1175 52.1025 ;
      RECT  70.1175 48.555 71.7275 50.21 ;
      RECT  70.1175 50.21 71.7275 50.56 ;
      RECT  70.1175 50.56 71.7275 52.1025 ;
      RECT  83.86 26.9275 84.275 29.5025 ;
      RECT  57.8375 0.14 68.8625 0.2775 ;
      RECT  46.3975 0.14 57.4225 0.2775 ;
      RECT  83.86 19.8425 84.275 20.5325 ;
      RECT  83.86 20.9475 84.275 23.5225 ;
      RECT  18.815 29.9175 19.23 32.4925 ;
      RECT  83.86 29.9175 84.275 32.4925 ;
      RECT  83.86 32.9075 84.275 35.4825 ;
      RECT  92.1575 0.14 103.1825 0.2775 ;
      RECT  103.5975 0.14 111.83 0.2775 ;
      RECT  69.2775 0.14 80.3025 0.2775 ;
      RECT  80.7175 0.14 91.7425 0.2775 ;
      RECT  15.22 2.7475 18.815 20.5325 ;
      RECT  15.22 20.5325 18.815 20.9475 ;
      RECT  15.22 20.9475 18.815 22.0275 ;
      RECT  18.815 2.7475 19.23 20.5325 ;
      RECT  18.815 20.9475 19.23 22.0275 ;
      RECT  19.23 2.7475 20.2425 20.5325 ;
      RECT  19.23 20.5325 20.2425 20.9475 ;
      RECT  19.23 20.9475 20.2425 22.0275 ;
      RECT  18.815 32.9075 19.23 35.4825 ;
      RECT  18.815 35.8975 19.23 36.5875 ;
      RECT  23.5175 0.14 34.5425 0.2775 ;
      RECT  34.9575 0.14 45.9825 0.2775 ;
      RECT  29.3875 11.58 43.1225 13.28 ;
      RECT  29.3875 13.63 43.1225 16.665 ;
      RECT  43.1225 11.58 43.5375 13.28 ;
      RECT  43.1225 13.63 43.5375 16.665 ;
      RECT  43.5375 11.58 70.0825 13.28 ;
      RECT  43.5375 13.63 70.0825 16.665 ;
   LAYER  metal4 ;
      RECT  74.29 0.14 74.99 20.39 ;
      RECT  74.29 45.01 74.99 62.61 ;
      RECT  17.1 0.14 17.8 2.19 ;
      RECT  17.1 17.71 17.8 20.39 ;
      RECT  17.8 0.14 74.29 2.19 ;
      RECT  24.85 45.08 25.55 62.61 ;
      RECT  0.14 2.19 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 17.71 ;
      RECT  0.4075 2.19 1.1075 9.5675 ;
      RECT  0.14 17.71 0.4075 20.39 ;
      RECT  0.14 20.39 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 45.01 ;
      RECT  0.4075 32.53 1.1075 45.01 ;
      RECT  74.99 45.08 77.54 62.61 ;
      RECT  77.54 45.08 78.24 62.61 ;
      RECT  78.24 45.08 85.485 49.98 ;
      RECT  78.24 49.98 85.485 60.56 ;
      RECT  78.24 60.56 85.485 62.61 ;
      RECT  85.485 45.08 86.185 49.98 ;
      RECT  85.485 60.56 86.185 62.61 ;
      RECT  17.8 2.19 29.18 17.22 ;
      RECT  17.8 17.22 29.18 17.71 ;
      RECT  29.18 2.19 29.88 17.22 ;
      RECT  29.88 2.19 74.29 17.22 ;
      RECT  25.55 45.08 29.18 47.93 ;
      RECT  25.55 47.93 29.18 62.61 ;
      RECT  29.18 47.93 29.88 62.61 ;
      RECT  29.88 47.93 74.29 62.61 ;
      RECT  28.8 20.39 29.18 45.01 ;
      RECT  102.3175 20.39 103.0175 30.22 ;
      RECT  103.0175 20.39 111.83 30.22 ;
      RECT  103.0175 30.22 111.83 45.01 ;
      RECT  103.0175 45.01 111.83 45.08 ;
      RECT  103.0175 45.08 111.83 49.98 ;
      RECT  102.3175 53.1825 103.0175 60.56 ;
      RECT  103.0175 49.98 111.83 53.1825 ;
      RECT  103.0175 53.1825 111.83 60.56 ;
      RECT  0.14 45.01 14.38 45.08 ;
      RECT  0.14 45.08 14.38 45.92 ;
      RECT  0.14 45.92 14.38 62.61 ;
      RECT  14.38 45.92 15.08 62.61 ;
      RECT  1.1075 35.34 14.38 45.01 ;
      RECT  14.38 32.53 15.08 35.34 ;
      RECT  88.205 0.14 88.905 10.51 ;
      RECT  88.905 0.14 111.83 10.51 ;
      RECT  88.905 10.51 111.83 20.39 ;
      RECT  88.205 21.09 88.905 30.22 ;
      RECT  88.905 20.39 102.3175 21.09 ;
      RECT  73.91 17.22 74.29 17.71 ;
      RECT  73.91 17.71 74.29 20.39 ;
      RECT  73.91 45.01 74.29 45.08 ;
      RECT  73.91 45.08 74.29 47.93 ;
      RECT  73.91 20.39 74.29 45.01 ;
      RECT  100.955 30.22 102.3175 45.01 ;
      RECT  100.955 45.01 102.3175 45.08 ;
      RECT  100.955 45.08 102.3175 49.98 ;
      RECT  100.255 53.15 100.955 53.1825 ;
      RECT  100.955 49.98 102.3175 53.15 ;
      RECT  100.955 53.15 102.3175 53.1825 ;
      RECT  88.905 21.09 100.255 30.1875 ;
      RECT  88.905 30.1875 100.255 30.22 ;
      RECT  100.255 21.09 100.955 30.1875 ;
      RECT  100.955 21.09 102.3175 30.1875 ;
      RECT  100.955 30.1875 102.3175 30.22 ;
      RECT  23.96 20.39 24.85 32.53 ;
      RECT  17.8 17.71 23.26 20.3575 ;
      RECT  17.8 20.3575 23.26 20.39 ;
      RECT  23.26 17.71 23.96 20.3575 ;
      RECT  23.96 17.71 29.18 20.3575 ;
      RECT  23.96 45.01 24.85 45.08 ;
      RECT  23.96 32.53 24.85 35.34 ;
      RECT  23.96 35.34 24.85 45.01 ;
      RECT  74.99 20.39 76.98 45.01 ;
      RECT  74.99 45.01 76.98 45.0425 ;
      RECT  74.99 45.0425 76.98 45.08 ;
      RECT  76.98 45.0425 77.54 45.08 ;
      RECT  74.99 10.51 76.98 20.3575 ;
      RECT  74.99 20.3575 76.98 20.39 ;
      RECT  76.98 10.51 77.68 20.3575 ;
      RECT  74.99 0.14 85.345 10.445 ;
      RECT  74.99 10.445 85.345 10.51 ;
      RECT  85.345 0.14 86.045 10.445 ;
      RECT  86.045 0.14 88.205 10.445 ;
      RECT  86.045 10.445 88.205 10.51 ;
      RECT  86.045 20.39 88.205 21.09 ;
      RECT  85.345 21.155 86.045 30.22 ;
      RECT  86.045 21.09 88.205 21.155 ;
      RECT  86.045 21.155 88.205 30.22 ;
      RECT  77.68 10.51 85.345 20.3575 ;
      RECT  86.045 10.51 88.205 20.3575 ;
      RECT  86.045 20.3575 88.205 20.39 ;
      RECT  86.185 60.56 96.76 62.61 ;
      RECT  97.46 60.56 111.83 62.61 ;
      RECT  86.185 53.1825 96.76 60.56 ;
      RECT  97.46 53.1825 102.3175 60.56 ;
      RECT  86.185 45.08 96.76 47.51 ;
      RECT  86.185 47.51 96.76 49.98 ;
      RECT  96.76 45.08 97.46 47.51 ;
      RECT  97.46 45.08 100.255 47.51 ;
      RECT  97.46 47.51 100.255 49.98 ;
      RECT  86.185 49.98 96.76 53.15 ;
      RECT  97.46 49.98 100.255 53.15 ;
      RECT  86.185 53.15 96.76 53.1825 ;
      RECT  97.46 53.15 100.255 53.1825 ;
      RECT  15.08 45.08 17.24 45.92 ;
      RECT  17.94 45.08 24.85 45.92 ;
      RECT  15.08 45.92 17.24 45.985 ;
      RECT  15.08 45.985 17.24 62.61 ;
      RECT  17.24 45.985 17.94 62.61 ;
      RECT  17.94 45.92 24.85 45.985 ;
      RECT  17.94 45.985 24.85 62.61 ;
      RECT  15.08 45.01 17.24 45.08 ;
      RECT  17.94 45.01 23.26 45.08 ;
      RECT  15.08 32.53 17.24 35.275 ;
      RECT  15.08 35.275 17.24 35.34 ;
      RECT  17.24 32.53 17.94 35.275 ;
      RECT  17.94 32.53 23.26 35.275 ;
      RECT  17.94 35.275 23.26 35.34 ;
      RECT  15.08 35.34 17.24 45.01 ;
      RECT  17.94 35.34 23.26 45.01 ;
      RECT  26.11 20.39 28.1 45.01 ;
      RECT  25.55 45.0425 26.11 45.08 ;
      RECT  26.11 45.01 29.18 45.0425 ;
      RECT  26.11 45.0425 29.18 45.08 ;
      RECT  23.96 20.3575 25.41 20.39 ;
      RECT  26.11 20.3575 29.18 20.39 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 17.71 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  1.1075 17.71 2.47 20.39 ;
      RECT  3.17 17.71 17.1 20.39 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 35.34 ;
      RECT  2.47 32.5625 3.17 35.34 ;
      RECT  3.17 32.53 14.38 32.5625 ;
      RECT  3.17 32.5625 14.38 35.34 ;
      RECT  1.1075 20.39 2.47 32.53 ;
      RECT  3.17 20.39 23.26 32.53 ;
      RECT  78.24 30.22 79.13 45.01 ;
      RECT  79.83 30.22 100.255 45.01 ;
      RECT  78.24 45.01 79.13 45.08 ;
      RECT  79.83 45.01 100.255 45.08 ;
      RECT  78.24 20.39 79.13 21.09 ;
      RECT  79.83 20.39 85.345 21.09 ;
      RECT  78.24 21.09 79.13 21.155 ;
      RECT  79.83 21.09 85.345 21.155 ;
      RECT  78.24 21.155 79.13 30.22 ;
      RECT  79.83 21.155 85.345 30.22 ;
      RECT  77.68 20.3575 79.13 20.39 ;
      RECT  79.83 20.3575 85.345 20.39 ;
      RECT  30.34 17.22 72.75 17.71 ;
      RECT  30.34 17.71 72.75 20.39 ;
      RECT  30.34 45.01 72.75 45.08 ;
      RECT  30.34 45.08 72.75 47.93 ;
      RECT  30.34 20.39 72.75 45.01 ;
      RECT  0.14 0.14 5.825 2.19 ;
      RECT  6.525 0.14 17.1 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 17.1 9.5675 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  6.525 9.5675 17.1 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  3.17 15.24 5.825 17.71 ;
      RECT  5.825 15.24 6.525 17.71 ;
      RECT  6.525 9.6 17.1 15.24 ;
      RECT  6.525 15.24 17.1 17.71 ;
   END
END    freepdk45_sram_1w1r_16x32_32
END    LIBRARY
