../macros/freepdk45_sram_1w1r_64x512/freepdk45_sram_1w1r_64x512.lef