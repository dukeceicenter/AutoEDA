VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1rw0r_64x44_22
   CLASS BLOCK ;
   SIZE 157.9 BY 74.4625 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.275 1.105 32.41 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.135 1.105 35.27 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.995 1.105 38.13 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.855 1.105 40.99 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.715 1.105 43.85 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.575 1.105 46.71 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.435 1.105 49.57 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.295 1.105 52.43 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.155 1.105 55.29 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.015 1.105 58.15 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.875 1.105 61.01 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.735 1.105 63.87 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.595 1.105 66.73 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.455 1.105 69.59 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.315 1.105 72.45 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.175 1.105 75.31 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.035 1.105 78.17 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.895 1.105 81.03 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.755 1.105 83.89 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.615 1.105 86.75 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.475 1.105 89.61 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.335 1.105 92.47 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.195 1.105 95.33 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.055 1.105 98.19 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.915 1.105 101.05 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.775 1.105 103.91 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.635 1.105 106.77 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.495 1.105 109.63 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.355 1.105 112.49 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.215 1.105 115.35 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.075 1.105 118.21 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.935 1.105 121.07 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.795 1.105 123.93 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.655 1.105 126.79 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.515 1.105 129.65 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.375 1.105 132.51 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.235 1.105 135.37 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.095 1.105 138.23 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.955 1.105 141.09 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.815 1.105 143.95 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.675 1.105 146.81 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.535 1.105 149.67 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.395 1.105 152.53 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.255 1.105 155.39 1.24 ;
      END
   END din0[43]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.695 1.105 23.83 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.975 49.3675 18.11 49.5025 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.975 52.0975 18.11 52.2325 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.975 54.3075 18.11 54.4425 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.975 57.0375 18.11 57.1725 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.975 59.2475 18.11 59.3825 ;
      END
   END addr0[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 7.3775 0.42 7.5125 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 10.1075 0.42 10.2425 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 7.4625 6.6625 7.5975 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.555 1.105 26.69 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.415 1.105 29.55 1.24 ;
      END
   END wmask0[1]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.5675 16.0725 39.7025 16.2075 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.9775 16.0725 41.1125 16.2075 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.3875 16.0725 42.5225 16.2075 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.7975 16.0725 43.9325 16.2075 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.2075 16.0725 45.3425 16.2075 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.6175 16.0725 46.7525 16.2075 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.0275 16.0725 48.1625 16.2075 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.4375 16.0725 49.5725 16.2075 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.8475 16.0725 50.9825 16.2075 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.2575 16.0725 52.3925 16.2075 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.6675 16.0725 53.8025 16.2075 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.0775 16.0725 55.2125 16.2075 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.4875 16.0725 56.6225 16.2075 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.8975 16.0725 58.0325 16.2075 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.3075 16.0725 59.4425 16.2075 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.7175 16.0725 60.8525 16.2075 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.1275 16.0725 62.2625 16.2075 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.5375 16.0725 63.6725 16.2075 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.9475 16.0725 65.0825 16.2075 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.3575 16.0725 66.4925 16.2075 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.7675 16.0725 67.9025 16.2075 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.1775 16.0725 69.3125 16.2075 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.5875 16.0725 70.7225 16.2075 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.9975 16.0725 72.1325 16.2075 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.4075 16.0725 73.5425 16.2075 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.8175 16.0725 74.9525 16.2075 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.2275 16.0725 76.3625 16.2075 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.6375 16.0725 77.7725 16.2075 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.0475 16.0725 79.1825 16.2075 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.4575 16.0725 80.5925 16.2075 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.8675 16.0725 82.0025 16.2075 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.2775 16.0725 83.4125 16.2075 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.6875 16.0725 84.8225 16.2075 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.0975 16.0725 86.2325 16.2075 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.5075 16.0725 87.6425 16.2075 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.9175 16.0725 89.0525 16.2075 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.3275 16.0725 90.4625 16.2075 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.7375 16.0725 91.8725 16.2075 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.1475 16.0725 93.2825 16.2075 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.5575 16.0725 94.6925 16.2075 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.9675 16.0725 96.1025 16.2075 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.3775 16.0725 97.5125 16.2075 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.7875 16.0725 98.9225 16.2075 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.1975 16.0725 100.3325 16.2075 ;
      END
   END dout0[43]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  37.1875 10.7975 37.3225 10.9325 ;
         LAYER metal3 ;
         RECT  24.0725 41.4375 24.2075 41.5725 ;
         LAYER metal3 ;
         RECT  24.0725 38.7075 24.2075 38.8425 ;
         LAYER metal3 ;
         RECT  77.7525 2.47 77.8875 2.605 ;
         LAYER metal3 ;
         RECT  24.0725 46.8975 24.2075 47.0325 ;
         LAYER metal3 ;
         RECT  89.1925 2.47 89.3275 2.605 ;
         LAYER metal3 ;
         RECT  100.6325 2.47 100.7675 2.605 ;
         LAYER metal3 ;
         RECT  31.9925 2.47 32.1275 2.605 ;
         LAYER metal3 ;
         RECT  43.4325 2.47 43.5675 2.605 ;
         LAYER metal3 ;
         RECT  24.4175 30.5175 24.5525 30.6525 ;
         LAYER metal3 ;
         RECT  101.5725 10.7975 101.7075 10.9325 ;
         LAYER metal4 ;
         RECT  0.6875 16.1175 0.8275 38.52 ;
         LAYER metal3 ;
         RECT  37.3225 25.545 101.7075 25.615 ;
         LAYER metal3 ;
         RECT  112.0725 2.47 112.2075 2.605 ;
         LAYER metal3 ;
         RECT  26.2725 2.47 26.4075 2.605 ;
         LAYER metal3 ;
         RECT  30.245 28.445 30.38 28.58 ;
         LAYER metal3 ;
         RECT  28.195 20.6475 28.33 20.7825 ;
         LAYER metal3 ;
         RECT  134.9525 2.47 135.0875 2.605 ;
         LAYER metal3 ;
         RECT  36.1775 27.7875 36.3125 27.9225 ;
         LAYER metal4 ;
         RECT  29.625 29.15 29.765 73.04 ;
         LAYER metal4 ;
         RECT  103.14 26.24 103.28 74.265 ;
         LAYER metal3 ;
         RECT  37.3225 18.6925 101.0025 18.7625 ;
         LAYER metal3 ;
         RECT  146.3925 2.47 146.5275 2.605 ;
         LAYER metal3 ;
         RECT  66.3125 2.47 66.4475 2.605 ;
         LAYER metal3 ;
         RECT  123.5125 2.47 123.6475 2.605 ;
         LAYER metal4 ;
         RECT  20.41 8.74 20.55 23.7 ;
         LAYER metal3 ;
         RECT  24.0725 44.1675 24.2075 44.3025 ;
         LAYER metal3 ;
         RECT  37.3225 11.765 101.0025 11.835 ;
         LAYER metal4 ;
         RECT  37.255 26.24 37.395 74.265 ;
         LAYER metal3 ;
         RECT  54.8725 2.47 55.0075 2.605 ;
         LAYER metal4 ;
         RECT  0.0 6.27 0.14 11.35 ;
         LAYER metal4 ;
         RECT  36.175 29.15 36.315 72.97 ;
         LAYER metal4 ;
         RECT  17.69 48.26 17.83 60.815 ;
         LAYER metal3 ;
         RECT  24.4175 33.2475 24.5525 33.3825 ;
         LAYER metal3 ;
         RECT  23.4125 2.47 23.5475 2.605 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  37.1875 8.9775 37.3225 9.1125 ;
         LAYER metal4 ;
         RECT  20.55 48.195 20.69 60.75 ;
         LAYER metal3 ;
         RECT  69.1725 0.0 69.3075 0.135 ;
         LAYER metal3 ;
         RECT  22.265 48.2625 22.4 48.3975 ;
         LAYER metal4 ;
         RECT  2.75 16.15 2.89 38.5525 ;
         LAYER metal3 ;
         RECT  34.8525 0.0 34.9875 0.135 ;
         LAYER metal3 ;
         RECT  22.89 31.8825 23.025 32.0175 ;
         LAYER metal3 ;
         RECT  22.265 37.3425 22.4 37.4775 ;
         LAYER metal3 ;
         RECT  28.195 18.1775 28.33 18.3125 ;
         LAYER metal3 ;
         RECT  22.89 34.6125 23.025 34.7475 ;
         LAYER metal3 ;
         RECT  37.3225 20.585 101.0375 20.655 ;
         LAYER metal3 ;
         RECT  22.89 29.1525 23.025 29.2875 ;
         LAYER metal3 ;
         RECT  26.2725 0.0 26.4075 0.135 ;
         LAYER metal4 ;
         RECT  37.715 26.24 37.855 74.265 ;
         LAYER metal4 ;
         RECT  6.385 6.27 6.525 26.17 ;
         LAYER metal3 ;
         RECT  37.3225 22.925 101.74 22.995 ;
         LAYER metal3 ;
         RECT  103.4925 0.0 103.6275 0.135 ;
         LAYER metal3 ;
         RECT  92.0525 0.0 92.1875 0.135 ;
         LAYER metal3 ;
         RECT  22.265 45.5325 22.4 45.6675 ;
         LAYER metal4 ;
         RECT  28.035 29.1175 28.175 73.04 ;
         LAYER metal3 ;
         RECT  126.3725 0.0 126.5075 0.135 ;
         LAYER metal4 ;
         RECT  4.845 6.205 4.985 11.415 ;
         LAYER metal3 ;
         RECT  22.265 40.0725 22.4 40.2075 ;
         LAYER metal3 ;
         RECT  29.1325 0.0 29.2675 0.135 ;
         LAYER metal3 ;
         RECT  149.2525 0.0 149.3875 0.135 ;
         LAYER metal4 ;
         RECT  102.68 26.24 102.82 74.265 ;
         LAYER metal3 ;
         RECT  46.2925 0.0 46.4275 0.135 ;
         LAYER metal3 ;
         RECT  37.3225 13.815 101.0025 13.885 ;
         LAYER metal3 ;
         RECT  114.9325 0.0 115.0675 0.135 ;
         LAYER metal3 ;
         RECT  137.8125 0.0 137.9475 0.135 ;
         LAYER metal4 ;
         RECT  30.185 29.1175 30.325 73.0025 ;
         LAYER metal3 ;
         RECT  28.195 23.1175 28.33 23.2525 ;
         LAYER metal3 ;
         RECT  101.5725 8.9775 101.7075 9.1125 ;
         LAYER metal3 ;
         RECT  80.6125 0.0 80.7475 0.135 ;
         LAYER metal3 ;
         RECT  57.7325 0.0 57.8675 0.135 ;
         LAYER metal3 ;
         RECT  22.265 42.8025 22.4 42.9375 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 157.76 74.3225 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 157.76 74.3225 ;
   LAYER  metal3 ;
      RECT  32.135 0.14 32.55 0.965 ;
      RECT  32.55 0.965 34.995 1.38 ;
      RECT  35.41 0.965 37.855 1.38 ;
      RECT  38.27 0.965 40.715 1.38 ;
      RECT  41.13 0.965 43.575 1.38 ;
      RECT  43.99 0.965 46.435 1.38 ;
      RECT  46.85 0.965 49.295 1.38 ;
      RECT  49.71 0.965 52.155 1.38 ;
      RECT  52.57 0.965 55.015 1.38 ;
      RECT  55.43 0.965 57.875 1.38 ;
      RECT  58.29 0.965 60.735 1.38 ;
      RECT  61.15 0.965 63.595 1.38 ;
      RECT  64.01 0.965 66.455 1.38 ;
      RECT  66.87 0.965 69.315 1.38 ;
      RECT  69.73 0.965 72.175 1.38 ;
      RECT  72.59 0.965 75.035 1.38 ;
      RECT  75.45 0.965 77.895 1.38 ;
      RECT  78.31 0.965 80.755 1.38 ;
      RECT  81.17 0.965 83.615 1.38 ;
      RECT  84.03 0.965 86.475 1.38 ;
      RECT  86.89 0.965 89.335 1.38 ;
      RECT  89.75 0.965 92.195 1.38 ;
      RECT  92.61 0.965 95.055 1.38 ;
      RECT  95.47 0.965 97.915 1.38 ;
      RECT  98.33 0.965 100.775 1.38 ;
      RECT  101.19 0.965 103.635 1.38 ;
      RECT  104.05 0.965 106.495 1.38 ;
      RECT  106.91 0.965 109.355 1.38 ;
      RECT  109.77 0.965 112.215 1.38 ;
      RECT  112.63 0.965 115.075 1.38 ;
      RECT  115.49 0.965 117.935 1.38 ;
      RECT  118.35 0.965 120.795 1.38 ;
      RECT  121.21 0.965 123.655 1.38 ;
      RECT  124.07 0.965 126.515 1.38 ;
      RECT  126.93 0.965 129.375 1.38 ;
      RECT  129.79 0.965 132.235 1.38 ;
      RECT  132.65 0.965 135.095 1.38 ;
      RECT  135.51 0.965 137.955 1.38 ;
      RECT  138.37 0.965 140.815 1.38 ;
      RECT  141.23 0.965 143.675 1.38 ;
      RECT  144.09 0.965 146.535 1.38 ;
      RECT  146.95 0.965 149.395 1.38 ;
      RECT  149.81 0.965 152.255 1.38 ;
      RECT  152.67 0.965 155.115 1.38 ;
      RECT  155.53 0.965 157.76 1.38 ;
      RECT  0.14 0.965 23.555 1.38 ;
      RECT  0.14 49.2275 17.835 49.6425 ;
      RECT  0.14 49.6425 17.835 74.3225 ;
      RECT  17.835 1.38 18.25 49.2275 ;
      RECT  18.25 49.2275 32.135 49.6425 ;
      RECT  18.25 49.6425 32.135 74.3225 ;
      RECT  17.835 49.6425 18.25 51.9575 ;
      RECT  17.835 52.3725 18.25 54.1675 ;
      RECT  17.835 54.5825 18.25 56.8975 ;
      RECT  17.835 57.3125 18.25 59.1075 ;
      RECT  17.835 59.5225 18.25 74.3225 ;
      RECT  0.14 1.38 0.145 7.2375 ;
      RECT  0.14 7.2375 0.145 7.6525 ;
      RECT  0.14 7.6525 0.145 49.2275 ;
      RECT  0.145 1.38 0.56 7.2375 ;
      RECT  0.56 1.38 17.835 7.2375 ;
      RECT  0.145 7.6525 0.56 9.9675 ;
      RECT  0.145 10.3825 0.56 49.2275 ;
      RECT  0.56 7.2375 6.3875 7.3225 ;
      RECT  0.56 7.3225 6.3875 7.6525 ;
      RECT  6.3875 7.2375 6.8025 7.3225 ;
      RECT  6.8025 7.2375 17.835 7.3225 ;
      RECT  6.8025 7.3225 17.835 7.6525 ;
      RECT  0.56 7.6525 6.3875 7.7375 ;
      RECT  0.56 7.7375 6.3875 49.2275 ;
      RECT  6.3875 7.7375 6.8025 49.2275 ;
      RECT  6.8025 7.6525 17.835 7.7375 ;
      RECT  6.8025 7.7375 17.835 49.2275 ;
      RECT  23.97 0.965 26.415 1.38 ;
      RECT  26.83 0.965 29.275 1.38 ;
      RECT  29.69 0.965 32.135 1.38 ;
      RECT  32.55 15.9325 39.4275 16.3475 ;
      RECT  39.8425 15.9325 40.8375 16.3475 ;
      RECT  41.2525 15.9325 42.2475 16.3475 ;
      RECT  42.6625 15.9325 43.6575 16.3475 ;
      RECT  44.0725 15.9325 45.0675 16.3475 ;
      RECT  45.4825 15.9325 46.4775 16.3475 ;
      RECT  46.8925 15.9325 47.8875 16.3475 ;
      RECT  48.3025 15.9325 49.2975 16.3475 ;
      RECT  49.7125 15.9325 50.7075 16.3475 ;
      RECT  51.1225 15.9325 52.1175 16.3475 ;
      RECT  52.5325 15.9325 53.5275 16.3475 ;
      RECT  53.9425 15.9325 54.9375 16.3475 ;
      RECT  55.3525 15.9325 56.3475 16.3475 ;
      RECT  56.7625 15.9325 57.7575 16.3475 ;
      RECT  58.1725 15.9325 59.1675 16.3475 ;
      RECT  59.5825 15.9325 60.5775 16.3475 ;
      RECT  60.9925 15.9325 61.9875 16.3475 ;
      RECT  62.4025 15.9325 63.3975 16.3475 ;
      RECT  63.8125 15.9325 64.8075 16.3475 ;
      RECT  65.2225 15.9325 66.2175 16.3475 ;
      RECT  66.6325 15.9325 67.6275 16.3475 ;
      RECT  68.0425 15.9325 69.0375 16.3475 ;
      RECT  69.4525 15.9325 70.4475 16.3475 ;
      RECT  70.8625 15.9325 71.8575 16.3475 ;
      RECT  72.2725 15.9325 73.2675 16.3475 ;
      RECT  73.6825 15.9325 74.6775 16.3475 ;
      RECT  75.0925 15.9325 76.0875 16.3475 ;
      RECT  76.5025 15.9325 77.4975 16.3475 ;
      RECT  77.9125 15.9325 78.9075 16.3475 ;
      RECT  79.3225 15.9325 80.3175 16.3475 ;
      RECT  80.7325 15.9325 81.7275 16.3475 ;
      RECT  82.1425 15.9325 83.1375 16.3475 ;
      RECT  83.5525 15.9325 84.5475 16.3475 ;
      RECT  84.9625 15.9325 85.9575 16.3475 ;
      RECT  86.3725 15.9325 87.3675 16.3475 ;
      RECT  87.7825 15.9325 88.7775 16.3475 ;
      RECT  89.1925 15.9325 90.1875 16.3475 ;
      RECT  90.6025 15.9325 91.5975 16.3475 ;
      RECT  92.0125 15.9325 93.0075 16.3475 ;
      RECT  93.4225 15.9325 94.4175 16.3475 ;
      RECT  94.8325 15.9325 95.8275 16.3475 ;
      RECT  96.2425 15.9325 97.2375 16.3475 ;
      RECT  97.6525 15.9325 98.6475 16.3475 ;
      RECT  99.0625 15.9325 100.0575 16.3475 ;
      RECT  100.4725 15.9325 157.76 16.3475 ;
      RECT  32.55 1.38 37.0475 10.6575 ;
      RECT  32.55 10.6575 37.0475 11.0725 ;
      RECT  32.55 11.0725 37.0475 15.9325 ;
      RECT  37.4625 1.38 39.4275 10.6575 ;
      RECT  37.4625 10.6575 39.4275 11.0725 ;
      RECT  18.25 41.2975 23.9325 41.7125 ;
      RECT  24.3475 41.2975 32.135 41.7125 ;
      RECT  24.3475 41.7125 32.135 49.2275 ;
      RECT  23.9325 38.9825 24.3475 41.2975 ;
      RECT  39.8425 1.38 77.6125 2.33 ;
      RECT  77.6125 1.38 78.0275 2.33 ;
      RECT  78.0275 1.38 157.76 2.33 ;
      RECT  23.9325 47.1725 24.3475 49.2275 ;
      RECT  78.0275 2.33 89.0525 2.745 ;
      RECT  89.4675 2.33 100.4925 2.745 ;
      RECT  32.135 1.38 32.2675 2.33 ;
      RECT  32.135 2.745 32.2675 74.3225 ;
      RECT  32.2675 1.38 32.55 2.33 ;
      RECT  32.2675 2.33 32.55 2.745 ;
      RECT  32.2675 2.745 32.55 74.3225 ;
      RECT  24.3475 1.38 31.8525 2.33 ;
      RECT  31.8525 1.38 32.135 2.33 ;
      RECT  31.8525 2.745 32.135 41.2975 ;
      RECT  39.8425 2.33 43.2925 2.745 ;
      RECT  23.9325 1.38 24.2775 30.3775 ;
      RECT  23.9325 30.3775 24.2775 30.7925 ;
      RECT  23.9325 30.7925 24.2775 38.5675 ;
      RECT  24.2775 1.38 24.3475 30.3775 ;
      RECT  24.3475 2.745 24.6925 30.3775 ;
      RECT  24.6925 30.3775 31.8525 30.7925 ;
      RECT  24.6925 30.7925 31.8525 41.2975 ;
      RECT  78.0275 2.745 101.4325 10.6575 ;
      RECT  78.0275 10.6575 101.4325 11.0725 ;
      RECT  101.4325 11.0725 101.8475 15.9325 ;
      RECT  101.8475 2.745 157.76 10.6575 ;
      RECT  101.8475 10.6575 157.76 11.0725 ;
      RECT  101.8475 11.0725 157.76 15.9325 ;
      RECT  32.55 16.3475 37.1825 25.405 ;
      RECT  32.55 25.405 37.1825 25.755 ;
      RECT  37.1825 25.755 39.4275 74.3225 ;
      RECT  39.4275 25.755 39.8425 74.3225 ;
      RECT  39.8425 25.755 101.8475 74.3225 ;
      RECT  101.8475 25.405 157.76 25.755 ;
      RECT  101.8475 25.755 157.76 74.3225 ;
      RECT  100.9075 2.33 111.9325 2.745 ;
      RECT  24.3475 2.33 26.1325 2.745 ;
      RECT  26.5475 2.33 31.8525 2.745 ;
      RECT  24.6925 28.305 30.105 28.72 ;
      RECT  24.6925 28.72 30.105 30.3775 ;
      RECT  30.105 2.745 30.52 28.305 ;
      RECT  30.105 28.72 30.52 30.3775 ;
      RECT  30.52 2.745 31.8525 28.305 ;
      RECT  30.52 28.305 31.8525 28.72 ;
      RECT  30.52 28.72 31.8525 30.3775 ;
      RECT  24.6925 2.745 28.055 20.5075 ;
      RECT  24.6925 20.5075 28.055 20.9225 ;
      RECT  24.6925 20.9225 28.055 28.305 ;
      RECT  28.47 2.745 30.105 20.5075 ;
      RECT  28.47 20.5075 30.105 20.9225 ;
      RECT  28.47 20.9225 30.105 28.305 ;
      RECT  32.55 25.755 36.0375 27.6475 ;
      RECT  32.55 27.6475 36.0375 28.0625 ;
      RECT  32.55 28.0625 36.0375 74.3225 ;
      RECT  36.0375 25.755 36.4525 27.6475 ;
      RECT  36.0375 28.0625 36.4525 74.3225 ;
      RECT  36.4525 25.755 37.1825 27.6475 ;
      RECT  36.4525 27.6475 37.1825 28.0625 ;
      RECT  36.4525 28.0625 37.1825 74.3225 ;
      RECT  37.1825 16.3475 39.4275 18.5525 ;
      RECT  39.4275 16.3475 39.8425 18.5525 ;
      RECT  39.8425 16.3475 101.1425 18.5525 ;
      RECT  101.1425 16.3475 101.8475 18.5525 ;
      RECT  101.1425 18.5525 101.8475 18.9025 ;
      RECT  135.2275 2.33 146.2525 2.745 ;
      RECT  146.6675 2.33 157.76 2.745 ;
      RECT  66.5875 2.33 77.6125 2.745 ;
      RECT  112.3475 2.33 123.3725 2.745 ;
      RECT  123.7875 2.33 134.8125 2.745 ;
      RECT  23.9325 41.7125 24.3475 44.0275 ;
      RECT  23.9325 44.4425 24.3475 46.7575 ;
      RECT  39.4275 1.38 39.8425 11.625 ;
      RECT  37.0475 11.0725 37.1825 11.625 ;
      RECT  37.0475 11.625 37.1825 11.975 ;
      RECT  37.0475 11.975 37.1825 15.9325 ;
      RECT  37.1825 11.0725 37.4625 11.625 ;
      RECT  37.4625 11.0725 39.4275 11.625 ;
      RECT  39.8425 2.745 77.6125 11.625 ;
      RECT  77.6125 2.745 78.0275 11.625 ;
      RECT  78.0275 11.0725 101.1425 11.625 ;
      RECT  101.1425 11.0725 101.4325 11.625 ;
      RECT  101.1425 11.625 101.4325 11.975 ;
      RECT  101.1425 11.975 101.4325 15.9325 ;
      RECT  43.7075 2.33 54.7325 2.745 ;
      RECT  55.1475 2.33 66.1725 2.745 ;
      RECT  24.2775 30.7925 24.3475 33.1075 ;
      RECT  24.2775 33.5225 24.3475 38.5675 ;
      RECT  24.3475 30.7925 24.6925 33.1075 ;
      RECT  24.3475 33.5225 24.6925 41.2975 ;
      RECT  18.25 1.38 23.2725 2.33 ;
      RECT  18.25 2.33 23.2725 2.745 ;
      RECT  23.2725 1.38 23.6875 2.33 ;
      RECT  23.2725 2.745 23.6875 41.2975 ;
      RECT  23.6875 1.38 23.9325 2.33 ;
      RECT  23.6875 2.33 23.9325 2.745 ;
      RECT  23.6875 2.745 23.9325 41.2975 ;
      RECT  37.0475 1.38 37.4625 8.8375 ;
      RECT  37.0475 9.2525 37.4625 10.6575 ;
      RECT  32.55 0.275 69.0325 0.965 ;
      RECT  69.0325 0.275 69.4475 0.965 ;
      RECT  69.4475 0.275 157.76 0.965 ;
      RECT  18.25 41.7125 22.125 48.1225 ;
      RECT  18.25 48.1225 22.125 48.5375 ;
      RECT  18.25 48.5375 22.125 49.2275 ;
      RECT  22.125 48.5375 22.54 49.2275 ;
      RECT  22.54 41.7125 23.9325 48.1225 ;
      RECT  22.54 48.1225 23.9325 48.5375 ;
      RECT  22.54 48.5375 23.9325 49.2275 ;
      RECT  32.55 0.14 34.7125 0.275 ;
      RECT  18.25 2.745 22.75 31.7425 ;
      RECT  18.25 31.7425 22.75 32.1575 ;
      RECT  23.165 2.745 23.2725 31.7425 ;
      RECT  23.165 31.7425 23.2725 32.1575 ;
      RECT  23.165 32.1575 23.2725 41.2975 ;
      RECT  18.25 32.1575 22.125 37.2025 ;
      RECT  18.25 37.2025 22.125 37.6175 ;
      RECT  18.25 37.6175 22.125 41.2975 ;
      RECT  22.125 32.1575 22.54 37.2025 ;
      RECT  22.54 32.1575 22.75 37.2025 ;
      RECT  22.54 37.2025 22.75 37.6175 ;
      RECT  22.54 37.6175 22.75 41.2975 ;
      RECT  28.055 2.745 28.47 18.0375 ;
      RECT  28.055 18.4525 28.47 20.5075 ;
      RECT  22.75 32.1575 23.165 34.4725 ;
      RECT  22.75 34.8875 23.165 41.2975 ;
      RECT  37.1825 18.9025 39.4275 20.445 ;
      RECT  39.4275 18.9025 39.8425 20.445 ;
      RECT  39.8425 18.9025 101.1425 20.445 ;
      RECT  101.1425 18.9025 101.1775 20.445 ;
      RECT  101.1775 18.9025 101.8475 20.445 ;
      RECT  101.1775 20.445 101.8475 20.795 ;
      RECT  22.75 2.745 23.165 29.0125 ;
      RECT  22.75 29.4275 23.165 31.7425 ;
      RECT  0.14 0.14 26.1325 0.275 ;
      RECT  0.14 0.275 26.1325 0.965 ;
      RECT  26.1325 0.275 26.5475 0.965 ;
      RECT  26.5475 0.275 32.135 0.965 ;
      RECT  101.8475 16.3475 101.88 22.785 ;
      RECT  101.8475 23.135 101.88 25.405 ;
      RECT  101.88 16.3475 157.76 22.785 ;
      RECT  101.88 22.785 157.76 23.135 ;
      RECT  101.88 23.135 157.76 25.405 ;
      RECT  37.1825 20.795 39.4275 22.785 ;
      RECT  37.1825 23.135 39.4275 25.405 ;
      RECT  39.4275 20.795 39.8425 22.785 ;
      RECT  39.4275 23.135 39.8425 25.405 ;
      RECT  39.8425 20.795 101.1425 22.785 ;
      RECT  39.8425 23.135 101.1425 25.405 ;
      RECT  101.1425 20.795 101.1775 22.785 ;
      RECT  101.1425 23.135 101.1775 25.405 ;
      RECT  101.1775 20.795 101.8475 22.785 ;
      RECT  101.1775 23.135 101.8475 25.405 ;
      RECT  92.3275 0.14 103.3525 0.275 ;
      RECT  22.125 45.8075 22.54 48.1225 ;
      RECT  22.125 37.6175 22.54 39.9325 ;
      RECT  22.125 40.3475 22.54 41.2975 ;
      RECT  26.5475 0.14 28.9925 0.275 ;
      RECT  29.4075 0.14 32.135 0.275 ;
      RECT  149.5275 0.14 157.76 0.275 ;
      RECT  35.1275 0.14 46.1525 0.275 ;
      RECT  39.4275 11.975 39.8425 13.675 ;
      RECT  39.4275 14.025 39.8425 15.9325 ;
      RECT  37.1825 11.975 37.4625 13.675 ;
      RECT  37.1825 14.025 37.4625 15.9325 ;
      RECT  37.4625 11.975 39.4275 13.675 ;
      RECT  37.4625 14.025 39.4275 15.9325 ;
      RECT  39.8425 11.975 77.6125 13.675 ;
      RECT  39.8425 14.025 77.6125 15.9325 ;
      RECT  77.6125 11.975 78.0275 13.675 ;
      RECT  77.6125 14.025 78.0275 15.9325 ;
      RECT  78.0275 11.975 101.1425 13.675 ;
      RECT  78.0275 14.025 101.1425 15.9325 ;
      RECT  103.7675 0.14 114.7925 0.275 ;
      RECT  115.2075 0.14 126.2325 0.275 ;
      RECT  126.6475 0.14 137.6725 0.275 ;
      RECT  138.0875 0.14 149.1125 0.275 ;
      RECT  28.055 20.9225 28.47 22.9775 ;
      RECT  28.055 23.3925 28.47 28.305 ;
      RECT  101.4325 2.745 101.8475 8.8375 ;
      RECT  101.4325 9.2525 101.8475 10.6575 ;
      RECT  69.4475 0.14 80.4725 0.275 ;
      RECT  80.8875 0.14 91.9125 0.275 ;
      RECT  46.5675 0.14 57.5925 0.275 ;
      RECT  58.0075 0.14 69.0325 0.275 ;
      RECT  22.125 41.7125 22.54 42.6625 ;
      RECT  22.125 43.0775 22.54 45.3925 ;
   LAYER  metal4 ;
      RECT  0.14 15.8375 0.4075 38.8 ;
      RECT  0.14 38.8 0.4075 74.3225 ;
      RECT  0.4075 38.8 1.1075 74.3225 ;
      RECT  1.1075 73.32 29.345 74.3225 ;
      RECT  29.345 73.32 30.045 74.3225 ;
      RECT  30.045 15.8375 102.86 25.96 ;
      RECT  102.86 15.8375 103.56 25.96 ;
      RECT  103.56 15.8375 157.76 25.96 ;
      RECT  103.56 25.96 157.76 28.87 ;
      RECT  103.56 28.87 157.76 38.8 ;
      RECT  103.56 38.8 157.76 73.32 ;
      RECT  103.56 73.32 157.76 74.3225 ;
      RECT  20.13 0.14 20.83 8.46 ;
      RECT  20.83 0.14 157.76 8.46 ;
      RECT  20.83 8.46 157.76 15.8375 ;
      RECT  20.13 23.98 20.83 28.87 ;
      RECT  20.83 15.8375 29.345 23.98 ;
      RECT  30.045 73.32 36.975 74.3225 ;
      RECT  0.14 0.14 0.4075 5.99 ;
      RECT  0.14 11.63 0.4075 15.8375 ;
      RECT  0.4075 0.14 0.42 5.99 ;
      RECT  0.4075 11.63 0.42 15.8375 ;
      RECT  0.42 0.14 1.1075 5.99 ;
      RECT  0.42 5.99 1.1075 11.63 ;
      RECT  0.42 11.63 1.1075 15.8375 ;
      RECT  36.595 28.87 36.975 38.8 ;
      RECT  35.895 73.25 36.595 73.32 ;
      RECT  36.595 38.8 36.975 73.25 ;
      RECT  36.595 73.25 36.975 73.32 ;
      RECT  1.1075 47.98 17.41 61.095 ;
      RECT  1.1075 61.095 17.41 73.32 ;
      RECT  17.41 38.8 18.11 47.98 ;
      RECT  17.41 61.095 18.11 73.32 ;
      RECT  18.11 38.8 20.27 47.915 ;
      RECT  18.11 47.915 20.27 47.98 ;
      RECT  20.27 38.8 20.97 47.915 ;
      RECT  18.11 47.98 20.27 61.03 ;
      RECT  18.11 61.03 20.27 61.095 ;
      RECT  20.27 61.03 20.97 61.095 ;
      RECT  1.1075 28.87 2.47 38.8 ;
      RECT  1.1075 15.8375 2.47 15.87 ;
      RECT  1.1075 15.87 2.47 23.98 ;
      RECT  2.47 15.8375 3.17 15.87 ;
      RECT  1.1075 23.98 2.47 28.87 ;
      RECT  1.1075 38.8 2.47 38.8325 ;
      RECT  1.1075 38.8325 2.47 47.98 ;
      RECT  2.47 38.8325 3.17 47.98 ;
      RECT  3.17 38.8 17.41 38.8325 ;
      RECT  3.17 38.8325 17.41 47.98 ;
      RECT  6.105 0.14 6.805 5.99 ;
      RECT  6.805 0.14 20.13 5.99 ;
      RECT  6.805 5.99 20.13 8.46 ;
      RECT  6.805 8.46 20.13 15.8375 ;
      RECT  3.17 15.8375 6.105 15.87 ;
      RECT  6.805 15.8375 20.13 15.87 ;
      RECT  3.17 15.87 6.105 23.98 ;
      RECT  6.805 15.87 20.13 23.98 ;
      RECT  3.17 23.98 6.105 26.45 ;
      RECT  3.17 26.45 6.105 28.87 ;
      RECT  6.105 26.45 6.805 28.87 ;
      RECT  6.805 23.98 20.13 26.45 ;
      RECT  6.805 26.45 20.13 28.87 ;
      RECT  20.83 23.98 27.755 28.8375 ;
      RECT  20.83 28.8375 27.755 28.87 ;
      RECT  27.755 23.98 28.455 28.8375 ;
      RECT  28.455 23.98 29.345 28.8375 ;
      RECT  28.455 28.8375 29.345 28.87 ;
      RECT  18.11 61.095 27.755 73.32 ;
      RECT  28.455 61.095 29.345 73.32 ;
      RECT  20.97 38.8 27.755 47.915 ;
      RECT  28.455 38.8 29.345 47.915 ;
      RECT  20.97 47.915 27.755 47.98 ;
      RECT  28.455 47.915 29.345 47.98 ;
      RECT  20.97 47.98 27.755 61.03 ;
      RECT  28.455 47.98 29.345 61.03 ;
      RECT  20.97 61.03 27.755 61.095 ;
      RECT  28.455 61.03 29.345 61.095 ;
      RECT  3.17 28.87 27.755 38.8 ;
      RECT  28.455 28.87 29.345 38.8 ;
      RECT  1.1075 0.14 4.565 5.925 ;
      RECT  1.1075 5.925 4.565 5.99 ;
      RECT  4.565 0.14 5.265 5.925 ;
      RECT  5.265 0.14 6.105 5.925 ;
      RECT  5.265 5.925 6.105 5.99 ;
      RECT  1.1075 5.99 4.565 8.46 ;
      RECT  5.265 5.99 6.105 8.46 ;
      RECT  1.1075 8.46 4.565 11.695 ;
      RECT  1.1075 11.695 4.565 15.8375 ;
      RECT  4.565 11.695 5.265 15.8375 ;
      RECT  5.265 8.46 6.105 11.695 ;
      RECT  5.265 11.695 6.105 15.8375 ;
      RECT  38.135 25.96 102.4 28.87 ;
      RECT  38.135 28.87 102.4 38.8 ;
      RECT  38.135 38.8 102.4 73.32 ;
      RECT  38.135 73.32 102.4 74.3225 ;
      RECT  29.345 15.8375 29.905 28.8375 ;
      RECT  29.345 28.8375 29.905 28.87 ;
      RECT  29.905 15.8375 30.045 28.8375 ;
      RECT  30.045 25.96 30.605 28.8375 ;
      RECT  30.605 25.96 36.975 28.8375 ;
      RECT  30.605 28.8375 36.975 28.87 ;
      RECT  30.605 28.87 35.895 38.8 ;
      RECT  30.605 38.8 35.895 73.25 ;
      RECT  30.045 73.2825 30.605 73.32 ;
      RECT  30.605 73.25 35.895 73.2825 ;
      RECT  30.605 73.2825 35.895 73.32 ;
   END
END    freepdk45_sram_1rw0r_64x44_22
END    LIBRARY
