../macros/freepdk45_sram_1w1r_128x52_13/freepdk45_sram_1w1r_128x52_13.lef