VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_31x128
   CLASS BLOCK ;
   SIZE 414.54 BY 103.18 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.425 4.2375 45.56 4.3725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.285 4.2375 48.42 4.3725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.145 4.2375 51.28 4.3725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.005 4.2375 54.14 4.3725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.865 4.2375 57.0 4.3725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.725 4.2375 59.86 4.3725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.585 4.2375 62.72 4.3725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.445 4.2375 65.58 4.3725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.305 4.2375 68.44 4.3725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.165 4.2375 71.3 4.3725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.025 4.2375 74.16 4.3725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.885 4.2375 77.02 4.3725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.745 4.2375 79.88 4.3725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.605 4.2375 82.74 4.3725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.465 4.2375 85.6 4.3725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.325 4.2375 88.46 4.3725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.185 4.2375 91.32 4.3725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.045 4.2375 94.18 4.3725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.905 4.2375 97.04 4.3725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.765 4.2375 99.9 4.3725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.625 4.2375 102.76 4.3725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.485 4.2375 105.62 4.3725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.345 4.2375 108.48 4.3725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.205 4.2375 111.34 4.3725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.065 4.2375 114.2 4.3725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.925 4.2375 117.06 4.3725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.785 4.2375 119.92 4.3725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.645 4.2375 122.78 4.3725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.505 4.2375 125.64 4.3725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.365 4.2375 128.5 4.3725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.225 4.2375 131.36 4.3725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.085 4.2375 134.22 4.3725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.945 4.2375 137.08 4.3725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.805 4.2375 139.94 4.3725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.665 4.2375 142.8 4.3725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.525 4.2375 145.66 4.3725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.385 4.2375 148.52 4.3725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.245 4.2375 151.38 4.3725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.105 4.2375 154.24 4.3725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.965 4.2375 157.1 4.3725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.825 4.2375 159.96 4.3725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.685 4.2375 162.82 4.3725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.545 4.2375 165.68 4.3725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.405 4.2375 168.54 4.3725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.265 4.2375 171.4 4.3725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.125 4.2375 174.26 4.3725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.985 4.2375 177.12 4.3725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.845 4.2375 179.98 4.3725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.705 4.2375 182.84 4.3725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.565 4.2375 185.7 4.3725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.425 4.2375 188.56 4.3725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.285 4.2375 191.42 4.3725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.145 4.2375 194.28 4.3725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.005 4.2375 197.14 4.3725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.865 4.2375 200.0 4.3725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.725 4.2375 202.86 4.3725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.585 4.2375 205.72 4.3725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.445 4.2375 208.58 4.3725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.305 4.2375 211.44 4.3725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.165 4.2375 214.3 4.3725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.025 4.2375 217.16 4.3725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.885 4.2375 220.02 4.3725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.745 4.2375 222.88 4.3725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.605 4.2375 225.74 4.3725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.465 4.2375 228.6 4.3725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.325 4.2375 231.46 4.3725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.185 4.2375 234.32 4.3725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.045 4.2375 237.18 4.3725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.905 4.2375 240.04 4.3725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.765 4.2375 242.9 4.3725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.625 4.2375 245.76 4.3725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.485 4.2375 248.62 4.3725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.345 4.2375 251.48 4.3725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.205 4.2375 254.34 4.3725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.065 4.2375 257.2 4.3725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.925 4.2375 260.06 4.3725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.785 4.2375 262.92 4.3725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.645 4.2375 265.78 4.3725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.505 4.2375 268.64 4.3725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.365 4.2375 271.5 4.3725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.225 4.2375 274.36 4.3725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.085 4.2375 277.22 4.3725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.945 4.2375 280.08 4.3725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  282.805 4.2375 282.94 4.3725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.665 4.2375 285.8 4.3725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.525 4.2375 288.66 4.3725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.385 4.2375 291.52 4.3725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.245 4.2375 294.38 4.3725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.105 4.2375 297.24 4.3725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.965 4.2375 300.1 4.3725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  302.825 4.2375 302.96 4.3725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.685 4.2375 305.82 4.3725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.545 4.2375 308.68 4.3725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.405 4.2375 311.54 4.3725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.265 4.2375 314.4 4.3725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.125 4.2375 317.26 4.3725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.985 4.2375 320.12 4.3725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  322.845 4.2375 322.98 4.3725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.705 4.2375 325.84 4.3725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.565 4.2375 328.7 4.3725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.425 4.2375 331.56 4.3725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.285 4.2375 334.42 4.3725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.145 4.2375 337.28 4.3725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.005 4.2375 340.14 4.3725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.865 4.2375 343.0 4.3725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.725 4.2375 345.86 4.3725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.585 4.2375 348.72 4.3725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  351.445 4.2375 351.58 4.3725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.305 4.2375 354.44 4.3725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.165 4.2375 357.3 4.3725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.025 4.2375 360.16 4.3725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.885 4.2375 363.02 4.3725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.745 4.2375 365.88 4.3725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.605 4.2375 368.74 4.3725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  371.465 4.2375 371.6 4.3725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.325 4.2375 374.46 4.3725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.185 4.2375 377.32 4.3725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.045 4.2375 380.18 4.3725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  382.905 4.2375 383.04 4.3725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  385.765 4.2375 385.9 4.3725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  388.625 4.2375 388.76 4.3725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  391.485 4.2375 391.62 4.3725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.345 4.2375 394.48 4.3725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.205 4.2375 397.34 4.3725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.065 4.2375 400.2 4.3725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  402.925 4.2375 403.06 4.3725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  405.785 4.2375 405.92 4.3725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  408.645 4.2375 408.78 4.3725 ;
      END
   END din0[127]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.705 57.5625 39.84 57.6975 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.705 60.2925 39.84 60.4275 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.705 62.5025 39.84 62.6375 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.705 65.2325 39.84 65.3675 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.705 67.4425 39.84 67.5775 ;
      END
   END addr0[4]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.945 34.4225 237.08 34.5575 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.945 31.6925 237.08 31.8275 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.945 29.4825 237.08 29.6175 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.945 26.7525 237.08 26.8875 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.945 24.5425 237.08 24.6775 ;
      END
   END addr1[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  3.32 15.9625 3.455 16.0975 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.47 98.7875 273.605 98.9225 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.2825 16.0475 9.4175 16.1825 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.3675 98.7025 267.5025 98.8375 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.0625 92.08 63.1975 92.215 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.2375 92.08 64.3725 92.215 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.4125 92.08 65.5475 92.215 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.5875 92.08 66.7225 92.215 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.7625 92.08 67.8975 92.215 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.9375 92.08 69.0725 92.215 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.1125 92.08 70.2475 92.215 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.2875 92.08 71.4225 92.215 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.4625 92.08 72.5975 92.215 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.6375 92.08 73.7725 92.215 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.8125 92.08 74.9475 92.215 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.9875 92.08 76.1225 92.215 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.1625 92.08 77.2975 92.215 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.3375 92.08 78.4725 92.215 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.5125 92.08 79.6475 92.215 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.6875 92.08 80.8225 92.215 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.8625 92.08 81.9975 92.215 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.0375 92.08 83.1725 92.215 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.2125 92.08 84.3475 92.215 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.3875 92.08 85.5225 92.215 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.5625 92.08 86.6975 92.215 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.7375 92.08 87.8725 92.215 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.9125 92.08 89.0475 92.215 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.0875 92.08 90.2225 92.215 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.2625 92.08 91.3975 92.215 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.4375 92.08 92.5725 92.215 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.6125 92.08 93.7475 92.215 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.7875 92.08 94.9225 92.215 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.9625 92.08 96.0975 92.215 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.1375 92.08 97.2725 92.215 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.3125 92.08 98.4475 92.215 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.4875 92.08 99.6225 92.215 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.6625 92.08 100.7975 92.215 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.8375 92.08 101.9725 92.215 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.0125 92.08 103.1475 92.215 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.1875 92.08 104.3225 92.215 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.3625 92.08 105.4975 92.215 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.5375 92.08 106.6725 92.215 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.7125 92.08 107.8475 92.215 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.8875 92.08 109.0225 92.215 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.0625 92.08 110.1975 92.215 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.2375 92.08 111.3725 92.215 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.4125 92.08 112.5475 92.215 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.5875 92.08 113.7225 92.215 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.7625 92.08 114.8975 92.215 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.9375 92.08 116.0725 92.215 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.1125 92.08 117.2475 92.215 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.2875 92.08 118.4225 92.215 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.4625 92.08 119.5975 92.215 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.6375 92.08 120.7725 92.215 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.8125 92.08 121.9475 92.215 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.9875 92.08 123.1225 92.215 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.1625 92.08 124.2975 92.215 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.3375 92.08 125.4725 92.215 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.5125 92.08 126.6475 92.215 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.6875 92.08 127.8225 92.215 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.8625 92.08 128.9975 92.215 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.0375 92.08 130.1725 92.215 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.2125 92.08 131.3475 92.215 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.3875 92.08 132.5225 92.215 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.5625 92.08 133.6975 92.215 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.7375 92.08 134.8725 92.215 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.9125 92.08 136.0475 92.215 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.0875 92.08 137.2225 92.215 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.2625 92.08 138.3975 92.215 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.4375 92.08 139.5725 92.215 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.6125 92.08 140.7475 92.215 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.7875 92.08 141.9225 92.215 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.9625 92.08 143.0975 92.215 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.1375 92.08 144.2725 92.215 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.3125 92.08 145.4475 92.215 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.4875 92.08 146.6225 92.215 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.6625 92.08 147.7975 92.215 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.8375 92.08 148.9725 92.215 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.0125 92.08 150.1475 92.215 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.1875 92.08 151.3225 92.215 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.3625 92.08 152.4975 92.215 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.5375 92.08 153.6725 92.215 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.7125 92.08 154.8475 92.215 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.8875 92.08 156.0225 92.215 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.0625 92.08 157.1975 92.215 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.2375 92.08 158.3725 92.215 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.4125 92.08 159.5475 92.215 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.5875 92.08 160.7225 92.215 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.7625 92.08 161.8975 92.215 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.9375 92.08 163.0725 92.215 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.1125 92.08 164.2475 92.215 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.2875 92.08 165.4225 92.215 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.4625 92.08 166.5975 92.215 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.6375 92.08 167.7725 92.215 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.8125 92.08 168.9475 92.215 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.9875 92.08 170.1225 92.215 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.1625 92.08 171.2975 92.215 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.3375 92.08 172.4725 92.215 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.5125 92.08 173.6475 92.215 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.6875 92.08 174.8225 92.215 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.8625 92.08 175.9975 92.215 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.0375 92.08 177.1725 92.215 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.2125 92.08 178.3475 92.215 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.3875 92.08 179.5225 92.215 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.5625 92.08 180.6975 92.215 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.7375 92.08 181.8725 92.215 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.9125 92.08 183.0475 92.215 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.0875 92.08 184.2225 92.215 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.2625 92.08 185.3975 92.215 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.4375 92.08 186.5725 92.215 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.6125 92.08 187.7475 92.215 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.7875 92.08 188.9225 92.215 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.9625 92.08 190.0975 92.215 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.1375 92.08 191.2725 92.215 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.3125 92.08 192.4475 92.215 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.4875 92.08 193.6225 92.215 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.6625 92.08 194.7975 92.215 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.8375 92.08 195.9725 92.215 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.0125 92.08 197.1475 92.215 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.1875 92.08 198.3225 92.215 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.3625 92.08 199.4975 92.215 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.5375 92.08 200.6725 92.215 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.7125 92.08 201.8475 92.215 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.8875 92.08 203.0225 92.215 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.0625 92.08 204.1975 92.215 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.2375 92.08 205.3725 92.215 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.4125 92.08 206.5475 92.215 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.5875 92.08 207.7225 92.215 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.7625 92.08 208.8975 92.215 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.9375 92.08 210.0725 92.215 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.1125 92.08 211.2475 92.215 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.2875 92.08 212.4225 92.215 ;
      END
   END dout1[127]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  1.4 101.08 413.14 101.78 ;
         LAYER metal3 ;
         RECT  1.4 1.4 413.14 2.1 ;
         LAYER metal4 ;
         RECT  412.44 1.4 413.14 101.78 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 101.78 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 0.0 414.54 0.7 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 103.18 ;
         LAYER metal3 ;
         RECT  0.0 102.48 414.54 103.18 ;
         LAYER metal4 ;
         RECT  413.84 0.0 414.54 103.18 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 414.4 103.04 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 414.4 103.04 ;
   LAYER  metal3 ;
      RECT  0.14 4.0975 45.285 4.5125 ;
      RECT  45.7 4.0975 48.145 4.5125 ;
      RECT  48.56 4.0975 51.005 4.5125 ;
      RECT  51.42 4.0975 53.865 4.5125 ;
      RECT  54.28 4.0975 56.725 4.5125 ;
      RECT  57.14 4.0975 59.585 4.5125 ;
      RECT  60.0 4.0975 62.445 4.5125 ;
      RECT  62.86 4.0975 65.305 4.5125 ;
      RECT  65.72 4.0975 68.165 4.5125 ;
      RECT  68.58 4.0975 71.025 4.5125 ;
      RECT  71.44 4.0975 73.885 4.5125 ;
      RECT  74.3 4.0975 76.745 4.5125 ;
      RECT  77.16 4.0975 79.605 4.5125 ;
      RECT  80.02 4.0975 82.465 4.5125 ;
      RECT  82.88 4.0975 85.325 4.5125 ;
      RECT  85.74 4.0975 88.185 4.5125 ;
      RECT  88.6 4.0975 91.045 4.5125 ;
      RECT  91.46 4.0975 93.905 4.5125 ;
      RECT  94.32 4.0975 96.765 4.5125 ;
      RECT  97.18 4.0975 99.625 4.5125 ;
      RECT  100.04 4.0975 102.485 4.5125 ;
      RECT  102.9 4.0975 105.345 4.5125 ;
      RECT  105.76 4.0975 108.205 4.5125 ;
      RECT  108.62 4.0975 111.065 4.5125 ;
      RECT  111.48 4.0975 113.925 4.5125 ;
      RECT  114.34 4.0975 116.785 4.5125 ;
      RECT  117.2 4.0975 119.645 4.5125 ;
      RECT  120.06 4.0975 122.505 4.5125 ;
      RECT  122.92 4.0975 125.365 4.5125 ;
      RECT  125.78 4.0975 128.225 4.5125 ;
      RECT  128.64 4.0975 131.085 4.5125 ;
      RECT  131.5 4.0975 133.945 4.5125 ;
      RECT  134.36 4.0975 136.805 4.5125 ;
      RECT  137.22 4.0975 139.665 4.5125 ;
      RECT  140.08 4.0975 142.525 4.5125 ;
      RECT  142.94 4.0975 145.385 4.5125 ;
      RECT  145.8 4.0975 148.245 4.5125 ;
      RECT  148.66 4.0975 151.105 4.5125 ;
      RECT  151.52 4.0975 153.965 4.5125 ;
      RECT  154.38 4.0975 156.825 4.5125 ;
      RECT  157.24 4.0975 159.685 4.5125 ;
      RECT  160.1 4.0975 162.545 4.5125 ;
      RECT  162.96 4.0975 165.405 4.5125 ;
      RECT  165.82 4.0975 168.265 4.5125 ;
      RECT  168.68 4.0975 171.125 4.5125 ;
      RECT  171.54 4.0975 173.985 4.5125 ;
      RECT  174.4 4.0975 176.845 4.5125 ;
      RECT  177.26 4.0975 179.705 4.5125 ;
      RECT  180.12 4.0975 182.565 4.5125 ;
      RECT  182.98 4.0975 185.425 4.5125 ;
      RECT  185.84 4.0975 188.285 4.5125 ;
      RECT  188.7 4.0975 191.145 4.5125 ;
      RECT  191.56 4.0975 194.005 4.5125 ;
      RECT  194.42 4.0975 196.865 4.5125 ;
      RECT  197.28 4.0975 199.725 4.5125 ;
      RECT  200.14 4.0975 202.585 4.5125 ;
      RECT  203.0 4.0975 205.445 4.5125 ;
      RECT  205.86 4.0975 208.305 4.5125 ;
      RECT  208.72 4.0975 211.165 4.5125 ;
      RECT  211.58 4.0975 214.025 4.5125 ;
      RECT  214.44 4.0975 216.885 4.5125 ;
      RECT  217.3 4.0975 219.745 4.5125 ;
      RECT  220.16 4.0975 222.605 4.5125 ;
      RECT  223.02 4.0975 225.465 4.5125 ;
      RECT  225.88 4.0975 228.325 4.5125 ;
      RECT  228.74 4.0975 231.185 4.5125 ;
      RECT  231.6 4.0975 234.045 4.5125 ;
      RECT  234.46 4.0975 236.905 4.5125 ;
      RECT  237.32 4.0975 239.765 4.5125 ;
      RECT  240.18 4.0975 242.625 4.5125 ;
      RECT  243.04 4.0975 245.485 4.5125 ;
      RECT  245.9 4.0975 248.345 4.5125 ;
      RECT  248.76 4.0975 251.205 4.5125 ;
      RECT  251.62 4.0975 254.065 4.5125 ;
      RECT  254.48 4.0975 256.925 4.5125 ;
      RECT  257.34 4.0975 259.785 4.5125 ;
      RECT  260.2 4.0975 262.645 4.5125 ;
      RECT  263.06 4.0975 265.505 4.5125 ;
      RECT  265.92 4.0975 268.365 4.5125 ;
      RECT  268.78 4.0975 271.225 4.5125 ;
      RECT  271.64 4.0975 274.085 4.5125 ;
      RECT  274.5 4.0975 276.945 4.5125 ;
      RECT  277.36 4.0975 279.805 4.5125 ;
      RECT  280.22 4.0975 282.665 4.5125 ;
      RECT  283.08 4.0975 285.525 4.5125 ;
      RECT  285.94 4.0975 288.385 4.5125 ;
      RECT  288.8 4.0975 291.245 4.5125 ;
      RECT  291.66 4.0975 294.105 4.5125 ;
      RECT  294.52 4.0975 296.965 4.5125 ;
      RECT  297.38 4.0975 299.825 4.5125 ;
      RECT  300.24 4.0975 302.685 4.5125 ;
      RECT  303.1 4.0975 305.545 4.5125 ;
      RECT  305.96 4.0975 308.405 4.5125 ;
      RECT  308.82 4.0975 311.265 4.5125 ;
      RECT  311.68 4.0975 314.125 4.5125 ;
      RECT  314.54 4.0975 316.985 4.5125 ;
      RECT  317.4 4.0975 319.845 4.5125 ;
      RECT  320.26 4.0975 322.705 4.5125 ;
      RECT  323.12 4.0975 325.565 4.5125 ;
      RECT  325.98 4.0975 328.425 4.5125 ;
      RECT  328.84 4.0975 331.285 4.5125 ;
      RECT  331.7 4.0975 334.145 4.5125 ;
      RECT  334.56 4.0975 337.005 4.5125 ;
      RECT  337.42 4.0975 339.865 4.5125 ;
      RECT  340.28 4.0975 342.725 4.5125 ;
      RECT  343.14 4.0975 345.585 4.5125 ;
      RECT  346.0 4.0975 348.445 4.5125 ;
      RECT  348.86 4.0975 351.305 4.5125 ;
      RECT  351.72 4.0975 354.165 4.5125 ;
      RECT  354.58 4.0975 357.025 4.5125 ;
      RECT  357.44 4.0975 359.885 4.5125 ;
      RECT  360.3 4.0975 362.745 4.5125 ;
      RECT  363.16 4.0975 365.605 4.5125 ;
      RECT  366.02 4.0975 368.465 4.5125 ;
      RECT  368.88 4.0975 371.325 4.5125 ;
      RECT  371.74 4.0975 374.185 4.5125 ;
      RECT  374.6 4.0975 377.045 4.5125 ;
      RECT  377.46 4.0975 379.905 4.5125 ;
      RECT  380.32 4.0975 382.765 4.5125 ;
      RECT  383.18 4.0975 385.625 4.5125 ;
      RECT  386.04 4.0975 388.485 4.5125 ;
      RECT  388.9 4.0975 391.345 4.5125 ;
      RECT  391.76 4.0975 394.205 4.5125 ;
      RECT  394.62 4.0975 397.065 4.5125 ;
      RECT  397.48 4.0975 399.925 4.5125 ;
      RECT  400.34 4.0975 402.785 4.5125 ;
      RECT  403.2 4.0975 405.645 4.5125 ;
      RECT  406.06 4.0975 408.505 4.5125 ;
      RECT  408.92 4.0975 414.4 4.5125 ;
      RECT  0.14 57.4225 39.565 57.8375 ;
      RECT  39.565 4.5125 39.98 57.4225 ;
      RECT  39.98 4.5125 45.285 57.4225 ;
      RECT  39.98 57.4225 45.285 57.8375 ;
      RECT  39.565 57.8375 39.98 60.1525 ;
      RECT  39.565 60.5675 39.98 62.3625 ;
      RECT  39.565 62.7775 39.98 65.0925 ;
      RECT  39.565 65.5075 39.98 67.3025 ;
      RECT  45.7 4.5125 236.805 34.2825 ;
      RECT  45.7 34.2825 236.805 34.6975 ;
      RECT  237.22 4.5125 414.4 34.2825 ;
      RECT  237.22 34.2825 414.4 34.6975 ;
      RECT  236.805 31.9675 237.22 34.2825 ;
      RECT  236.805 29.7575 237.22 31.5525 ;
      RECT  236.805 27.0275 237.22 29.3425 ;
      RECT  236.805 4.5125 237.22 24.4025 ;
      RECT  236.805 24.8175 237.22 26.6125 ;
      RECT  0.14 4.5125 3.18 15.8225 ;
      RECT  0.14 15.8225 3.18 16.2375 ;
      RECT  0.14 16.2375 3.18 57.4225 ;
      RECT  3.18 4.5125 3.595 15.8225 ;
      RECT  3.18 16.2375 3.595 57.4225 ;
      RECT  3.595 4.5125 39.565 15.8225 ;
      RECT  273.33 34.6975 273.745 98.6475 ;
      RECT  273.745 34.6975 414.4 98.6475 ;
      RECT  273.745 98.6475 414.4 99.0625 ;
      RECT  3.595 15.8225 9.1425 15.9075 ;
      RECT  3.595 15.9075 9.1425 16.2375 ;
      RECT  9.1425 15.8225 9.5575 15.9075 ;
      RECT  9.5575 15.8225 39.565 15.9075 ;
      RECT  9.5575 15.9075 39.565 16.2375 ;
      RECT  3.595 16.2375 9.1425 16.3225 ;
      RECT  3.595 16.3225 9.1425 57.4225 ;
      RECT  9.1425 16.3225 9.5575 57.4225 ;
      RECT  9.5575 16.2375 39.565 16.3225 ;
      RECT  9.5575 16.3225 39.565 57.4225 ;
      RECT  237.22 34.6975 267.2275 98.5625 ;
      RECT  237.22 98.5625 267.2275 98.6475 ;
      RECT  267.2275 34.6975 267.6425 98.5625 ;
      RECT  267.6425 34.6975 273.33 98.5625 ;
      RECT  267.6425 98.5625 273.33 98.6475 ;
      RECT  237.22 98.6475 267.2275 98.9775 ;
      RECT  237.22 98.9775 267.2275 99.0625 ;
      RECT  267.2275 98.9775 267.6425 99.0625 ;
      RECT  267.6425 98.6475 273.33 98.9775 ;
      RECT  267.6425 98.9775 273.33 99.0625 ;
      RECT  45.7 34.6975 62.9225 91.94 ;
      RECT  45.7 91.94 62.9225 92.355 ;
      RECT  62.9225 34.6975 63.3375 91.94 ;
      RECT  63.3375 34.6975 236.805 91.94 ;
      RECT  63.3375 91.94 64.0975 92.355 ;
      RECT  64.5125 91.94 65.2725 92.355 ;
      RECT  65.6875 91.94 66.4475 92.355 ;
      RECT  66.8625 91.94 67.6225 92.355 ;
      RECT  68.0375 91.94 68.7975 92.355 ;
      RECT  69.2125 91.94 69.9725 92.355 ;
      RECT  70.3875 91.94 71.1475 92.355 ;
      RECT  71.5625 91.94 72.3225 92.355 ;
      RECT  72.7375 91.94 73.4975 92.355 ;
      RECT  73.9125 91.94 74.6725 92.355 ;
      RECT  75.0875 91.94 75.8475 92.355 ;
      RECT  76.2625 91.94 77.0225 92.355 ;
      RECT  77.4375 91.94 78.1975 92.355 ;
      RECT  78.6125 91.94 79.3725 92.355 ;
      RECT  79.7875 91.94 80.5475 92.355 ;
      RECT  80.9625 91.94 81.7225 92.355 ;
      RECT  82.1375 91.94 82.8975 92.355 ;
      RECT  83.3125 91.94 84.0725 92.355 ;
      RECT  84.4875 91.94 85.2475 92.355 ;
      RECT  85.6625 91.94 86.4225 92.355 ;
      RECT  86.8375 91.94 87.5975 92.355 ;
      RECT  88.0125 91.94 88.7725 92.355 ;
      RECT  89.1875 91.94 89.9475 92.355 ;
      RECT  90.3625 91.94 91.1225 92.355 ;
      RECT  91.5375 91.94 92.2975 92.355 ;
      RECT  92.7125 91.94 93.4725 92.355 ;
      RECT  93.8875 91.94 94.6475 92.355 ;
      RECT  95.0625 91.94 95.8225 92.355 ;
      RECT  96.2375 91.94 96.9975 92.355 ;
      RECT  97.4125 91.94 98.1725 92.355 ;
      RECT  98.5875 91.94 99.3475 92.355 ;
      RECT  99.7625 91.94 100.5225 92.355 ;
      RECT  100.9375 91.94 101.6975 92.355 ;
      RECT  102.1125 91.94 102.8725 92.355 ;
      RECT  103.2875 91.94 104.0475 92.355 ;
      RECT  104.4625 91.94 105.2225 92.355 ;
      RECT  105.6375 91.94 106.3975 92.355 ;
      RECT  106.8125 91.94 107.5725 92.355 ;
      RECT  107.9875 91.94 108.7475 92.355 ;
      RECT  109.1625 91.94 109.9225 92.355 ;
      RECT  110.3375 91.94 111.0975 92.355 ;
      RECT  111.5125 91.94 112.2725 92.355 ;
      RECT  112.6875 91.94 113.4475 92.355 ;
      RECT  113.8625 91.94 114.6225 92.355 ;
      RECT  115.0375 91.94 115.7975 92.355 ;
      RECT  116.2125 91.94 116.9725 92.355 ;
      RECT  117.3875 91.94 118.1475 92.355 ;
      RECT  118.5625 91.94 119.3225 92.355 ;
      RECT  119.7375 91.94 120.4975 92.355 ;
      RECT  120.9125 91.94 121.6725 92.355 ;
      RECT  122.0875 91.94 122.8475 92.355 ;
      RECT  123.2625 91.94 124.0225 92.355 ;
      RECT  124.4375 91.94 125.1975 92.355 ;
      RECT  125.6125 91.94 126.3725 92.355 ;
      RECT  126.7875 91.94 127.5475 92.355 ;
      RECT  127.9625 91.94 128.7225 92.355 ;
      RECT  129.1375 91.94 129.8975 92.355 ;
      RECT  130.3125 91.94 131.0725 92.355 ;
      RECT  131.4875 91.94 132.2475 92.355 ;
      RECT  132.6625 91.94 133.4225 92.355 ;
      RECT  133.8375 91.94 134.5975 92.355 ;
      RECT  135.0125 91.94 135.7725 92.355 ;
      RECT  136.1875 91.94 136.9475 92.355 ;
      RECT  137.3625 91.94 138.1225 92.355 ;
      RECT  138.5375 91.94 139.2975 92.355 ;
      RECT  139.7125 91.94 140.4725 92.355 ;
      RECT  140.8875 91.94 141.6475 92.355 ;
      RECT  142.0625 91.94 142.8225 92.355 ;
      RECT  143.2375 91.94 143.9975 92.355 ;
      RECT  144.4125 91.94 145.1725 92.355 ;
      RECT  145.5875 91.94 146.3475 92.355 ;
      RECT  146.7625 91.94 147.5225 92.355 ;
      RECT  147.9375 91.94 148.6975 92.355 ;
      RECT  149.1125 91.94 149.8725 92.355 ;
      RECT  150.2875 91.94 151.0475 92.355 ;
      RECT  151.4625 91.94 152.2225 92.355 ;
      RECT  152.6375 91.94 153.3975 92.355 ;
      RECT  153.8125 91.94 154.5725 92.355 ;
      RECT  154.9875 91.94 155.7475 92.355 ;
      RECT  156.1625 91.94 156.9225 92.355 ;
      RECT  157.3375 91.94 158.0975 92.355 ;
      RECT  158.5125 91.94 159.2725 92.355 ;
      RECT  159.6875 91.94 160.4475 92.355 ;
      RECT  160.8625 91.94 161.6225 92.355 ;
      RECT  162.0375 91.94 162.7975 92.355 ;
      RECT  163.2125 91.94 163.9725 92.355 ;
      RECT  164.3875 91.94 165.1475 92.355 ;
      RECT  165.5625 91.94 166.3225 92.355 ;
      RECT  166.7375 91.94 167.4975 92.355 ;
      RECT  167.9125 91.94 168.6725 92.355 ;
      RECT  169.0875 91.94 169.8475 92.355 ;
      RECT  170.2625 91.94 171.0225 92.355 ;
      RECT  171.4375 91.94 172.1975 92.355 ;
      RECT  172.6125 91.94 173.3725 92.355 ;
      RECT  173.7875 91.94 174.5475 92.355 ;
      RECT  174.9625 91.94 175.7225 92.355 ;
      RECT  176.1375 91.94 176.8975 92.355 ;
      RECT  177.3125 91.94 178.0725 92.355 ;
      RECT  178.4875 91.94 179.2475 92.355 ;
      RECT  179.6625 91.94 180.4225 92.355 ;
      RECT  180.8375 91.94 181.5975 92.355 ;
      RECT  182.0125 91.94 182.7725 92.355 ;
      RECT  183.1875 91.94 183.9475 92.355 ;
      RECT  184.3625 91.94 185.1225 92.355 ;
      RECT  185.5375 91.94 186.2975 92.355 ;
      RECT  186.7125 91.94 187.4725 92.355 ;
      RECT  187.8875 91.94 188.6475 92.355 ;
      RECT  189.0625 91.94 189.8225 92.355 ;
      RECT  190.2375 91.94 190.9975 92.355 ;
      RECT  191.4125 91.94 192.1725 92.355 ;
      RECT  192.5875 91.94 193.3475 92.355 ;
      RECT  193.7625 91.94 194.5225 92.355 ;
      RECT  194.9375 91.94 195.6975 92.355 ;
      RECT  196.1125 91.94 196.8725 92.355 ;
      RECT  197.2875 91.94 198.0475 92.355 ;
      RECT  198.4625 91.94 199.2225 92.355 ;
      RECT  199.6375 91.94 200.3975 92.355 ;
      RECT  200.8125 91.94 201.5725 92.355 ;
      RECT  201.9875 91.94 202.7475 92.355 ;
      RECT  203.1625 91.94 203.9225 92.355 ;
      RECT  204.3375 91.94 205.0975 92.355 ;
      RECT  205.5125 91.94 206.2725 92.355 ;
      RECT  206.6875 91.94 207.4475 92.355 ;
      RECT  207.8625 91.94 208.6225 92.355 ;
      RECT  209.0375 91.94 209.7975 92.355 ;
      RECT  210.2125 91.94 210.9725 92.355 ;
      RECT  211.3875 91.94 212.1475 92.355 ;
      RECT  212.5625 91.94 236.805 92.355 ;
      RECT  45.285 4.5125 45.7 100.94 ;
      RECT  0.14 57.8375 1.26 100.94 ;
      RECT  0.14 100.94 1.26 101.92 ;
      RECT  1.26 57.8375 39.565 100.94 ;
      RECT  39.98 57.8375 45.285 100.94 ;
      RECT  39.565 67.7175 39.98 100.94 ;
      RECT  236.805 34.6975 237.22 100.94 ;
      RECT  237.22 99.0625 273.33 100.94 ;
      RECT  273.33 99.0625 273.745 100.94 ;
      RECT  273.745 99.0625 413.28 100.94 ;
      RECT  413.28 99.0625 414.4 100.94 ;
      RECT  413.28 100.94 414.4 101.92 ;
      RECT  45.7 92.355 62.9225 100.94 ;
      RECT  62.9225 92.355 63.3375 100.94 ;
      RECT  63.3375 92.355 236.805 100.94 ;
      RECT  0.14 1.26 1.26 2.24 ;
      RECT  0.14 2.24 1.26 4.0975 ;
      RECT  1.26 2.24 45.285 4.0975 ;
      RECT  45.285 2.24 45.7 4.0975 ;
      RECT  45.7 2.24 413.28 4.0975 ;
      RECT  413.28 1.26 414.4 2.24 ;
      RECT  413.28 2.24 414.4 4.0975 ;
      RECT  0.14 0.84 1.26 1.26 ;
      RECT  1.26 0.84 45.285 1.26 ;
      RECT  45.285 0.84 45.7 1.26 ;
      RECT  45.7 0.84 413.28 1.26 ;
      RECT  413.28 0.84 414.4 1.26 ;
      RECT  45.285 101.92 45.7 102.34 ;
      RECT  0.14 101.92 1.26 102.34 ;
      RECT  1.26 101.92 39.565 102.34 ;
      RECT  39.98 101.92 45.285 102.34 ;
      RECT  39.565 101.92 39.98 102.34 ;
      RECT  236.805 101.92 237.22 102.34 ;
      RECT  237.22 101.92 273.33 102.34 ;
      RECT  273.33 101.92 273.745 102.34 ;
      RECT  273.745 101.92 413.28 102.34 ;
      RECT  413.28 101.92 414.4 102.34 ;
      RECT  45.7 101.92 62.9225 102.34 ;
      RECT  62.9225 101.92 63.3375 102.34 ;
      RECT  63.3375 101.92 236.805 102.34 ;
   LAYER  metal4 ;
      RECT  412.16 0.14 413.42 1.12 ;
      RECT  412.16 102.06 413.42 103.04 ;
      RECT  2.38 1.12 412.16 102.06 ;
      RECT  0.98 0.14 412.16 1.12 ;
      RECT  0.98 102.06 412.16 103.04 ;
      RECT  0.98 1.12 1.12 102.06 ;
      RECT  413.42 0.14 413.56 1.12 ;
      RECT  413.42 1.12 413.56 102.06 ;
      RECT  413.42 102.06 413.56 103.04 ;
   END
END    freepdk45_sram_1w1r_31x128
END    LIBRARY
