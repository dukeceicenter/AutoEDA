VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_64x512
   CLASS BLOCK ;
   SIZE 1593.34 BY 214.34 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.065 4.2375 126.2 4.3725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.925 4.2375 129.06 4.3725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.785 4.2375 131.92 4.3725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.645 4.2375 134.78 4.3725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.505 4.2375 137.64 4.3725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.365 4.2375 140.5 4.3725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.225 4.2375 143.36 4.3725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.085 4.2375 146.22 4.3725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.945 4.2375 149.08 4.3725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.805 4.2375 151.94 4.3725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.665 4.2375 154.8 4.3725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.525 4.2375 157.66 4.3725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.385 4.2375 160.52 4.3725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.245 4.2375 163.38 4.3725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.105 4.2375 166.24 4.3725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.965 4.2375 169.1 4.3725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.825 4.2375 171.96 4.3725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.685 4.2375 174.82 4.3725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.545 4.2375 177.68 4.3725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.405 4.2375 180.54 4.3725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.265 4.2375 183.4 4.3725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.125 4.2375 186.26 4.3725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.985 4.2375 189.12 4.3725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.845 4.2375 191.98 4.3725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.705 4.2375 194.84 4.3725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.565 4.2375 197.7 4.3725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.425 4.2375 200.56 4.3725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.285 4.2375 203.42 4.3725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.145 4.2375 206.28 4.3725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.005 4.2375 209.14 4.3725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.865 4.2375 212.0 4.3725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.725 4.2375 214.86 4.3725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.585 4.2375 217.72 4.3725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.445 4.2375 220.58 4.3725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.305 4.2375 223.44 4.3725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.165 4.2375 226.3 4.3725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.025 4.2375 229.16 4.3725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.885 4.2375 232.02 4.3725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.745 4.2375 234.88 4.3725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.605 4.2375 237.74 4.3725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.465 4.2375 240.6 4.3725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.325 4.2375 243.46 4.3725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.185 4.2375 246.32 4.3725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.045 4.2375 249.18 4.3725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.905 4.2375 252.04 4.3725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.765 4.2375 254.9 4.3725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.625 4.2375 257.76 4.3725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.485 4.2375 260.62 4.3725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.345 4.2375 263.48 4.3725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.205 4.2375 266.34 4.3725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.065 4.2375 269.2 4.3725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.925 4.2375 272.06 4.3725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.785 4.2375 274.92 4.3725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.645 4.2375 277.78 4.3725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.505 4.2375 280.64 4.3725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.365 4.2375 283.5 4.3725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.225 4.2375 286.36 4.3725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.085 4.2375 289.22 4.3725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.945 4.2375 292.08 4.3725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.805 4.2375 294.94 4.3725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.665 4.2375 297.8 4.3725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.525 4.2375 300.66 4.3725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.385 4.2375 303.52 4.3725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.245 4.2375 306.38 4.3725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.105 4.2375 309.24 4.3725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.965 4.2375 312.1 4.3725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.825 4.2375 314.96 4.3725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.685 4.2375 317.82 4.3725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.545 4.2375 320.68 4.3725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.405 4.2375 323.54 4.3725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.265 4.2375 326.4 4.3725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.125 4.2375 329.26 4.3725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.985 4.2375 332.12 4.3725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.845 4.2375 334.98 4.3725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.705 4.2375 337.84 4.3725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.565 4.2375 340.7 4.3725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.425 4.2375 343.56 4.3725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.285 4.2375 346.42 4.3725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.145 4.2375 349.28 4.3725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.005 4.2375 352.14 4.3725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.865 4.2375 355.0 4.3725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.725 4.2375 357.86 4.3725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.585 4.2375 360.72 4.3725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.445 4.2375 363.58 4.3725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.305 4.2375 366.44 4.3725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.165 4.2375 369.3 4.3725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.025 4.2375 372.16 4.3725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.885 4.2375 375.02 4.3725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.745 4.2375 377.88 4.3725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.605 4.2375 380.74 4.3725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.465 4.2375 383.6 4.3725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.325 4.2375 386.46 4.3725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.185 4.2375 389.32 4.3725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.045 4.2375 392.18 4.3725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.905 4.2375 395.04 4.3725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.765 4.2375 397.9 4.3725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.625 4.2375 400.76 4.3725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.485 4.2375 403.62 4.3725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.345 4.2375 406.48 4.3725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.205 4.2375 409.34 4.3725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.065 4.2375 412.2 4.3725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  414.925 4.2375 415.06 4.3725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.785 4.2375 417.92 4.3725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.645 4.2375 420.78 4.3725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.505 4.2375 423.64 4.3725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.365 4.2375 426.5 4.3725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.225 4.2375 429.36 4.3725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.085 4.2375 432.22 4.3725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  434.945 4.2375 435.08 4.3725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  437.805 4.2375 437.94 4.3725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.665 4.2375 440.8 4.3725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.525 4.2375 443.66 4.3725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.385 4.2375 446.52 4.3725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.245 4.2375 449.38 4.3725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.105 4.2375 452.24 4.3725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  454.965 4.2375 455.1 4.3725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  457.825 4.2375 457.96 4.3725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  460.685 4.2375 460.82 4.3725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  463.545 4.2375 463.68 4.3725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.405 4.2375 466.54 4.3725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.265 4.2375 469.4 4.3725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.125 4.2375 472.26 4.3725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  474.985 4.2375 475.12 4.3725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  477.845 4.2375 477.98 4.3725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  480.705 4.2375 480.84 4.3725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  483.565 4.2375 483.7 4.3725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.425 4.2375 486.56 4.3725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.285 4.2375 489.42 4.3725 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.145 4.2375 492.28 4.3725 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.005 4.2375 495.14 4.3725 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  497.865 4.2375 498.0 4.3725 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  500.725 4.2375 500.86 4.3725 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  503.585 4.2375 503.72 4.3725 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  506.445 4.2375 506.58 4.3725 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.305 4.2375 509.44 4.3725 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.165 4.2375 512.3 4.3725 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.025 4.2375 515.16 4.3725 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  517.885 4.2375 518.02 4.3725 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  520.745 4.2375 520.88 4.3725 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  523.605 4.2375 523.74 4.3725 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  526.465 4.2375 526.6 4.3725 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  529.325 4.2375 529.46 4.3725 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  532.185 4.2375 532.32 4.3725 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  535.045 4.2375 535.18 4.3725 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  537.905 4.2375 538.04 4.3725 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  540.765 4.2375 540.9 4.3725 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  543.625 4.2375 543.76 4.3725 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  546.485 4.2375 546.62 4.3725 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  549.345 4.2375 549.48 4.3725 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  552.205 4.2375 552.34 4.3725 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  555.065 4.2375 555.2 4.3725 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  557.925 4.2375 558.06 4.3725 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  560.785 4.2375 560.92 4.3725 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  563.645 4.2375 563.78 4.3725 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  566.505 4.2375 566.64 4.3725 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  569.365 4.2375 569.5 4.3725 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  572.225 4.2375 572.36 4.3725 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  575.085 4.2375 575.22 4.3725 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  577.945 4.2375 578.08 4.3725 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  580.805 4.2375 580.94 4.3725 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  583.665 4.2375 583.8 4.3725 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  586.525 4.2375 586.66 4.3725 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  589.385 4.2375 589.52 4.3725 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  592.245 4.2375 592.38 4.3725 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  595.105 4.2375 595.24 4.3725 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  597.965 4.2375 598.1 4.3725 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  600.825 4.2375 600.96 4.3725 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  603.685 4.2375 603.82 4.3725 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  606.545 4.2375 606.68 4.3725 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  609.405 4.2375 609.54 4.3725 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  612.265 4.2375 612.4 4.3725 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  615.125 4.2375 615.26 4.3725 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  617.985 4.2375 618.12 4.3725 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  620.845 4.2375 620.98 4.3725 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  623.705 4.2375 623.84 4.3725 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  626.565 4.2375 626.7 4.3725 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  629.425 4.2375 629.56 4.3725 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  632.285 4.2375 632.42 4.3725 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  635.145 4.2375 635.28 4.3725 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  638.005 4.2375 638.14 4.3725 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  640.865 4.2375 641.0 4.3725 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  643.725 4.2375 643.86 4.3725 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  646.585 4.2375 646.72 4.3725 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  649.445 4.2375 649.58 4.3725 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  652.305 4.2375 652.44 4.3725 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  655.165 4.2375 655.3 4.3725 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  658.025 4.2375 658.16 4.3725 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  660.885 4.2375 661.02 4.3725 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  663.745 4.2375 663.88 4.3725 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  666.605 4.2375 666.74 4.3725 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  669.465 4.2375 669.6 4.3725 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  672.325 4.2375 672.46 4.3725 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  675.185 4.2375 675.32 4.3725 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  678.045 4.2375 678.18 4.3725 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  680.905 4.2375 681.04 4.3725 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  683.765 4.2375 683.9 4.3725 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  686.625 4.2375 686.76 4.3725 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  689.485 4.2375 689.62 4.3725 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  692.345 4.2375 692.48 4.3725 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  695.205 4.2375 695.34 4.3725 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  698.065 4.2375 698.2 4.3725 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  700.925 4.2375 701.06 4.3725 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  703.785 4.2375 703.92 4.3725 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  706.645 4.2375 706.78 4.3725 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  709.505 4.2375 709.64 4.3725 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  712.365 4.2375 712.5 4.3725 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  715.225 4.2375 715.36 4.3725 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  718.085 4.2375 718.22 4.3725 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  720.945 4.2375 721.08 4.3725 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  723.805 4.2375 723.94 4.3725 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  726.665 4.2375 726.8 4.3725 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  729.525 4.2375 729.66 4.3725 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  732.385 4.2375 732.52 4.3725 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  735.245 4.2375 735.38 4.3725 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  738.105 4.2375 738.24 4.3725 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  740.965 4.2375 741.1 4.3725 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  743.825 4.2375 743.96 4.3725 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  746.685 4.2375 746.82 4.3725 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  749.545 4.2375 749.68 4.3725 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  752.405 4.2375 752.54 4.3725 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  755.265 4.2375 755.4 4.3725 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  758.125 4.2375 758.26 4.3725 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  760.985 4.2375 761.12 4.3725 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  763.845 4.2375 763.98 4.3725 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  766.705 4.2375 766.84 4.3725 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  769.565 4.2375 769.7 4.3725 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  772.425 4.2375 772.56 4.3725 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  775.285 4.2375 775.42 4.3725 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  778.145 4.2375 778.28 4.3725 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  781.005 4.2375 781.14 4.3725 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  783.865 4.2375 784.0 4.3725 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  786.725 4.2375 786.86 4.3725 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  789.585 4.2375 789.72 4.3725 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  792.445 4.2375 792.58 4.3725 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  795.305 4.2375 795.44 4.3725 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  798.165 4.2375 798.3 4.3725 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.025 4.2375 801.16 4.3725 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  803.885 4.2375 804.02 4.3725 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  806.745 4.2375 806.88 4.3725 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  809.605 4.2375 809.74 4.3725 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  812.465 4.2375 812.6 4.3725 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  815.325 4.2375 815.46 4.3725 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  818.185 4.2375 818.32 4.3725 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  821.045 4.2375 821.18 4.3725 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  823.905 4.2375 824.04 4.3725 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  826.765 4.2375 826.9 4.3725 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  829.625 4.2375 829.76 4.3725 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  832.485 4.2375 832.62 4.3725 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  835.345 4.2375 835.48 4.3725 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  838.205 4.2375 838.34 4.3725 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  841.065 4.2375 841.2 4.3725 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  843.925 4.2375 844.06 4.3725 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  846.785 4.2375 846.92 4.3725 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  849.645 4.2375 849.78 4.3725 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  852.505 4.2375 852.64 4.3725 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  855.365 4.2375 855.5 4.3725 ;
      END
   END din0[255]
   PIN din0[256]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  858.225 4.2375 858.36 4.3725 ;
      END
   END din0[256]
   PIN din0[257]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  861.085 4.2375 861.22 4.3725 ;
      END
   END din0[257]
   PIN din0[258]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  863.945 4.2375 864.08 4.3725 ;
      END
   END din0[258]
   PIN din0[259]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  866.805 4.2375 866.94 4.3725 ;
      END
   END din0[259]
   PIN din0[260]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  869.665 4.2375 869.8 4.3725 ;
      END
   END din0[260]
   PIN din0[261]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  872.525 4.2375 872.66 4.3725 ;
      END
   END din0[261]
   PIN din0[262]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  875.385 4.2375 875.52 4.3725 ;
      END
   END din0[262]
   PIN din0[263]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  878.245 4.2375 878.38 4.3725 ;
      END
   END din0[263]
   PIN din0[264]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  881.105 4.2375 881.24 4.3725 ;
      END
   END din0[264]
   PIN din0[265]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  883.965 4.2375 884.1 4.3725 ;
      END
   END din0[265]
   PIN din0[266]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  886.825 4.2375 886.96 4.3725 ;
      END
   END din0[266]
   PIN din0[267]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  889.685 4.2375 889.82 4.3725 ;
      END
   END din0[267]
   PIN din0[268]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  892.545 4.2375 892.68 4.3725 ;
      END
   END din0[268]
   PIN din0[269]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  895.405 4.2375 895.54 4.3725 ;
      END
   END din0[269]
   PIN din0[270]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  898.265 4.2375 898.4 4.3725 ;
      END
   END din0[270]
   PIN din0[271]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  901.125 4.2375 901.26 4.3725 ;
      END
   END din0[271]
   PIN din0[272]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  903.985 4.2375 904.12 4.3725 ;
      END
   END din0[272]
   PIN din0[273]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  906.845 4.2375 906.98 4.3725 ;
      END
   END din0[273]
   PIN din0[274]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  909.705 4.2375 909.84 4.3725 ;
      END
   END din0[274]
   PIN din0[275]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  912.565 4.2375 912.7 4.3725 ;
      END
   END din0[275]
   PIN din0[276]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  915.425 4.2375 915.56 4.3725 ;
      END
   END din0[276]
   PIN din0[277]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  918.285 4.2375 918.42 4.3725 ;
      END
   END din0[277]
   PIN din0[278]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  921.145 4.2375 921.28 4.3725 ;
      END
   END din0[278]
   PIN din0[279]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  924.005 4.2375 924.14 4.3725 ;
      END
   END din0[279]
   PIN din0[280]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  926.865 4.2375 927.0 4.3725 ;
      END
   END din0[280]
   PIN din0[281]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  929.725 4.2375 929.86 4.3725 ;
      END
   END din0[281]
   PIN din0[282]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  932.585 4.2375 932.72 4.3725 ;
      END
   END din0[282]
   PIN din0[283]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  935.445 4.2375 935.58 4.3725 ;
      END
   END din0[283]
   PIN din0[284]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  938.305 4.2375 938.44 4.3725 ;
      END
   END din0[284]
   PIN din0[285]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  941.165 4.2375 941.3 4.3725 ;
      END
   END din0[285]
   PIN din0[286]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  944.025 4.2375 944.16 4.3725 ;
      END
   END din0[286]
   PIN din0[287]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  946.885 4.2375 947.02 4.3725 ;
      END
   END din0[287]
   PIN din0[288]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  949.745 4.2375 949.88 4.3725 ;
      END
   END din0[288]
   PIN din0[289]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  952.605 4.2375 952.74 4.3725 ;
      END
   END din0[289]
   PIN din0[290]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  955.465 4.2375 955.6 4.3725 ;
      END
   END din0[290]
   PIN din0[291]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  958.325 4.2375 958.46 4.3725 ;
      END
   END din0[291]
   PIN din0[292]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  961.185 4.2375 961.32 4.3725 ;
      END
   END din0[292]
   PIN din0[293]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  964.045 4.2375 964.18 4.3725 ;
      END
   END din0[293]
   PIN din0[294]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  966.905 4.2375 967.04 4.3725 ;
      END
   END din0[294]
   PIN din0[295]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  969.765 4.2375 969.9 4.3725 ;
      END
   END din0[295]
   PIN din0[296]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  972.625 4.2375 972.76 4.3725 ;
      END
   END din0[296]
   PIN din0[297]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  975.485 4.2375 975.62 4.3725 ;
      END
   END din0[297]
   PIN din0[298]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  978.345 4.2375 978.48 4.3725 ;
      END
   END din0[298]
   PIN din0[299]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  981.205 4.2375 981.34 4.3725 ;
      END
   END din0[299]
   PIN din0[300]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  984.065 4.2375 984.2 4.3725 ;
      END
   END din0[300]
   PIN din0[301]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  986.925 4.2375 987.06 4.3725 ;
      END
   END din0[301]
   PIN din0[302]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  989.785 4.2375 989.92 4.3725 ;
      END
   END din0[302]
   PIN din0[303]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  992.645 4.2375 992.78 4.3725 ;
      END
   END din0[303]
   PIN din0[304]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  995.505 4.2375 995.64 4.3725 ;
      END
   END din0[304]
   PIN din0[305]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  998.365 4.2375 998.5 4.3725 ;
      END
   END din0[305]
   PIN din0[306]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1001.225 4.2375 1001.36 4.3725 ;
      END
   END din0[306]
   PIN din0[307]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1004.085 4.2375 1004.22 4.3725 ;
      END
   END din0[307]
   PIN din0[308]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1006.945 4.2375 1007.08 4.3725 ;
      END
   END din0[308]
   PIN din0[309]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1009.805 4.2375 1009.94 4.3725 ;
      END
   END din0[309]
   PIN din0[310]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1012.665 4.2375 1012.8 4.3725 ;
      END
   END din0[310]
   PIN din0[311]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1015.525 4.2375 1015.66 4.3725 ;
      END
   END din0[311]
   PIN din0[312]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1018.385 4.2375 1018.52 4.3725 ;
      END
   END din0[312]
   PIN din0[313]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1021.245 4.2375 1021.38 4.3725 ;
      END
   END din0[313]
   PIN din0[314]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1024.105 4.2375 1024.24 4.3725 ;
      END
   END din0[314]
   PIN din0[315]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1026.965 4.2375 1027.1 4.3725 ;
      END
   END din0[315]
   PIN din0[316]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1029.825 4.2375 1029.96 4.3725 ;
      END
   END din0[316]
   PIN din0[317]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1032.685 4.2375 1032.82 4.3725 ;
      END
   END din0[317]
   PIN din0[318]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1035.545 4.2375 1035.68 4.3725 ;
      END
   END din0[318]
   PIN din0[319]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1038.405 4.2375 1038.54 4.3725 ;
      END
   END din0[319]
   PIN din0[320]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1041.265 4.2375 1041.4 4.3725 ;
      END
   END din0[320]
   PIN din0[321]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1044.125 4.2375 1044.26 4.3725 ;
      END
   END din0[321]
   PIN din0[322]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1046.985 4.2375 1047.12 4.3725 ;
      END
   END din0[322]
   PIN din0[323]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1049.845 4.2375 1049.98 4.3725 ;
      END
   END din0[323]
   PIN din0[324]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1052.705 4.2375 1052.84 4.3725 ;
      END
   END din0[324]
   PIN din0[325]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1055.565 4.2375 1055.7 4.3725 ;
      END
   END din0[325]
   PIN din0[326]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1058.425 4.2375 1058.56 4.3725 ;
      END
   END din0[326]
   PIN din0[327]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1061.285 4.2375 1061.42 4.3725 ;
      END
   END din0[327]
   PIN din0[328]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1064.145 4.2375 1064.28 4.3725 ;
      END
   END din0[328]
   PIN din0[329]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1067.005 4.2375 1067.14 4.3725 ;
      END
   END din0[329]
   PIN din0[330]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1069.865 4.2375 1070.0 4.3725 ;
      END
   END din0[330]
   PIN din0[331]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1072.725 4.2375 1072.86 4.3725 ;
      END
   END din0[331]
   PIN din0[332]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1075.585 4.2375 1075.72 4.3725 ;
      END
   END din0[332]
   PIN din0[333]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1078.445 4.2375 1078.58 4.3725 ;
      END
   END din0[333]
   PIN din0[334]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1081.305 4.2375 1081.44 4.3725 ;
      END
   END din0[334]
   PIN din0[335]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1084.165 4.2375 1084.3 4.3725 ;
      END
   END din0[335]
   PIN din0[336]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1087.025 4.2375 1087.16 4.3725 ;
      END
   END din0[336]
   PIN din0[337]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1089.885 4.2375 1090.02 4.3725 ;
      END
   END din0[337]
   PIN din0[338]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1092.745 4.2375 1092.88 4.3725 ;
      END
   END din0[338]
   PIN din0[339]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1095.605 4.2375 1095.74 4.3725 ;
      END
   END din0[339]
   PIN din0[340]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1098.465 4.2375 1098.6 4.3725 ;
      END
   END din0[340]
   PIN din0[341]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1101.325 4.2375 1101.46 4.3725 ;
      END
   END din0[341]
   PIN din0[342]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1104.185 4.2375 1104.32 4.3725 ;
      END
   END din0[342]
   PIN din0[343]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1107.045 4.2375 1107.18 4.3725 ;
      END
   END din0[343]
   PIN din0[344]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1109.905 4.2375 1110.04 4.3725 ;
      END
   END din0[344]
   PIN din0[345]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1112.765 4.2375 1112.9 4.3725 ;
      END
   END din0[345]
   PIN din0[346]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1115.625 4.2375 1115.76 4.3725 ;
      END
   END din0[346]
   PIN din0[347]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1118.485 4.2375 1118.62 4.3725 ;
      END
   END din0[347]
   PIN din0[348]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1121.345 4.2375 1121.48 4.3725 ;
      END
   END din0[348]
   PIN din0[349]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1124.205 4.2375 1124.34 4.3725 ;
      END
   END din0[349]
   PIN din0[350]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1127.065 4.2375 1127.2 4.3725 ;
      END
   END din0[350]
   PIN din0[351]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1129.925 4.2375 1130.06 4.3725 ;
      END
   END din0[351]
   PIN din0[352]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1132.785 4.2375 1132.92 4.3725 ;
      END
   END din0[352]
   PIN din0[353]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1135.645 4.2375 1135.78 4.3725 ;
      END
   END din0[353]
   PIN din0[354]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1138.505 4.2375 1138.64 4.3725 ;
      END
   END din0[354]
   PIN din0[355]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1141.365 4.2375 1141.5 4.3725 ;
      END
   END din0[355]
   PIN din0[356]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1144.225 4.2375 1144.36 4.3725 ;
      END
   END din0[356]
   PIN din0[357]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1147.085 4.2375 1147.22 4.3725 ;
      END
   END din0[357]
   PIN din0[358]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1149.945 4.2375 1150.08 4.3725 ;
      END
   END din0[358]
   PIN din0[359]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1152.805 4.2375 1152.94 4.3725 ;
      END
   END din0[359]
   PIN din0[360]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1155.665 4.2375 1155.8 4.3725 ;
      END
   END din0[360]
   PIN din0[361]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1158.525 4.2375 1158.66 4.3725 ;
      END
   END din0[361]
   PIN din0[362]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1161.385 4.2375 1161.52 4.3725 ;
      END
   END din0[362]
   PIN din0[363]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1164.245 4.2375 1164.38 4.3725 ;
      END
   END din0[363]
   PIN din0[364]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1167.105 4.2375 1167.24 4.3725 ;
      END
   END din0[364]
   PIN din0[365]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1169.965 4.2375 1170.1 4.3725 ;
      END
   END din0[365]
   PIN din0[366]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1172.825 4.2375 1172.96 4.3725 ;
      END
   END din0[366]
   PIN din0[367]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1175.685 4.2375 1175.82 4.3725 ;
      END
   END din0[367]
   PIN din0[368]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1178.545 4.2375 1178.68 4.3725 ;
      END
   END din0[368]
   PIN din0[369]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1181.405 4.2375 1181.54 4.3725 ;
      END
   END din0[369]
   PIN din0[370]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1184.265 4.2375 1184.4 4.3725 ;
      END
   END din0[370]
   PIN din0[371]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1187.125 4.2375 1187.26 4.3725 ;
      END
   END din0[371]
   PIN din0[372]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1189.985 4.2375 1190.12 4.3725 ;
      END
   END din0[372]
   PIN din0[373]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1192.845 4.2375 1192.98 4.3725 ;
      END
   END din0[373]
   PIN din0[374]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1195.705 4.2375 1195.84 4.3725 ;
      END
   END din0[374]
   PIN din0[375]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1198.565 4.2375 1198.7 4.3725 ;
      END
   END din0[375]
   PIN din0[376]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1201.425 4.2375 1201.56 4.3725 ;
      END
   END din0[376]
   PIN din0[377]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1204.285 4.2375 1204.42 4.3725 ;
      END
   END din0[377]
   PIN din0[378]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1207.145 4.2375 1207.28 4.3725 ;
      END
   END din0[378]
   PIN din0[379]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1210.005 4.2375 1210.14 4.3725 ;
      END
   END din0[379]
   PIN din0[380]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1212.865 4.2375 1213.0 4.3725 ;
      END
   END din0[380]
   PIN din0[381]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1215.725 4.2375 1215.86 4.3725 ;
      END
   END din0[381]
   PIN din0[382]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1218.585 4.2375 1218.72 4.3725 ;
      END
   END din0[382]
   PIN din0[383]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1221.445 4.2375 1221.58 4.3725 ;
      END
   END din0[383]
   PIN din0[384]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1224.305 4.2375 1224.44 4.3725 ;
      END
   END din0[384]
   PIN din0[385]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1227.165 4.2375 1227.3 4.3725 ;
      END
   END din0[385]
   PIN din0[386]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1230.025 4.2375 1230.16 4.3725 ;
      END
   END din0[386]
   PIN din0[387]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1232.885 4.2375 1233.02 4.3725 ;
      END
   END din0[387]
   PIN din0[388]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1235.745 4.2375 1235.88 4.3725 ;
      END
   END din0[388]
   PIN din0[389]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1238.605 4.2375 1238.74 4.3725 ;
      END
   END din0[389]
   PIN din0[390]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1241.465 4.2375 1241.6 4.3725 ;
      END
   END din0[390]
   PIN din0[391]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1244.325 4.2375 1244.46 4.3725 ;
      END
   END din0[391]
   PIN din0[392]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1247.185 4.2375 1247.32 4.3725 ;
      END
   END din0[392]
   PIN din0[393]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1250.045 4.2375 1250.18 4.3725 ;
      END
   END din0[393]
   PIN din0[394]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1252.905 4.2375 1253.04 4.3725 ;
      END
   END din0[394]
   PIN din0[395]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1255.765 4.2375 1255.9 4.3725 ;
      END
   END din0[395]
   PIN din0[396]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1258.625 4.2375 1258.76 4.3725 ;
      END
   END din0[396]
   PIN din0[397]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1261.485 4.2375 1261.62 4.3725 ;
      END
   END din0[397]
   PIN din0[398]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1264.345 4.2375 1264.48 4.3725 ;
      END
   END din0[398]
   PIN din0[399]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1267.205 4.2375 1267.34 4.3725 ;
      END
   END din0[399]
   PIN din0[400]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1270.065 4.2375 1270.2 4.3725 ;
      END
   END din0[400]
   PIN din0[401]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1272.925 4.2375 1273.06 4.3725 ;
      END
   END din0[401]
   PIN din0[402]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1275.785 4.2375 1275.92 4.3725 ;
      END
   END din0[402]
   PIN din0[403]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1278.645 4.2375 1278.78 4.3725 ;
      END
   END din0[403]
   PIN din0[404]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1281.505 4.2375 1281.64 4.3725 ;
      END
   END din0[404]
   PIN din0[405]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1284.365 4.2375 1284.5 4.3725 ;
      END
   END din0[405]
   PIN din0[406]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1287.225 4.2375 1287.36 4.3725 ;
      END
   END din0[406]
   PIN din0[407]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1290.085 4.2375 1290.22 4.3725 ;
      END
   END din0[407]
   PIN din0[408]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1292.945 4.2375 1293.08 4.3725 ;
      END
   END din0[408]
   PIN din0[409]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1295.805 4.2375 1295.94 4.3725 ;
      END
   END din0[409]
   PIN din0[410]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1298.665 4.2375 1298.8 4.3725 ;
      END
   END din0[410]
   PIN din0[411]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1301.525 4.2375 1301.66 4.3725 ;
      END
   END din0[411]
   PIN din0[412]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1304.385 4.2375 1304.52 4.3725 ;
      END
   END din0[412]
   PIN din0[413]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1307.245 4.2375 1307.38 4.3725 ;
      END
   END din0[413]
   PIN din0[414]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1310.105 4.2375 1310.24 4.3725 ;
      END
   END din0[414]
   PIN din0[415]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1312.965 4.2375 1313.1 4.3725 ;
      END
   END din0[415]
   PIN din0[416]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1315.825 4.2375 1315.96 4.3725 ;
      END
   END din0[416]
   PIN din0[417]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1318.685 4.2375 1318.82 4.3725 ;
      END
   END din0[417]
   PIN din0[418]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1321.545 4.2375 1321.68 4.3725 ;
      END
   END din0[418]
   PIN din0[419]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1324.405 4.2375 1324.54 4.3725 ;
      END
   END din0[419]
   PIN din0[420]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1327.265 4.2375 1327.4 4.3725 ;
      END
   END din0[420]
   PIN din0[421]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1330.125 4.2375 1330.26 4.3725 ;
      END
   END din0[421]
   PIN din0[422]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1332.985 4.2375 1333.12 4.3725 ;
      END
   END din0[422]
   PIN din0[423]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1335.845 4.2375 1335.98 4.3725 ;
      END
   END din0[423]
   PIN din0[424]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1338.705 4.2375 1338.84 4.3725 ;
      END
   END din0[424]
   PIN din0[425]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1341.565 4.2375 1341.7 4.3725 ;
      END
   END din0[425]
   PIN din0[426]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1344.425 4.2375 1344.56 4.3725 ;
      END
   END din0[426]
   PIN din0[427]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1347.285 4.2375 1347.42 4.3725 ;
      END
   END din0[427]
   PIN din0[428]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1350.145 4.2375 1350.28 4.3725 ;
      END
   END din0[428]
   PIN din0[429]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1353.005 4.2375 1353.14 4.3725 ;
      END
   END din0[429]
   PIN din0[430]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1355.865 4.2375 1356.0 4.3725 ;
      END
   END din0[430]
   PIN din0[431]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1358.725 4.2375 1358.86 4.3725 ;
      END
   END din0[431]
   PIN din0[432]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1361.585 4.2375 1361.72 4.3725 ;
      END
   END din0[432]
   PIN din0[433]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1364.445 4.2375 1364.58 4.3725 ;
      END
   END din0[433]
   PIN din0[434]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1367.305 4.2375 1367.44 4.3725 ;
      END
   END din0[434]
   PIN din0[435]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1370.165 4.2375 1370.3 4.3725 ;
      END
   END din0[435]
   PIN din0[436]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1373.025 4.2375 1373.16 4.3725 ;
      END
   END din0[436]
   PIN din0[437]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1375.885 4.2375 1376.02 4.3725 ;
      END
   END din0[437]
   PIN din0[438]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1378.745 4.2375 1378.88 4.3725 ;
      END
   END din0[438]
   PIN din0[439]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1381.605 4.2375 1381.74 4.3725 ;
      END
   END din0[439]
   PIN din0[440]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1384.465 4.2375 1384.6 4.3725 ;
      END
   END din0[440]
   PIN din0[441]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1387.325 4.2375 1387.46 4.3725 ;
      END
   END din0[441]
   PIN din0[442]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1390.185 4.2375 1390.32 4.3725 ;
      END
   END din0[442]
   PIN din0[443]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1393.045 4.2375 1393.18 4.3725 ;
      END
   END din0[443]
   PIN din0[444]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1395.905 4.2375 1396.04 4.3725 ;
      END
   END din0[444]
   PIN din0[445]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1398.765 4.2375 1398.9 4.3725 ;
      END
   END din0[445]
   PIN din0[446]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1401.625 4.2375 1401.76 4.3725 ;
      END
   END din0[446]
   PIN din0[447]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1404.485 4.2375 1404.62 4.3725 ;
      END
   END din0[447]
   PIN din0[448]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1407.345 4.2375 1407.48 4.3725 ;
      END
   END din0[448]
   PIN din0[449]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1410.205 4.2375 1410.34 4.3725 ;
      END
   END din0[449]
   PIN din0[450]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1413.065 4.2375 1413.2 4.3725 ;
      END
   END din0[450]
   PIN din0[451]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1415.925 4.2375 1416.06 4.3725 ;
      END
   END din0[451]
   PIN din0[452]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1418.785 4.2375 1418.92 4.3725 ;
      END
   END din0[452]
   PIN din0[453]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1421.645 4.2375 1421.78 4.3725 ;
      END
   END din0[453]
   PIN din0[454]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1424.505 4.2375 1424.64 4.3725 ;
      END
   END din0[454]
   PIN din0[455]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1427.365 4.2375 1427.5 4.3725 ;
      END
   END din0[455]
   PIN din0[456]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1430.225 4.2375 1430.36 4.3725 ;
      END
   END din0[456]
   PIN din0[457]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1433.085 4.2375 1433.22 4.3725 ;
      END
   END din0[457]
   PIN din0[458]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1435.945 4.2375 1436.08 4.3725 ;
      END
   END din0[458]
   PIN din0[459]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1438.805 4.2375 1438.94 4.3725 ;
      END
   END din0[459]
   PIN din0[460]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1441.665 4.2375 1441.8 4.3725 ;
      END
   END din0[460]
   PIN din0[461]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1444.525 4.2375 1444.66 4.3725 ;
      END
   END din0[461]
   PIN din0[462]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1447.385 4.2375 1447.52 4.3725 ;
      END
   END din0[462]
   PIN din0[463]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1450.245 4.2375 1450.38 4.3725 ;
      END
   END din0[463]
   PIN din0[464]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1453.105 4.2375 1453.24 4.3725 ;
      END
   END din0[464]
   PIN din0[465]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1455.965 4.2375 1456.1 4.3725 ;
      END
   END din0[465]
   PIN din0[466]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1458.825 4.2375 1458.96 4.3725 ;
      END
   END din0[466]
   PIN din0[467]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1461.685 4.2375 1461.82 4.3725 ;
      END
   END din0[467]
   PIN din0[468]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1464.545 4.2375 1464.68 4.3725 ;
      END
   END din0[468]
   PIN din0[469]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1467.405 4.2375 1467.54 4.3725 ;
      END
   END din0[469]
   PIN din0[470]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1470.265 4.2375 1470.4 4.3725 ;
      END
   END din0[470]
   PIN din0[471]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1473.125 4.2375 1473.26 4.3725 ;
      END
   END din0[471]
   PIN din0[472]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1475.985 4.2375 1476.12 4.3725 ;
      END
   END din0[472]
   PIN din0[473]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1478.845 4.2375 1478.98 4.3725 ;
      END
   END din0[473]
   PIN din0[474]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1481.705 4.2375 1481.84 4.3725 ;
      END
   END din0[474]
   PIN din0[475]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1484.565 4.2375 1484.7 4.3725 ;
      END
   END din0[475]
   PIN din0[476]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1487.425 4.2375 1487.56 4.3725 ;
      END
   END din0[476]
   PIN din0[477]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1490.285 4.2375 1490.42 4.3725 ;
      END
   END din0[477]
   PIN din0[478]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1493.145 4.2375 1493.28 4.3725 ;
      END
   END din0[478]
   PIN din0[479]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1496.005 4.2375 1496.14 4.3725 ;
      END
   END din0[479]
   PIN din0[480]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1498.865 4.2375 1499.0 4.3725 ;
      END
   END din0[480]
   PIN din0[481]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1501.725 4.2375 1501.86 4.3725 ;
      END
   END din0[481]
   PIN din0[482]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1504.585 4.2375 1504.72 4.3725 ;
      END
   END din0[482]
   PIN din0[483]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1507.445 4.2375 1507.58 4.3725 ;
      END
   END din0[483]
   PIN din0[484]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1510.305 4.2375 1510.44 4.3725 ;
      END
   END din0[484]
   PIN din0[485]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1513.165 4.2375 1513.3 4.3725 ;
      END
   END din0[485]
   PIN din0[486]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1516.025 4.2375 1516.16 4.3725 ;
      END
   END din0[486]
   PIN din0[487]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1518.885 4.2375 1519.02 4.3725 ;
      END
   END din0[487]
   PIN din0[488]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1521.745 4.2375 1521.88 4.3725 ;
      END
   END din0[488]
   PIN din0[489]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1524.605 4.2375 1524.74 4.3725 ;
      END
   END din0[489]
   PIN din0[490]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1527.465 4.2375 1527.6 4.3725 ;
      END
   END din0[490]
   PIN din0[491]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1530.325 4.2375 1530.46 4.3725 ;
      END
   END din0[491]
   PIN din0[492]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1533.185 4.2375 1533.32 4.3725 ;
      END
   END din0[492]
   PIN din0[493]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1536.045 4.2375 1536.18 4.3725 ;
      END
   END din0[493]
   PIN din0[494]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1538.905 4.2375 1539.04 4.3725 ;
      END
   END din0[494]
   PIN din0[495]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1541.765 4.2375 1541.9 4.3725 ;
      END
   END din0[495]
   PIN din0[496]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1544.625 4.2375 1544.76 4.3725 ;
      END
   END din0[496]
   PIN din0[497]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1547.485 4.2375 1547.62 4.3725 ;
      END
   END din0[497]
   PIN din0[498]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1550.345 4.2375 1550.48 4.3725 ;
      END
   END din0[498]
   PIN din0[499]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1553.205 4.2375 1553.34 4.3725 ;
      END
   END din0[499]
   PIN din0[500]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1556.065 4.2375 1556.2 4.3725 ;
      END
   END din0[500]
   PIN din0[501]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1558.925 4.2375 1559.06 4.3725 ;
      END
   END din0[501]
   PIN din0[502]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1561.785 4.2375 1561.92 4.3725 ;
      END
   END din0[502]
   PIN din0[503]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1564.645 4.2375 1564.78 4.3725 ;
      END
   END din0[503]
   PIN din0[504]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1567.505 4.2375 1567.64 4.3725 ;
      END
   END din0[504]
   PIN din0[505]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1570.365 4.2375 1570.5 4.3725 ;
      END
   END din0[505]
   PIN din0[506]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1573.225 4.2375 1573.36 4.3725 ;
      END
   END din0[506]
   PIN din0[507]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1576.085 4.2375 1576.22 4.3725 ;
      END
   END din0[507]
   PIN din0[508]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1578.945 4.2375 1579.08 4.3725 ;
      END
   END din0[508]
   PIN din0[509]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1581.805 4.2375 1581.94 4.3725 ;
      END
   END din0[509]
   PIN din0[510]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1584.665 4.2375 1584.8 4.3725 ;
      END
   END din0[510]
   PIN din0[511]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1587.525 4.2375 1587.66 4.3725 ;
      END
   END din0[511]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.345 122.4325 120.48 122.5675 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.345 125.1625 120.48 125.2975 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.345 127.3725 120.48 127.5075 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.345 130.1025 120.48 130.2375 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.345 132.3125 120.48 132.4475 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.345 135.0425 120.48 135.1775 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.225 96.3025 801.36 96.4375 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.225 93.5725 801.36 93.7075 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.225 91.3625 801.36 91.4975 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.225 88.6325 801.36 88.7675 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.225 86.4225 801.36 86.5575 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.225 83.6925 801.36 83.8275 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  3.385 77.8425 3.52 77.9775 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  918.325 210.0025 918.46 210.1375 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.3475 77.9275 9.4825 78.0625 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  912.2225 209.9175 912.3575 210.0525 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.9225 203.295 160.0575 203.43 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.0975 203.295 161.2325 203.43 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.2725 203.295 162.4075 203.43 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.4475 203.295 163.5825 203.43 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.6225 203.295 164.7575 203.43 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.7975 203.295 165.9325 203.43 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.9725 203.295 167.1075 203.43 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.1475 203.295 168.2825 203.43 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.3225 203.295 169.4575 203.43 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.4975 203.295 170.6325 203.43 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.6725 203.295 171.8075 203.43 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.8475 203.295 172.9825 203.43 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.0225 203.295 174.1575 203.43 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.1975 203.295 175.3325 203.43 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.3725 203.295 176.5075 203.43 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.5475 203.295 177.6825 203.43 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.7225 203.295 178.8575 203.43 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.8975 203.295 180.0325 203.43 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.0725 203.295 181.2075 203.43 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.2475 203.295 182.3825 203.43 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.4225 203.295 183.5575 203.43 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.5975 203.295 184.7325 203.43 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.7725 203.295 185.9075 203.43 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.9475 203.295 187.0825 203.43 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.1225 203.295 188.2575 203.43 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.2975 203.295 189.4325 203.43 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.4725 203.295 190.6075 203.43 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.6475 203.295 191.7825 203.43 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.8225 203.295 192.9575 203.43 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.9975 203.295 194.1325 203.43 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.1725 203.295 195.3075 203.43 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.3475 203.295 196.4825 203.43 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.5225 203.295 197.6575 203.43 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.6975 203.295 198.8325 203.43 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.8725 203.295 200.0075 203.43 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.0475 203.295 201.1825 203.43 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.2225 203.295 202.3575 203.43 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.3975 203.295 203.5325 203.43 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.5725 203.295 204.7075 203.43 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.7475 203.295 205.8825 203.43 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.9225 203.295 207.0575 203.43 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.0975 203.295 208.2325 203.43 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.2725 203.295 209.4075 203.43 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.4475 203.295 210.5825 203.43 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.6225 203.295 211.7575 203.43 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.7975 203.295 212.9325 203.43 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.9725 203.295 214.1075 203.43 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.1475 203.295 215.2825 203.43 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.3225 203.295 216.4575 203.43 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.4975 203.295 217.6325 203.43 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.6725 203.295 218.8075 203.43 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.8475 203.295 219.9825 203.43 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.0225 203.295 221.1575 203.43 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.1975 203.295 222.3325 203.43 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.3725 203.295 223.5075 203.43 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.5475 203.295 224.6825 203.43 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.7225 203.295 225.8575 203.43 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.8975 203.295 227.0325 203.43 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.0725 203.295 228.2075 203.43 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.2475 203.295 229.3825 203.43 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.4225 203.295 230.5575 203.43 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.5975 203.295 231.7325 203.43 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.7725 203.295 232.9075 203.43 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.9475 203.295 234.0825 203.43 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.1225 203.295 235.2575 203.43 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.2975 203.295 236.4325 203.43 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.4725 203.295 237.6075 203.43 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.6475 203.295 238.7825 203.43 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.8225 203.295 239.9575 203.43 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.9975 203.295 241.1325 203.43 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.1725 203.295 242.3075 203.43 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.3475 203.295 243.4825 203.43 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.5225 203.295 244.6575 203.43 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.6975 203.295 245.8325 203.43 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.8725 203.295 247.0075 203.43 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.0475 203.295 248.1825 203.43 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.2225 203.295 249.3575 203.43 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.3975 203.295 250.5325 203.43 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.5725 203.295 251.7075 203.43 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.7475 203.295 252.8825 203.43 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.9225 203.295 254.0575 203.43 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.0975 203.295 255.2325 203.43 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.2725 203.295 256.4075 203.43 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.4475 203.295 257.5825 203.43 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.6225 203.295 258.7575 203.43 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.7975 203.295 259.9325 203.43 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.9725 203.295 261.1075 203.43 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.1475 203.295 262.2825 203.43 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.3225 203.295 263.4575 203.43 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.4975 203.295 264.6325 203.43 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.6725 203.295 265.8075 203.43 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.8475 203.295 266.9825 203.43 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.0225 203.295 268.1575 203.43 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.1975 203.295 269.3325 203.43 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.3725 203.295 270.5075 203.43 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.5475 203.295 271.6825 203.43 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.7225 203.295 272.8575 203.43 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.8975 203.295 274.0325 203.43 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.0725 203.295 275.2075 203.43 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.2475 203.295 276.3825 203.43 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.4225 203.295 277.5575 203.43 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.5975 203.295 278.7325 203.43 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.7725 203.295 279.9075 203.43 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.9475 203.295 281.0825 203.43 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  282.1225 203.295 282.2575 203.43 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.2975 203.295 283.4325 203.43 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.4725 203.295 284.6075 203.43 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.6475 203.295 285.7825 203.43 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.8225 203.295 286.9575 203.43 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.9975 203.295 288.1325 203.43 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.1725 203.295 289.3075 203.43 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.3475 203.295 290.4825 203.43 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.5225 203.295 291.6575 203.43 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.6975 203.295 292.8325 203.43 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.8725 203.295 294.0075 203.43 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.0475 203.295 295.1825 203.43 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.2225 203.295 296.3575 203.43 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.3975 203.295 297.5325 203.43 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.5725 203.295 298.7075 203.43 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.7475 203.295 299.8825 203.43 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.9225 203.295 301.0575 203.43 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  302.0975 203.295 302.2325 203.43 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.2725 203.295 303.4075 203.43 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.4475 203.295 304.5825 203.43 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.6225 203.295 305.7575 203.43 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.7975 203.295 306.9325 203.43 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.9725 203.295 308.1075 203.43 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.1475 203.295 309.2825 203.43 ;
      END
   END dout1[127]
   PIN dout1[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.3225 203.295 310.4575 203.43 ;
      END
   END dout1[128]
   PIN dout1[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.4975 203.295 311.6325 203.43 ;
      END
   END dout1[129]
   PIN dout1[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.6725 203.295 312.8075 203.43 ;
      END
   END dout1[130]
   PIN dout1[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.8475 203.295 313.9825 203.43 ;
      END
   END dout1[131]
   PIN dout1[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.0225 203.295 315.1575 203.43 ;
      END
   END dout1[132]
   PIN dout1[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.1975 203.295 316.3325 203.43 ;
      END
   END dout1[133]
   PIN dout1[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.3725 203.295 317.5075 203.43 ;
      END
   END dout1[134]
   PIN dout1[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.5475 203.295 318.6825 203.43 ;
      END
   END dout1[135]
   PIN dout1[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.7225 203.295 319.8575 203.43 ;
      END
   END dout1[136]
   PIN dout1[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.8975 203.295 321.0325 203.43 ;
      END
   END dout1[137]
   PIN dout1[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  322.0725 203.295 322.2075 203.43 ;
      END
   END dout1[138]
   PIN dout1[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.2475 203.295 323.3825 203.43 ;
      END
   END dout1[139]
   PIN dout1[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.4225 203.295 324.5575 203.43 ;
      END
   END dout1[140]
   PIN dout1[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.5975 203.295 325.7325 203.43 ;
      END
   END dout1[141]
   PIN dout1[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.7725 203.295 326.9075 203.43 ;
      END
   END dout1[142]
   PIN dout1[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.9475 203.295 328.0825 203.43 ;
      END
   END dout1[143]
   PIN dout1[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.1225 203.295 329.2575 203.43 ;
      END
   END dout1[144]
   PIN dout1[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.2975 203.295 330.4325 203.43 ;
      END
   END dout1[145]
   PIN dout1[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.4725 203.295 331.6075 203.43 ;
      END
   END dout1[146]
   PIN dout1[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.6475 203.295 332.7825 203.43 ;
      END
   END dout1[147]
   PIN dout1[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.8225 203.295 333.9575 203.43 ;
      END
   END dout1[148]
   PIN dout1[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.9975 203.295 335.1325 203.43 ;
      END
   END dout1[149]
   PIN dout1[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.1725 203.295 336.3075 203.43 ;
      END
   END dout1[150]
   PIN dout1[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.3475 203.295 337.4825 203.43 ;
      END
   END dout1[151]
   PIN dout1[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.5225 203.295 338.6575 203.43 ;
      END
   END dout1[152]
   PIN dout1[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.6975 203.295 339.8325 203.43 ;
      END
   END dout1[153]
   PIN dout1[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.8725 203.295 341.0075 203.43 ;
      END
   END dout1[154]
   PIN dout1[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.0475 203.295 342.1825 203.43 ;
      END
   END dout1[155]
   PIN dout1[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.2225 203.295 343.3575 203.43 ;
      END
   END dout1[156]
   PIN dout1[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.3975 203.295 344.5325 203.43 ;
      END
   END dout1[157]
   PIN dout1[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.5725 203.295 345.7075 203.43 ;
      END
   END dout1[158]
   PIN dout1[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.7475 203.295 346.8825 203.43 ;
      END
   END dout1[159]
   PIN dout1[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.9225 203.295 348.0575 203.43 ;
      END
   END dout1[160]
   PIN dout1[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.0975 203.295 349.2325 203.43 ;
      END
   END dout1[161]
   PIN dout1[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.2725 203.295 350.4075 203.43 ;
      END
   END dout1[162]
   PIN dout1[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  351.4475 203.295 351.5825 203.43 ;
      END
   END dout1[163]
   PIN dout1[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.6225 203.295 352.7575 203.43 ;
      END
   END dout1[164]
   PIN dout1[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.7975 203.295 353.9325 203.43 ;
      END
   END dout1[165]
   PIN dout1[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.9725 203.295 355.1075 203.43 ;
      END
   END dout1[166]
   PIN dout1[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.1475 203.295 356.2825 203.43 ;
      END
   END dout1[167]
   PIN dout1[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.3225 203.295 357.4575 203.43 ;
      END
   END dout1[168]
   PIN dout1[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.4975 203.295 358.6325 203.43 ;
      END
   END dout1[169]
   PIN dout1[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.6725 203.295 359.8075 203.43 ;
      END
   END dout1[170]
   PIN dout1[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.8475 203.295 360.9825 203.43 ;
      END
   END dout1[171]
   PIN dout1[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.0225 203.295 362.1575 203.43 ;
      END
   END dout1[172]
   PIN dout1[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.1975 203.295 363.3325 203.43 ;
      END
   END dout1[173]
   PIN dout1[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.3725 203.295 364.5075 203.43 ;
      END
   END dout1[174]
   PIN dout1[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.5475 203.295 365.6825 203.43 ;
      END
   END dout1[175]
   PIN dout1[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.7225 203.295 366.8575 203.43 ;
      END
   END dout1[176]
   PIN dout1[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.8975 203.295 368.0325 203.43 ;
      END
   END dout1[177]
   PIN dout1[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.0725 203.295 369.2075 203.43 ;
      END
   END dout1[178]
   PIN dout1[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.2475 203.295 370.3825 203.43 ;
      END
   END dout1[179]
   PIN dout1[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  371.4225 203.295 371.5575 203.43 ;
      END
   END dout1[180]
   PIN dout1[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.5975 203.295 372.7325 203.43 ;
      END
   END dout1[181]
   PIN dout1[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.7725 203.295 373.9075 203.43 ;
      END
   END dout1[182]
   PIN dout1[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.9475 203.295 375.0825 203.43 ;
      END
   END dout1[183]
   PIN dout1[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  376.1225 203.295 376.2575 203.43 ;
      END
   END dout1[184]
   PIN dout1[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.2975 203.295 377.4325 203.43 ;
      END
   END dout1[185]
   PIN dout1[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.4725 203.295 378.6075 203.43 ;
      END
   END dout1[186]
   PIN dout1[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  379.6475 203.295 379.7825 203.43 ;
      END
   END dout1[187]
   PIN dout1[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.8225 203.295 380.9575 203.43 ;
      END
   END dout1[188]
   PIN dout1[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.9975 203.295 382.1325 203.43 ;
      END
   END dout1[189]
   PIN dout1[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.1725 203.295 383.3075 203.43 ;
      END
   END dout1[190]
   PIN dout1[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.3475 203.295 384.4825 203.43 ;
      END
   END dout1[191]
   PIN dout1[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  385.5225 203.295 385.6575 203.43 ;
      END
   END dout1[192]
   PIN dout1[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.6975 203.295 386.8325 203.43 ;
      END
   END dout1[193]
   PIN dout1[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  387.8725 203.295 388.0075 203.43 ;
      END
   END dout1[194]
   PIN dout1[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.0475 203.295 389.1825 203.43 ;
      END
   END dout1[195]
   PIN dout1[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  390.2225 203.295 390.3575 203.43 ;
      END
   END dout1[196]
   PIN dout1[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  391.3975 203.295 391.5325 203.43 ;
      END
   END dout1[197]
   PIN dout1[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.5725 203.295 392.7075 203.43 ;
      END
   END dout1[198]
   PIN dout1[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.7475 203.295 393.8825 203.43 ;
      END
   END dout1[199]
   PIN dout1[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.9225 203.295 395.0575 203.43 ;
      END
   END dout1[200]
   PIN dout1[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.0975 203.295 396.2325 203.43 ;
      END
   END dout1[201]
   PIN dout1[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.2725 203.295 397.4075 203.43 ;
      END
   END dout1[202]
   PIN dout1[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.4475 203.295 398.5825 203.43 ;
      END
   END dout1[203]
   PIN dout1[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.6225 203.295 399.7575 203.43 ;
      END
   END dout1[204]
   PIN dout1[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.7975 203.295 400.9325 203.43 ;
      END
   END dout1[205]
   PIN dout1[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.9725 203.295 402.1075 203.43 ;
      END
   END dout1[206]
   PIN dout1[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.1475 203.295 403.2825 203.43 ;
      END
   END dout1[207]
   PIN dout1[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.3225 203.295 404.4575 203.43 ;
      END
   END dout1[208]
   PIN dout1[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  405.4975 203.295 405.6325 203.43 ;
      END
   END dout1[209]
   PIN dout1[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.6725 203.295 406.8075 203.43 ;
      END
   END dout1[210]
   PIN dout1[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.8475 203.295 407.9825 203.43 ;
      END
   END dout1[211]
   PIN dout1[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.0225 203.295 409.1575 203.43 ;
      END
   END dout1[212]
   PIN dout1[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.1975 203.295 410.3325 203.43 ;
      END
   END dout1[213]
   PIN dout1[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  411.3725 203.295 411.5075 203.43 ;
      END
   END dout1[214]
   PIN dout1[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.5475 203.295 412.6825 203.43 ;
      END
   END dout1[215]
   PIN dout1[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  413.7225 203.295 413.8575 203.43 ;
      END
   END dout1[216]
   PIN dout1[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  414.8975 203.295 415.0325 203.43 ;
      END
   END dout1[217]
   PIN dout1[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  416.0725 203.295 416.2075 203.43 ;
      END
   END dout1[218]
   PIN dout1[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.2475 203.295 417.3825 203.43 ;
      END
   END dout1[219]
   PIN dout1[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.4225 203.295 418.5575 203.43 ;
      END
   END dout1[220]
   PIN dout1[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  419.5975 203.295 419.7325 203.43 ;
      END
   END dout1[221]
   PIN dout1[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.7725 203.295 420.9075 203.43 ;
      END
   END dout1[222]
   PIN dout1[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.9475 203.295 422.0825 203.43 ;
      END
   END dout1[223]
   PIN dout1[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.1225 203.295 423.2575 203.43 ;
      END
   END dout1[224]
   PIN dout1[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.2975 203.295 424.4325 203.43 ;
      END
   END dout1[225]
   PIN dout1[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  425.4725 203.295 425.6075 203.43 ;
      END
   END dout1[226]
   PIN dout1[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.6475 203.295 426.7825 203.43 ;
      END
   END dout1[227]
   PIN dout1[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.8225 203.295 427.9575 203.43 ;
      END
   END dout1[228]
   PIN dout1[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  428.9975 203.295 429.1325 203.43 ;
      END
   END dout1[229]
   PIN dout1[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  430.1725 203.295 430.3075 203.43 ;
      END
   END dout1[230]
   PIN dout1[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  431.3475 203.295 431.4825 203.43 ;
      END
   END dout1[231]
   PIN dout1[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.5225 203.295 432.6575 203.43 ;
      END
   END dout1[232]
   PIN dout1[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  433.6975 203.295 433.8325 203.43 ;
      END
   END dout1[233]
   PIN dout1[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  434.8725 203.295 435.0075 203.43 ;
      END
   END dout1[234]
   PIN dout1[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  436.0475 203.295 436.1825 203.43 ;
      END
   END dout1[235]
   PIN dout1[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  437.2225 203.295 437.3575 203.43 ;
      END
   END dout1[236]
   PIN dout1[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.3975 203.295 438.5325 203.43 ;
      END
   END dout1[237]
   PIN dout1[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  439.5725 203.295 439.7075 203.43 ;
      END
   END dout1[238]
   PIN dout1[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.7475 203.295 440.8825 203.43 ;
      END
   END dout1[239]
   PIN dout1[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.9225 203.295 442.0575 203.43 ;
      END
   END dout1[240]
   PIN dout1[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.0975 203.295 443.2325 203.43 ;
      END
   END dout1[241]
   PIN dout1[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.2725 203.295 444.4075 203.43 ;
      END
   END dout1[242]
   PIN dout1[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  445.4475 203.295 445.5825 203.43 ;
      END
   END dout1[243]
   PIN dout1[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.6225 203.295 446.7575 203.43 ;
      END
   END dout1[244]
   PIN dout1[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.7975 203.295 447.9325 203.43 ;
      END
   END dout1[245]
   PIN dout1[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  448.9725 203.295 449.1075 203.43 ;
      END
   END dout1[246]
   PIN dout1[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  450.1475 203.295 450.2825 203.43 ;
      END
   END dout1[247]
   PIN dout1[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  451.3225 203.295 451.4575 203.43 ;
      END
   END dout1[248]
   PIN dout1[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.4975 203.295 452.6325 203.43 ;
      END
   END dout1[249]
   PIN dout1[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.6725 203.295 453.8075 203.43 ;
      END
   END dout1[250]
   PIN dout1[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  454.8475 203.295 454.9825 203.43 ;
      END
   END dout1[251]
   PIN dout1[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  456.0225 203.295 456.1575 203.43 ;
      END
   END dout1[252]
   PIN dout1[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  457.1975 203.295 457.3325 203.43 ;
      END
   END dout1[253]
   PIN dout1[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.3725 203.295 458.5075 203.43 ;
      END
   END dout1[254]
   PIN dout1[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  459.5475 203.295 459.6825 203.43 ;
      END
   END dout1[255]
   PIN dout1[256]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  460.7225 203.295 460.8575 203.43 ;
      END
   END dout1[256]
   PIN dout1[257]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.8975 203.295 462.0325 203.43 ;
      END
   END dout1[257]
   PIN dout1[258]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  463.0725 203.295 463.2075 203.43 ;
      END
   END dout1[258]
   PIN dout1[259]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.2475 203.295 464.3825 203.43 ;
      END
   END dout1[259]
   PIN dout1[260]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  465.4225 203.295 465.5575 203.43 ;
      END
   END dout1[260]
   PIN dout1[261]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.5975 203.295 466.7325 203.43 ;
      END
   END dout1[261]
   PIN dout1[262]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.7725 203.295 467.9075 203.43 ;
      END
   END dout1[262]
   PIN dout1[263]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  468.9475 203.295 469.0825 203.43 ;
      END
   END dout1[263]
   PIN dout1[264]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.1225 203.295 470.2575 203.43 ;
      END
   END dout1[264]
   PIN dout1[265]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  471.2975 203.295 471.4325 203.43 ;
      END
   END dout1[265]
   PIN dout1[266]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.4725 203.295 472.6075 203.43 ;
      END
   END dout1[266]
   PIN dout1[267]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  473.6475 203.295 473.7825 203.43 ;
      END
   END dout1[267]
   PIN dout1[268]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  474.8225 203.295 474.9575 203.43 ;
      END
   END dout1[268]
   PIN dout1[269]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.9975 203.295 476.1325 203.43 ;
      END
   END dout1[269]
   PIN dout1[270]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  477.1725 203.295 477.3075 203.43 ;
      END
   END dout1[270]
   PIN dout1[271]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.3475 203.295 478.4825 203.43 ;
      END
   END dout1[271]
   PIN dout1[272]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  479.5225 203.295 479.6575 203.43 ;
      END
   END dout1[272]
   PIN dout1[273]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  480.6975 203.295 480.8325 203.43 ;
      END
   END dout1[273]
   PIN dout1[274]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.8725 203.295 482.0075 203.43 ;
      END
   END dout1[274]
   PIN dout1[275]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  483.0475 203.295 483.1825 203.43 ;
      END
   END dout1[275]
   PIN dout1[276]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.2225 203.295 484.3575 203.43 ;
      END
   END dout1[276]
   PIN dout1[277]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  485.3975 203.295 485.5325 203.43 ;
      END
   END dout1[277]
   PIN dout1[278]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.5725 203.295 486.7075 203.43 ;
      END
   END dout1[278]
   PIN dout1[279]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.7475 203.295 487.8825 203.43 ;
      END
   END dout1[279]
   PIN dout1[280]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  488.9225 203.295 489.0575 203.43 ;
      END
   END dout1[280]
   PIN dout1[281]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  490.0975 203.295 490.2325 203.43 ;
      END
   END dout1[281]
   PIN dout1[282]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  491.2725 203.295 491.4075 203.43 ;
      END
   END dout1[282]
   PIN dout1[283]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.4475 203.295 492.5825 203.43 ;
      END
   END dout1[283]
   PIN dout1[284]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  493.6225 203.295 493.7575 203.43 ;
      END
   END dout1[284]
   PIN dout1[285]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  494.7975 203.295 494.9325 203.43 ;
      END
   END dout1[285]
   PIN dout1[286]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.9725 203.295 496.1075 203.43 ;
      END
   END dout1[286]
   PIN dout1[287]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  497.1475 203.295 497.2825 203.43 ;
      END
   END dout1[287]
   PIN dout1[288]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.3225 203.295 498.4575 203.43 ;
      END
   END dout1[288]
   PIN dout1[289]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  499.4975 203.295 499.6325 203.43 ;
      END
   END dout1[289]
   PIN dout1[290]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  500.6725 203.295 500.8075 203.43 ;
      END
   END dout1[290]
   PIN dout1[291]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.8475 203.295 501.9825 203.43 ;
      END
   END dout1[291]
   PIN dout1[292]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  503.0225 203.295 503.1575 203.43 ;
      END
   END dout1[292]
   PIN dout1[293]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.1975 203.295 504.3325 203.43 ;
      END
   END dout1[293]
   PIN dout1[294]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  505.3725 203.295 505.5075 203.43 ;
      END
   END dout1[294]
   PIN dout1[295]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  506.5475 203.295 506.6825 203.43 ;
      END
   END dout1[295]
   PIN dout1[296]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.7225 203.295 507.8575 203.43 ;
      END
   END dout1[296]
   PIN dout1[297]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  508.8975 203.295 509.0325 203.43 ;
      END
   END dout1[297]
   PIN dout1[298]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.0725 203.295 510.2075 203.43 ;
      END
   END dout1[298]
   PIN dout1[299]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  511.2475 203.295 511.3825 203.43 ;
      END
   END dout1[299]
   PIN dout1[300]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.4225 203.295 512.5575 203.43 ;
      END
   END dout1[300]
   PIN dout1[301]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  513.5975 203.295 513.7325 203.43 ;
      END
   END dout1[301]
   PIN dout1[302]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.7725 203.295 514.9075 203.43 ;
      END
   END dout1[302]
   PIN dout1[303]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.9475 203.295 516.0825 203.43 ;
      END
   END dout1[303]
   PIN dout1[304]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  517.1225 203.295 517.2575 203.43 ;
      END
   END dout1[304]
   PIN dout1[305]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.2975 203.295 518.4325 203.43 ;
      END
   END dout1[305]
   PIN dout1[306]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  519.4725 203.295 519.6075 203.43 ;
      END
   END dout1[306]
   PIN dout1[307]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  520.6475 203.295 520.7825 203.43 ;
      END
   END dout1[307]
   PIN dout1[308]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.8225 203.295 521.9575 203.43 ;
      END
   END dout1[308]
   PIN dout1[309]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  522.9975 203.295 523.1325 203.43 ;
      END
   END dout1[309]
   PIN dout1[310]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  524.1725 203.295 524.3075 203.43 ;
      END
   END dout1[310]
   PIN dout1[311]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  525.3475 203.295 525.4825 203.43 ;
      END
   END dout1[311]
   PIN dout1[312]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  526.5225 203.295 526.6575 203.43 ;
      END
   END dout1[312]
   PIN dout1[313]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.6975 203.295 527.8325 203.43 ;
      END
   END dout1[313]
   PIN dout1[314]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  528.8725 203.295 529.0075 203.43 ;
      END
   END dout1[314]
   PIN dout1[315]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  530.0475 203.295 530.1825 203.43 ;
      END
   END dout1[315]
   PIN dout1[316]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  531.2225 203.295 531.3575 203.43 ;
      END
   END dout1[316]
   PIN dout1[317]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  532.3975 203.295 532.5325 203.43 ;
      END
   END dout1[317]
   PIN dout1[318]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  533.5725 203.295 533.7075 203.43 ;
      END
   END dout1[318]
   PIN dout1[319]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  534.7475 203.295 534.8825 203.43 ;
      END
   END dout1[319]
   PIN dout1[320]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  535.9225 203.295 536.0575 203.43 ;
      END
   END dout1[320]
   PIN dout1[321]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  537.0975 203.295 537.2325 203.43 ;
      END
   END dout1[321]
   PIN dout1[322]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  538.2725 203.295 538.4075 203.43 ;
      END
   END dout1[322]
   PIN dout1[323]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  539.4475 203.295 539.5825 203.43 ;
      END
   END dout1[323]
   PIN dout1[324]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  540.6225 203.295 540.7575 203.43 ;
      END
   END dout1[324]
   PIN dout1[325]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  541.7975 203.295 541.9325 203.43 ;
      END
   END dout1[325]
   PIN dout1[326]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  542.9725 203.295 543.1075 203.43 ;
      END
   END dout1[326]
   PIN dout1[327]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  544.1475 203.295 544.2825 203.43 ;
      END
   END dout1[327]
   PIN dout1[328]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  545.3225 203.295 545.4575 203.43 ;
      END
   END dout1[328]
   PIN dout1[329]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  546.4975 203.295 546.6325 203.43 ;
      END
   END dout1[329]
   PIN dout1[330]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  547.6725 203.295 547.8075 203.43 ;
      END
   END dout1[330]
   PIN dout1[331]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  548.8475 203.295 548.9825 203.43 ;
      END
   END dout1[331]
   PIN dout1[332]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  550.0225 203.295 550.1575 203.43 ;
      END
   END dout1[332]
   PIN dout1[333]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  551.1975 203.295 551.3325 203.43 ;
      END
   END dout1[333]
   PIN dout1[334]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  552.3725 203.295 552.5075 203.43 ;
      END
   END dout1[334]
   PIN dout1[335]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  553.5475 203.295 553.6825 203.43 ;
      END
   END dout1[335]
   PIN dout1[336]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  554.7225 203.295 554.8575 203.43 ;
      END
   END dout1[336]
   PIN dout1[337]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  555.8975 203.295 556.0325 203.43 ;
      END
   END dout1[337]
   PIN dout1[338]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  557.0725 203.295 557.2075 203.43 ;
      END
   END dout1[338]
   PIN dout1[339]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  558.2475 203.295 558.3825 203.43 ;
      END
   END dout1[339]
   PIN dout1[340]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  559.4225 203.295 559.5575 203.43 ;
      END
   END dout1[340]
   PIN dout1[341]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  560.5975 203.295 560.7325 203.43 ;
      END
   END dout1[341]
   PIN dout1[342]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  561.7725 203.295 561.9075 203.43 ;
      END
   END dout1[342]
   PIN dout1[343]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  562.9475 203.295 563.0825 203.43 ;
      END
   END dout1[343]
   PIN dout1[344]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  564.1225 203.295 564.2575 203.43 ;
      END
   END dout1[344]
   PIN dout1[345]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  565.2975 203.295 565.4325 203.43 ;
      END
   END dout1[345]
   PIN dout1[346]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  566.4725 203.295 566.6075 203.43 ;
      END
   END dout1[346]
   PIN dout1[347]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  567.6475 203.295 567.7825 203.43 ;
      END
   END dout1[347]
   PIN dout1[348]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  568.8225 203.295 568.9575 203.43 ;
      END
   END dout1[348]
   PIN dout1[349]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  569.9975 203.295 570.1325 203.43 ;
      END
   END dout1[349]
   PIN dout1[350]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  571.1725 203.295 571.3075 203.43 ;
      END
   END dout1[350]
   PIN dout1[351]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  572.3475 203.295 572.4825 203.43 ;
      END
   END dout1[351]
   PIN dout1[352]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  573.5225 203.295 573.6575 203.43 ;
      END
   END dout1[352]
   PIN dout1[353]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  574.6975 203.295 574.8325 203.43 ;
      END
   END dout1[353]
   PIN dout1[354]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  575.8725 203.295 576.0075 203.43 ;
      END
   END dout1[354]
   PIN dout1[355]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  577.0475 203.295 577.1825 203.43 ;
      END
   END dout1[355]
   PIN dout1[356]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  578.2225 203.295 578.3575 203.43 ;
      END
   END dout1[356]
   PIN dout1[357]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  579.3975 203.295 579.5325 203.43 ;
      END
   END dout1[357]
   PIN dout1[358]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  580.5725 203.295 580.7075 203.43 ;
      END
   END dout1[358]
   PIN dout1[359]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  581.7475 203.295 581.8825 203.43 ;
      END
   END dout1[359]
   PIN dout1[360]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  582.9225 203.295 583.0575 203.43 ;
      END
   END dout1[360]
   PIN dout1[361]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  584.0975 203.295 584.2325 203.43 ;
      END
   END dout1[361]
   PIN dout1[362]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  585.2725 203.295 585.4075 203.43 ;
      END
   END dout1[362]
   PIN dout1[363]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  586.4475 203.295 586.5825 203.43 ;
      END
   END dout1[363]
   PIN dout1[364]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  587.6225 203.295 587.7575 203.43 ;
      END
   END dout1[364]
   PIN dout1[365]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  588.7975 203.295 588.9325 203.43 ;
      END
   END dout1[365]
   PIN dout1[366]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  589.9725 203.295 590.1075 203.43 ;
      END
   END dout1[366]
   PIN dout1[367]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  591.1475 203.295 591.2825 203.43 ;
      END
   END dout1[367]
   PIN dout1[368]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  592.3225 203.295 592.4575 203.43 ;
      END
   END dout1[368]
   PIN dout1[369]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  593.4975 203.295 593.6325 203.43 ;
      END
   END dout1[369]
   PIN dout1[370]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  594.6725 203.295 594.8075 203.43 ;
      END
   END dout1[370]
   PIN dout1[371]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  595.8475 203.295 595.9825 203.43 ;
      END
   END dout1[371]
   PIN dout1[372]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  597.0225 203.295 597.1575 203.43 ;
      END
   END dout1[372]
   PIN dout1[373]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  598.1975 203.295 598.3325 203.43 ;
      END
   END dout1[373]
   PIN dout1[374]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  599.3725 203.295 599.5075 203.43 ;
      END
   END dout1[374]
   PIN dout1[375]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  600.5475 203.295 600.6825 203.43 ;
      END
   END dout1[375]
   PIN dout1[376]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  601.7225 203.295 601.8575 203.43 ;
      END
   END dout1[376]
   PIN dout1[377]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  602.8975 203.295 603.0325 203.43 ;
      END
   END dout1[377]
   PIN dout1[378]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  604.0725 203.295 604.2075 203.43 ;
      END
   END dout1[378]
   PIN dout1[379]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  605.2475 203.295 605.3825 203.43 ;
      END
   END dout1[379]
   PIN dout1[380]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  606.4225 203.295 606.5575 203.43 ;
      END
   END dout1[380]
   PIN dout1[381]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  607.5975 203.295 607.7325 203.43 ;
      END
   END dout1[381]
   PIN dout1[382]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  608.7725 203.295 608.9075 203.43 ;
      END
   END dout1[382]
   PIN dout1[383]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  609.9475 203.295 610.0825 203.43 ;
      END
   END dout1[383]
   PIN dout1[384]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  611.1225 203.295 611.2575 203.43 ;
      END
   END dout1[384]
   PIN dout1[385]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  612.2975 203.295 612.4325 203.43 ;
      END
   END dout1[385]
   PIN dout1[386]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  613.4725 203.295 613.6075 203.43 ;
      END
   END dout1[386]
   PIN dout1[387]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  614.6475 203.295 614.7825 203.43 ;
      END
   END dout1[387]
   PIN dout1[388]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  615.8225 203.295 615.9575 203.43 ;
      END
   END dout1[388]
   PIN dout1[389]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  616.9975 203.295 617.1325 203.43 ;
      END
   END dout1[389]
   PIN dout1[390]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  618.1725 203.295 618.3075 203.43 ;
      END
   END dout1[390]
   PIN dout1[391]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  619.3475 203.295 619.4825 203.43 ;
      END
   END dout1[391]
   PIN dout1[392]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  620.5225 203.295 620.6575 203.43 ;
      END
   END dout1[392]
   PIN dout1[393]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  621.6975 203.295 621.8325 203.43 ;
      END
   END dout1[393]
   PIN dout1[394]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  622.8725 203.295 623.0075 203.43 ;
      END
   END dout1[394]
   PIN dout1[395]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  624.0475 203.295 624.1825 203.43 ;
      END
   END dout1[395]
   PIN dout1[396]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  625.2225 203.295 625.3575 203.43 ;
      END
   END dout1[396]
   PIN dout1[397]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  626.3975 203.295 626.5325 203.43 ;
      END
   END dout1[397]
   PIN dout1[398]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  627.5725 203.295 627.7075 203.43 ;
      END
   END dout1[398]
   PIN dout1[399]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  628.7475 203.295 628.8825 203.43 ;
      END
   END dout1[399]
   PIN dout1[400]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  629.9225 203.295 630.0575 203.43 ;
      END
   END dout1[400]
   PIN dout1[401]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  631.0975 203.295 631.2325 203.43 ;
      END
   END dout1[401]
   PIN dout1[402]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  632.2725 203.295 632.4075 203.43 ;
      END
   END dout1[402]
   PIN dout1[403]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  633.4475 203.295 633.5825 203.43 ;
      END
   END dout1[403]
   PIN dout1[404]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  634.6225 203.295 634.7575 203.43 ;
      END
   END dout1[404]
   PIN dout1[405]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  635.7975 203.295 635.9325 203.43 ;
      END
   END dout1[405]
   PIN dout1[406]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  636.9725 203.295 637.1075 203.43 ;
      END
   END dout1[406]
   PIN dout1[407]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  638.1475 203.295 638.2825 203.43 ;
      END
   END dout1[407]
   PIN dout1[408]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  639.3225 203.295 639.4575 203.43 ;
      END
   END dout1[408]
   PIN dout1[409]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  640.4975 203.295 640.6325 203.43 ;
      END
   END dout1[409]
   PIN dout1[410]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  641.6725 203.295 641.8075 203.43 ;
      END
   END dout1[410]
   PIN dout1[411]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  642.8475 203.295 642.9825 203.43 ;
      END
   END dout1[411]
   PIN dout1[412]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  644.0225 203.295 644.1575 203.43 ;
      END
   END dout1[412]
   PIN dout1[413]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  645.1975 203.295 645.3325 203.43 ;
      END
   END dout1[413]
   PIN dout1[414]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  646.3725 203.295 646.5075 203.43 ;
      END
   END dout1[414]
   PIN dout1[415]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  647.5475 203.295 647.6825 203.43 ;
      END
   END dout1[415]
   PIN dout1[416]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  648.7225 203.295 648.8575 203.43 ;
      END
   END dout1[416]
   PIN dout1[417]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  649.8975 203.295 650.0325 203.43 ;
      END
   END dout1[417]
   PIN dout1[418]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  651.0725 203.295 651.2075 203.43 ;
      END
   END dout1[418]
   PIN dout1[419]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  652.2475 203.295 652.3825 203.43 ;
      END
   END dout1[419]
   PIN dout1[420]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  653.4225 203.295 653.5575 203.43 ;
      END
   END dout1[420]
   PIN dout1[421]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  654.5975 203.295 654.7325 203.43 ;
      END
   END dout1[421]
   PIN dout1[422]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  655.7725 203.295 655.9075 203.43 ;
      END
   END dout1[422]
   PIN dout1[423]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  656.9475 203.295 657.0825 203.43 ;
      END
   END dout1[423]
   PIN dout1[424]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  658.1225 203.295 658.2575 203.43 ;
      END
   END dout1[424]
   PIN dout1[425]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  659.2975 203.295 659.4325 203.43 ;
      END
   END dout1[425]
   PIN dout1[426]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  660.4725 203.295 660.6075 203.43 ;
      END
   END dout1[426]
   PIN dout1[427]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  661.6475 203.295 661.7825 203.43 ;
      END
   END dout1[427]
   PIN dout1[428]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  662.8225 203.295 662.9575 203.43 ;
      END
   END dout1[428]
   PIN dout1[429]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  663.9975 203.295 664.1325 203.43 ;
      END
   END dout1[429]
   PIN dout1[430]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  665.1725 203.295 665.3075 203.43 ;
      END
   END dout1[430]
   PIN dout1[431]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  666.3475 203.295 666.4825 203.43 ;
      END
   END dout1[431]
   PIN dout1[432]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  667.5225 203.295 667.6575 203.43 ;
      END
   END dout1[432]
   PIN dout1[433]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  668.6975 203.295 668.8325 203.43 ;
      END
   END dout1[433]
   PIN dout1[434]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  669.8725 203.295 670.0075 203.43 ;
      END
   END dout1[434]
   PIN dout1[435]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  671.0475 203.295 671.1825 203.43 ;
      END
   END dout1[435]
   PIN dout1[436]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  672.2225 203.295 672.3575 203.43 ;
      END
   END dout1[436]
   PIN dout1[437]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  673.3975 203.295 673.5325 203.43 ;
      END
   END dout1[437]
   PIN dout1[438]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  674.5725 203.295 674.7075 203.43 ;
      END
   END dout1[438]
   PIN dout1[439]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  675.7475 203.295 675.8825 203.43 ;
      END
   END dout1[439]
   PIN dout1[440]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  676.9225 203.295 677.0575 203.43 ;
      END
   END dout1[440]
   PIN dout1[441]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  678.0975 203.295 678.2325 203.43 ;
      END
   END dout1[441]
   PIN dout1[442]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  679.2725 203.295 679.4075 203.43 ;
      END
   END dout1[442]
   PIN dout1[443]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  680.4475 203.295 680.5825 203.43 ;
      END
   END dout1[443]
   PIN dout1[444]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  681.6225 203.295 681.7575 203.43 ;
      END
   END dout1[444]
   PIN dout1[445]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  682.7975 203.295 682.9325 203.43 ;
      END
   END dout1[445]
   PIN dout1[446]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  683.9725 203.295 684.1075 203.43 ;
      END
   END dout1[446]
   PIN dout1[447]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  685.1475 203.295 685.2825 203.43 ;
      END
   END dout1[447]
   PIN dout1[448]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  686.3225 203.295 686.4575 203.43 ;
      END
   END dout1[448]
   PIN dout1[449]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  687.4975 203.295 687.6325 203.43 ;
      END
   END dout1[449]
   PIN dout1[450]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  688.6725 203.295 688.8075 203.43 ;
      END
   END dout1[450]
   PIN dout1[451]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  689.8475 203.295 689.9825 203.43 ;
      END
   END dout1[451]
   PIN dout1[452]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  691.0225 203.295 691.1575 203.43 ;
      END
   END dout1[452]
   PIN dout1[453]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  692.1975 203.295 692.3325 203.43 ;
      END
   END dout1[453]
   PIN dout1[454]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  693.3725 203.295 693.5075 203.43 ;
      END
   END dout1[454]
   PIN dout1[455]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  694.5475 203.295 694.6825 203.43 ;
      END
   END dout1[455]
   PIN dout1[456]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  695.7225 203.295 695.8575 203.43 ;
      END
   END dout1[456]
   PIN dout1[457]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  696.8975 203.295 697.0325 203.43 ;
      END
   END dout1[457]
   PIN dout1[458]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  698.0725 203.295 698.2075 203.43 ;
      END
   END dout1[458]
   PIN dout1[459]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  699.2475 203.295 699.3825 203.43 ;
      END
   END dout1[459]
   PIN dout1[460]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  700.4225 203.295 700.5575 203.43 ;
      END
   END dout1[460]
   PIN dout1[461]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  701.5975 203.295 701.7325 203.43 ;
      END
   END dout1[461]
   PIN dout1[462]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  702.7725 203.295 702.9075 203.43 ;
      END
   END dout1[462]
   PIN dout1[463]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  703.9475 203.295 704.0825 203.43 ;
      END
   END dout1[463]
   PIN dout1[464]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  705.1225 203.295 705.2575 203.43 ;
      END
   END dout1[464]
   PIN dout1[465]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  706.2975 203.295 706.4325 203.43 ;
      END
   END dout1[465]
   PIN dout1[466]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  707.4725 203.295 707.6075 203.43 ;
      END
   END dout1[466]
   PIN dout1[467]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  708.6475 203.295 708.7825 203.43 ;
      END
   END dout1[467]
   PIN dout1[468]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  709.8225 203.295 709.9575 203.43 ;
      END
   END dout1[468]
   PIN dout1[469]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  710.9975 203.295 711.1325 203.43 ;
      END
   END dout1[469]
   PIN dout1[470]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  712.1725 203.295 712.3075 203.43 ;
      END
   END dout1[470]
   PIN dout1[471]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  713.3475 203.295 713.4825 203.43 ;
      END
   END dout1[471]
   PIN dout1[472]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  714.5225 203.295 714.6575 203.43 ;
      END
   END dout1[472]
   PIN dout1[473]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  715.6975 203.295 715.8325 203.43 ;
      END
   END dout1[473]
   PIN dout1[474]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  716.8725 203.295 717.0075 203.43 ;
      END
   END dout1[474]
   PIN dout1[475]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  718.0475 203.295 718.1825 203.43 ;
      END
   END dout1[475]
   PIN dout1[476]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  719.2225 203.295 719.3575 203.43 ;
      END
   END dout1[476]
   PIN dout1[477]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  720.3975 203.295 720.5325 203.43 ;
      END
   END dout1[477]
   PIN dout1[478]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  721.5725 203.295 721.7075 203.43 ;
      END
   END dout1[478]
   PIN dout1[479]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  722.7475 203.295 722.8825 203.43 ;
      END
   END dout1[479]
   PIN dout1[480]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  723.9225 203.295 724.0575 203.43 ;
      END
   END dout1[480]
   PIN dout1[481]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  725.0975 203.295 725.2325 203.43 ;
      END
   END dout1[481]
   PIN dout1[482]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  726.2725 203.295 726.4075 203.43 ;
      END
   END dout1[482]
   PIN dout1[483]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  727.4475 203.295 727.5825 203.43 ;
      END
   END dout1[483]
   PIN dout1[484]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  728.6225 203.295 728.7575 203.43 ;
      END
   END dout1[484]
   PIN dout1[485]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  729.7975 203.295 729.9325 203.43 ;
      END
   END dout1[485]
   PIN dout1[486]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  730.9725 203.295 731.1075 203.43 ;
      END
   END dout1[486]
   PIN dout1[487]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  732.1475 203.295 732.2825 203.43 ;
      END
   END dout1[487]
   PIN dout1[488]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  733.3225 203.295 733.4575 203.43 ;
      END
   END dout1[488]
   PIN dout1[489]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  734.4975 203.295 734.6325 203.43 ;
      END
   END dout1[489]
   PIN dout1[490]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  735.6725 203.295 735.8075 203.43 ;
      END
   END dout1[490]
   PIN dout1[491]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  736.8475 203.295 736.9825 203.43 ;
      END
   END dout1[491]
   PIN dout1[492]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  738.0225 203.295 738.1575 203.43 ;
      END
   END dout1[492]
   PIN dout1[493]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  739.1975 203.295 739.3325 203.43 ;
      END
   END dout1[493]
   PIN dout1[494]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  740.3725 203.295 740.5075 203.43 ;
      END
   END dout1[494]
   PIN dout1[495]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  741.5475 203.295 741.6825 203.43 ;
      END
   END dout1[495]
   PIN dout1[496]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  742.7225 203.295 742.8575 203.43 ;
      END
   END dout1[496]
   PIN dout1[497]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  743.8975 203.295 744.0325 203.43 ;
      END
   END dout1[497]
   PIN dout1[498]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  745.0725 203.295 745.2075 203.43 ;
      END
   END dout1[498]
   PIN dout1[499]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  746.2475 203.295 746.3825 203.43 ;
      END
   END dout1[499]
   PIN dout1[500]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  747.4225 203.295 747.5575 203.43 ;
      END
   END dout1[500]
   PIN dout1[501]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  748.5975 203.295 748.7325 203.43 ;
      END
   END dout1[501]
   PIN dout1[502]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  749.7725 203.295 749.9075 203.43 ;
      END
   END dout1[502]
   PIN dout1[503]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  750.9475 203.295 751.0825 203.43 ;
      END
   END dout1[503]
   PIN dout1[504]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  752.1225 203.295 752.2575 203.43 ;
      END
   END dout1[504]
   PIN dout1[505]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  753.2975 203.295 753.4325 203.43 ;
      END
   END dout1[505]
   PIN dout1[506]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  754.4725 203.295 754.6075 203.43 ;
      END
   END dout1[506]
   PIN dout1[507]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  755.6475 203.295 755.7825 203.43 ;
      END
   END dout1[507]
   PIN dout1[508]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  756.8225 203.295 756.9575 203.43 ;
      END
   END dout1[508]
   PIN dout1[509]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  757.9975 203.295 758.1325 203.43 ;
      END
   END dout1[509]
   PIN dout1[510]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  759.1725 203.295 759.3075 203.43 ;
      END
   END dout1[510]
   PIN dout1[511]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  760.3475 203.295 760.4825 203.43 ;
      END
   END dout1[511]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  1.4 1.4 1591.94 2.1 ;
         LAYER metal3 ;
         RECT  1.4 212.24 1591.94 212.94 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 212.94 ;
         LAYER metal4 ;
         RECT  1591.24 1.4 1591.94 212.94 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  1592.64 0.0 1593.34 214.34 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 214.34 ;
         LAYER metal3 ;
         RECT  0.0 0.0 1593.34 0.7 ;
         LAYER metal3 ;
         RECT  0.0 213.64 1593.34 214.34 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 1593.2 214.2 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 1593.2 214.2 ;
   LAYER  metal3 ;
      RECT  0.14 4.0975 125.925 4.5125 ;
      RECT  126.34 4.0975 128.785 4.5125 ;
      RECT  129.2 4.0975 131.645 4.5125 ;
      RECT  132.06 4.0975 134.505 4.5125 ;
      RECT  134.92 4.0975 137.365 4.5125 ;
      RECT  137.78 4.0975 140.225 4.5125 ;
      RECT  140.64 4.0975 143.085 4.5125 ;
      RECT  143.5 4.0975 145.945 4.5125 ;
      RECT  146.36 4.0975 148.805 4.5125 ;
      RECT  149.22 4.0975 151.665 4.5125 ;
      RECT  152.08 4.0975 154.525 4.5125 ;
      RECT  154.94 4.0975 157.385 4.5125 ;
      RECT  157.8 4.0975 160.245 4.5125 ;
      RECT  160.66 4.0975 163.105 4.5125 ;
      RECT  163.52 4.0975 165.965 4.5125 ;
      RECT  166.38 4.0975 168.825 4.5125 ;
      RECT  169.24 4.0975 171.685 4.5125 ;
      RECT  172.1 4.0975 174.545 4.5125 ;
      RECT  174.96 4.0975 177.405 4.5125 ;
      RECT  177.82 4.0975 180.265 4.5125 ;
      RECT  180.68 4.0975 183.125 4.5125 ;
      RECT  183.54 4.0975 185.985 4.5125 ;
      RECT  186.4 4.0975 188.845 4.5125 ;
      RECT  189.26 4.0975 191.705 4.5125 ;
      RECT  192.12 4.0975 194.565 4.5125 ;
      RECT  194.98 4.0975 197.425 4.5125 ;
      RECT  197.84 4.0975 200.285 4.5125 ;
      RECT  200.7 4.0975 203.145 4.5125 ;
      RECT  203.56 4.0975 206.005 4.5125 ;
      RECT  206.42 4.0975 208.865 4.5125 ;
      RECT  209.28 4.0975 211.725 4.5125 ;
      RECT  212.14 4.0975 214.585 4.5125 ;
      RECT  215.0 4.0975 217.445 4.5125 ;
      RECT  217.86 4.0975 220.305 4.5125 ;
      RECT  220.72 4.0975 223.165 4.5125 ;
      RECT  223.58 4.0975 226.025 4.5125 ;
      RECT  226.44 4.0975 228.885 4.5125 ;
      RECT  229.3 4.0975 231.745 4.5125 ;
      RECT  232.16 4.0975 234.605 4.5125 ;
      RECT  235.02 4.0975 237.465 4.5125 ;
      RECT  237.88 4.0975 240.325 4.5125 ;
      RECT  240.74 4.0975 243.185 4.5125 ;
      RECT  243.6 4.0975 246.045 4.5125 ;
      RECT  246.46 4.0975 248.905 4.5125 ;
      RECT  249.32 4.0975 251.765 4.5125 ;
      RECT  252.18 4.0975 254.625 4.5125 ;
      RECT  255.04 4.0975 257.485 4.5125 ;
      RECT  257.9 4.0975 260.345 4.5125 ;
      RECT  260.76 4.0975 263.205 4.5125 ;
      RECT  263.62 4.0975 266.065 4.5125 ;
      RECT  266.48 4.0975 268.925 4.5125 ;
      RECT  269.34 4.0975 271.785 4.5125 ;
      RECT  272.2 4.0975 274.645 4.5125 ;
      RECT  275.06 4.0975 277.505 4.5125 ;
      RECT  277.92 4.0975 280.365 4.5125 ;
      RECT  280.78 4.0975 283.225 4.5125 ;
      RECT  283.64 4.0975 286.085 4.5125 ;
      RECT  286.5 4.0975 288.945 4.5125 ;
      RECT  289.36 4.0975 291.805 4.5125 ;
      RECT  292.22 4.0975 294.665 4.5125 ;
      RECT  295.08 4.0975 297.525 4.5125 ;
      RECT  297.94 4.0975 300.385 4.5125 ;
      RECT  300.8 4.0975 303.245 4.5125 ;
      RECT  303.66 4.0975 306.105 4.5125 ;
      RECT  306.52 4.0975 308.965 4.5125 ;
      RECT  309.38 4.0975 311.825 4.5125 ;
      RECT  312.24 4.0975 314.685 4.5125 ;
      RECT  315.1 4.0975 317.545 4.5125 ;
      RECT  317.96 4.0975 320.405 4.5125 ;
      RECT  320.82 4.0975 323.265 4.5125 ;
      RECT  323.68 4.0975 326.125 4.5125 ;
      RECT  326.54 4.0975 328.985 4.5125 ;
      RECT  329.4 4.0975 331.845 4.5125 ;
      RECT  332.26 4.0975 334.705 4.5125 ;
      RECT  335.12 4.0975 337.565 4.5125 ;
      RECT  337.98 4.0975 340.425 4.5125 ;
      RECT  340.84 4.0975 343.285 4.5125 ;
      RECT  343.7 4.0975 346.145 4.5125 ;
      RECT  346.56 4.0975 349.005 4.5125 ;
      RECT  349.42 4.0975 351.865 4.5125 ;
      RECT  352.28 4.0975 354.725 4.5125 ;
      RECT  355.14 4.0975 357.585 4.5125 ;
      RECT  358.0 4.0975 360.445 4.5125 ;
      RECT  360.86 4.0975 363.305 4.5125 ;
      RECT  363.72 4.0975 366.165 4.5125 ;
      RECT  366.58 4.0975 369.025 4.5125 ;
      RECT  369.44 4.0975 371.885 4.5125 ;
      RECT  372.3 4.0975 374.745 4.5125 ;
      RECT  375.16 4.0975 377.605 4.5125 ;
      RECT  378.02 4.0975 380.465 4.5125 ;
      RECT  380.88 4.0975 383.325 4.5125 ;
      RECT  383.74 4.0975 386.185 4.5125 ;
      RECT  386.6 4.0975 389.045 4.5125 ;
      RECT  389.46 4.0975 391.905 4.5125 ;
      RECT  392.32 4.0975 394.765 4.5125 ;
      RECT  395.18 4.0975 397.625 4.5125 ;
      RECT  398.04 4.0975 400.485 4.5125 ;
      RECT  400.9 4.0975 403.345 4.5125 ;
      RECT  403.76 4.0975 406.205 4.5125 ;
      RECT  406.62 4.0975 409.065 4.5125 ;
      RECT  409.48 4.0975 411.925 4.5125 ;
      RECT  412.34 4.0975 414.785 4.5125 ;
      RECT  415.2 4.0975 417.645 4.5125 ;
      RECT  418.06 4.0975 420.505 4.5125 ;
      RECT  420.92 4.0975 423.365 4.5125 ;
      RECT  423.78 4.0975 426.225 4.5125 ;
      RECT  426.64 4.0975 429.085 4.5125 ;
      RECT  429.5 4.0975 431.945 4.5125 ;
      RECT  432.36 4.0975 434.805 4.5125 ;
      RECT  435.22 4.0975 437.665 4.5125 ;
      RECT  438.08 4.0975 440.525 4.5125 ;
      RECT  440.94 4.0975 443.385 4.5125 ;
      RECT  443.8 4.0975 446.245 4.5125 ;
      RECT  446.66 4.0975 449.105 4.5125 ;
      RECT  449.52 4.0975 451.965 4.5125 ;
      RECT  452.38 4.0975 454.825 4.5125 ;
      RECT  455.24 4.0975 457.685 4.5125 ;
      RECT  458.1 4.0975 460.545 4.5125 ;
      RECT  460.96 4.0975 463.405 4.5125 ;
      RECT  463.82 4.0975 466.265 4.5125 ;
      RECT  466.68 4.0975 469.125 4.5125 ;
      RECT  469.54 4.0975 471.985 4.5125 ;
      RECT  472.4 4.0975 474.845 4.5125 ;
      RECT  475.26 4.0975 477.705 4.5125 ;
      RECT  478.12 4.0975 480.565 4.5125 ;
      RECT  480.98 4.0975 483.425 4.5125 ;
      RECT  483.84 4.0975 486.285 4.5125 ;
      RECT  486.7 4.0975 489.145 4.5125 ;
      RECT  489.56 4.0975 492.005 4.5125 ;
      RECT  492.42 4.0975 494.865 4.5125 ;
      RECT  495.28 4.0975 497.725 4.5125 ;
      RECT  498.14 4.0975 500.585 4.5125 ;
      RECT  501.0 4.0975 503.445 4.5125 ;
      RECT  503.86 4.0975 506.305 4.5125 ;
      RECT  506.72 4.0975 509.165 4.5125 ;
      RECT  509.58 4.0975 512.025 4.5125 ;
      RECT  512.44 4.0975 514.885 4.5125 ;
      RECT  515.3 4.0975 517.745 4.5125 ;
      RECT  518.16 4.0975 520.605 4.5125 ;
      RECT  521.02 4.0975 523.465 4.5125 ;
      RECT  523.88 4.0975 526.325 4.5125 ;
      RECT  526.74 4.0975 529.185 4.5125 ;
      RECT  529.6 4.0975 532.045 4.5125 ;
      RECT  532.46 4.0975 534.905 4.5125 ;
      RECT  535.32 4.0975 537.765 4.5125 ;
      RECT  538.18 4.0975 540.625 4.5125 ;
      RECT  541.04 4.0975 543.485 4.5125 ;
      RECT  543.9 4.0975 546.345 4.5125 ;
      RECT  546.76 4.0975 549.205 4.5125 ;
      RECT  549.62 4.0975 552.065 4.5125 ;
      RECT  552.48 4.0975 554.925 4.5125 ;
      RECT  555.34 4.0975 557.785 4.5125 ;
      RECT  558.2 4.0975 560.645 4.5125 ;
      RECT  561.06 4.0975 563.505 4.5125 ;
      RECT  563.92 4.0975 566.365 4.5125 ;
      RECT  566.78 4.0975 569.225 4.5125 ;
      RECT  569.64 4.0975 572.085 4.5125 ;
      RECT  572.5 4.0975 574.945 4.5125 ;
      RECT  575.36 4.0975 577.805 4.5125 ;
      RECT  578.22 4.0975 580.665 4.5125 ;
      RECT  581.08 4.0975 583.525 4.5125 ;
      RECT  583.94 4.0975 586.385 4.5125 ;
      RECT  586.8 4.0975 589.245 4.5125 ;
      RECT  589.66 4.0975 592.105 4.5125 ;
      RECT  592.52 4.0975 594.965 4.5125 ;
      RECT  595.38 4.0975 597.825 4.5125 ;
      RECT  598.24 4.0975 600.685 4.5125 ;
      RECT  601.1 4.0975 603.545 4.5125 ;
      RECT  603.96 4.0975 606.405 4.5125 ;
      RECT  606.82 4.0975 609.265 4.5125 ;
      RECT  609.68 4.0975 612.125 4.5125 ;
      RECT  612.54 4.0975 614.985 4.5125 ;
      RECT  615.4 4.0975 617.845 4.5125 ;
      RECT  618.26 4.0975 620.705 4.5125 ;
      RECT  621.12 4.0975 623.565 4.5125 ;
      RECT  623.98 4.0975 626.425 4.5125 ;
      RECT  626.84 4.0975 629.285 4.5125 ;
      RECT  629.7 4.0975 632.145 4.5125 ;
      RECT  632.56 4.0975 635.005 4.5125 ;
      RECT  635.42 4.0975 637.865 4.5125 ;
      RECT  638.28 4.0975 640.725 4.5125 ;
      RECT  641.14 4.0975 643.585 4.5125 ;
      RECT  644.0 4.0975 646.445 4.5125 ;
      RECT  646.86 4.0975 649.305 4.5125 ;
      RECT  649.72 4.0975 652.165 4.5125 ;
      RECT  652.58 4.0975 655.025 4.5125 ;
      RECT  655.44 4.0975 657.885 4.5125 ;
      RECT  658.3 4.0975 660.745 4.5125 ;
      RECT  661.16 4.0975 663.605 4.5125 ;
      RECT  664.02 4.0975 666.465 4.5125 ;
      RECT  666.88 4.0975 669.325 4.5125 ;
      RECT  669.74 4.0975 672.185 4.5125 ;
      RECT  672.6 4.0975 675.045 4.5125 ;
      RECT  675.46 4.0975 677.905 4.5125 ;
      RECT  678.32 4.0975 680.765 4.5125 ;
      RECT  681.18 4.0975 683.625 4.5125 ;
      RECT  684.04 4.0975 686.485 4.5125 ;
      RECT  686.9 4.0975 689.345 4.5125 ;
      RECT  689.76 4.0975 692.205 4.5125 ;
      RECT  692.62 4.0975 695.065 4.5125 ;
      RECT  695.48 4.0975 697.925 4.5125 ;
      RECT  698.34 4.0975 700.785 4.5125 ;
      RECT  701.2 4.0975 703.645 4.5125 ;
      RECT  704.06 4.0975 706.505 4.5125 ;
      RECT  706.92 4.0975 709.365 4.5125 ;
      RECT  709.78 4.0975 712.225 4.5125 ;
      RECT  712.64 4.0975 715.085 4.5125 ;
      RECT  715.5 4.0975 717.945 4.5125 ;
      RECT  718.36 4.0975 720.805 4.5125 ;
      RECT  721.22 4.0975 723.665 4.5125 ;
      RECT  724.08 4.0975 726.525 4.5125 ;
      RECT  726.94 4.0975 729.385 4.5125 ;
      RECT  729.8 4.0975 732.245 4.5125 ;
      RECT  732.66 4.0975 735.105 4.5125 ;
      RECT  735.52 4.0975 737.965 4.5125 ;
      RECT  738.38 4.0975 740.825 4.5125 ;
      RECT  741.24 4.0975 743.685 4.5125 ;
      RECT  744.1 4.0975 746.545 4.5125 ;
      RECT  746.96 4.0975 749.405 4.5125 ;
      RECT  749.82 4.0975 752.265 4.5125 ;
      RECT  752.68 4.0975 755.125 4.5125 ;
      RECT  755.54 4.0975 757.985 4.5125 ;
      RECT  758.4 4.0975 760.845 4.5125 ;
      RECT  761.26 4.0975 763.705 4.5125 ;
      RECT  764.12 4.0975 766.565 4.5125 ;
      RECT  766.98 4.0975 769.425 4.5125 ;
      RECT  769.84 4.0975 772.285 4.5125 ;
      RECT  772.7 4.0975 775.145 4.5125 ;
      RECT  775.56 4.0975 778.005 4.5125 ;
      RECT  778.42 4.0975 780.865 4.5125 ;
      RECT  781.28 4.0975 783.725 4.5125 ;
      RECT  784.14 4.0975 786.585 4.5125 ;
      RECT  787.0 4.0975 789.445 4.5125 ;
      RECT  789.86 4.0975 792.305 4.5125 ;
      RECT  792.72 4.0975 795.165 4.5125 ;
      RECT  795.58 4.0975 798.025 4.5125 ;
      RECT  798.44 4.0975 800.885 4.5125 ;
      RECT  801.3 4.0975 803.745 4.5125 ;
      RECT  804.16 4.0975 806.605 4.5125 ;
      RECT  807.02 4.0975 809.465 4.5125 ;
      RECT  809.88 4.0975 812.325 4.5125 ;
      RECT  812.74 4.0975 815.185 4.5125 ;
      RECT  815.6 4.0975 818.045 4.5125 ;
      RECT  818.46 4.0975 820.905 4.5125 ;
      RECT  821.32 4.0975 823.765 4.5125 ;
      RECT  824.18 4.0975 826.625 4.5125 ;
      RECT  827.04 4.0975 829.485 4.5125 ;
      RECT  829.9 4.0975 832.345 4.5125 ;
      RECT  832.76 4.0975 835.205 4.5125 ;
      RECT  835.62 4.0975 838.065 4.5125 ;
      RECT  838.48 4.0975 840.925 4.5125 ;
      RECT  841.34 4.0975 843.785 4.5125 ;
      RECT  844.2 4.0975 846.645 4.5125 ;
      RECT  847.06 4.0975 849.505 4.5125 ;
      RECT  849.92 4.0975 852.365 4.5125 ;
      RECT  852.78 4.0975 855.225 4.5125 ;
      RECT  855.64 4.0975 858.085 4.5125 ;
      RECT  858.5 4.0975 860.945 4.5125 ;
      RECT  861.36 4.0975 863.805 4.5125 ;
      RECT  864.22 4.0975 866.665 4.5125 ;
      RECT  867.08 4.0975 869.525 4.5125 ;
      RECT  869.94 4.0975 872.385 4.5125 ;
      RECT  872.8 4.0975 875.245 4.5125 ;
      RECT  875.66 4.0975 878.105 4.5125 ;
      RECT  878.52 4.0975 880.965 4.5125 ;
      RECT  881.38 4.0975 883.825 4.5125 ;
      RECT  884.24 4.0975 886.685 4.5125 ;
      RECT  887.1 4.0975 889.545 4.5125 ;
      RECT  889.96 4.0975 892.405 4.5125 ;
      RECT  892.82 4.0975 895.265 4.5125 ;
      RECT  895.68 4.0975 898.125 4.5125 ;
      RECT  898.54 4.0975 900.985 4.5125 ;
      RECT  901.4 4.0975 903.845 4.5125 ;
      RECT  904.26 4.0975 906.705 4.5125 ;
      RECT  907.12 4.0975 909.565 4.5125 ;
      RECT  909.98 4.0975 912.425 4.5125 ;
      RECT  912.84 4.0975 915.285 4.5125 ;
      RECT  915.7 4.0975 918.145 4.5125 ;
      RECT  918.56 4.0975 921.005 4.5125 ;
      RECT  921.42 4.0975 923.865 4.5125 ;
      RECT  924.28 4.0975 926.725 4.5125 ;
      RECT  927.14 4.0975 929.585 4.5125 ;
      RECT  930.0 4.0975 932.445 4.5125 ;
      RECT  932.86 4.0975 935.305 4.5125 ;
      RECT  935.72 4.0975 938.165 4.5125 ;
      RECT  938.58 4.0975 941.025 4.5125 ;
      RECT  941.44 4.0975 943.885 4.5125 ;
      RECT  944.3 4.0975 946.745 4.5125 ;
      RECT  947.16 4.0975 949.605 4.5125 ;
      RECT  950.02 4.0975 952.465 4.5125 ;
      RECT  952.88 4.0975 955.325 4.5125 ;
      RECT  955.74 4.0975 958.185 4.5125 ;
      RECT  958.6 4.0975 961.045 4.5125 ;
      RECT  961.46 4.0975 963.905 4.5125 ;
      RECT  964.32 4.0975 966.765 4.5125 ;
      RECT  967.18 4.0975 969.625 4.5125 ;
      RECT  970.04 4.0975 972.485 4.5125 ;
      RECT  972.9 4.0975 975.345 4.5125 ;
      RECT  975.76 4.0975 978.205 4.5125 ;
      RECT  978.62 4.0975 981.065 4.5125 ;
      RECT  981.48 4.0975 983.925 4.5125 ;
      RECT  984.34 4.0975 986.785 4.5125 ;
      RECT  987.2 4.0975 989.645 4.5125 ;
      RECT  990.06 4.0975 992.505 4.5125 ;
      RECT  992.92 4.0975 995.365 4.5125 ;
      RECT  995.78 4.0975 998.225 4.5125 ;
      RECT  998.64 4.0975 1001.085 4.5125 ;
      RECT  1001.5 4.0975 1003.945 4.5125 ;
      RECT  1004.36 4.0975 1006.805 4.5125 ;
      RECT  1007.22 4.0975 1009.665 4.5125 ;
      RECT  1010.08 4.0975 1012.525 4.5125 ;
      RECT  1012.94 4.0975 1015.385 4.5125 ;
      RECT  1015.8 4.0975 1018.245 4.5125 ;
      RECT  1018.66 4.0975 1021.105 4.5125 ;
      RECT  1021.52 4.0975 1023.965 4.5125 ;
      RECT  1024.38 4.0975 1026.825 4.5125 ;
      RECT  1027.24 4.0975 1029.685 4.5125 ;
      RECT  1030.1 4.0975 1032.545 4.5125 ;
      RECT  1032.96 4.0975 1035.405 4.5125 ;
      RECT  1035.82 4.0975 1038.265 4.5125 ;
      RECT  1038.68 4.0975 1041.125 4.5125 ;
      RECT  1041.54 4.0975 1043.985 4.5125 ;
      RECT  1044.4 4.0975 1046.845 4.5125 ;
      RECT  1047.26 4.0975 1049.705 4.5125 ;
      RECT  1050.12 4.0975 1052.565 4.5125 ;
      RECT  1052.98 4.0975 1055.425 4.5125 ;
      RECT  1055.84 4.0975 1058.285 4.5125 ;
      RECT  1058.7 4.0975 1061.145 4.5125 ;
      RECT  1061.56 4.0975 1064.005 4.5125 ;
      RECT  1064.42 4.0975 1066.865 4.5125 ;
      RECT  1067.28 4.0975 1069.725 4.5125 ;
      RECT  1070.14 4.0975 1072.585 4.5125 ;
      RECT  1073.0 4.0975 1075.445 4.5125 ;
      RECT  1075.86 4.0975 1078.305 4.5125 ;
      RECT  1078.72 4.0975 1081.165 4.5125 ;
      RECT  1081.58 4.0975 1084.025 4.5125 ;
      RECT  1084.44 4.0975 1086.885 4.5125 ;
      RECT  1087.3 4.0975 1089.745 4.5125 ;
      RECT  1090.16 4.0975 1092.605 4.5125 ;
      RECT  1093.02 4.0975 1095.465 4.5125 ;
      RECT  1095.88 4.0975 1098.325 4.5125 ;
      RECT  1098.74 4.0975 1101.185 4.5125 ;
      RECT  1101.6 4.0975 1104.045 4.5125 ;
      RECT  1104.46 4.0975 1106.905 4.5125 ;
      RECT  1107.32 4.0975 1109.765 4.5125 ;
      RECT  1110.18 4.0975 1112.625 4.5125 ;
      RECT  1113.04 4.0975 1115.485 4.5125 ;
      RECT  1115.9 4.0975 1118.345 4.5125 ;
      RECT  1118.76 4.0975 1121.205 4.5125 ;
      RECT  1121.62 4.0975 1124.065 4.5125 ;
      RECT  1124.48 4.0975 1126.925 4.5125 ;
      RECT  1127.34 4.0975 1129.785 4.5125 ;
      RECT  1130.2 4.0975 1132.645 4.5125 ;
      RECT  1133.06 4.0975 1135.505 4.5125 ;
      RECT  1135.92 4.0975 1138.365 4.5125 ;
      RECT  1138.78 4.0975 1141.225 4.5125 ;
      RECT  1141.64 4.0975 1144.085 4.5125 ;
      RECT  1144.5 4.0975 1146.945 4.5125 ;
      RECT  1147.36 4.0975 1149.805 4.5125 ;
      RECT  1150.22 4.0975 1152.665 4.5125 ;
      RECT  1153.08 4.0975 1155.525 4.5125 ;
      RECT  1155.94 4.0975 1158.385 4.5125 ;
      RECT  1158.8 4.0975 1161.245 4.5125 ;
      RECT  1161.66 4.0975 1164.105 4.5125 ;
      RECT  1164.52 4.0975 1166.965 4.5125 ;
      RECT  1167.38 4.0975 1169.825 4.5125 ;
      RECT  1170.24 4.0975 1172.685 4.5125 ;
      RECT  1173.1 4.0975 1175.545 4.5125 ;
      RECT  1175.96 4.0975 1178.405 4.5125 ;
      RECT  1178.82 4.0975 1181.265 4.5125 ;
      RECT  1181.68 4.0975 1184.125 4.5125 ;
      RECT  1184.54 4.0975 1186.985 4.5125 ;
      RECT  1187.4 4.0975 1189.845 4.5125 ;
      RECT  1190.26 4.0975 1192.705 4.5125 ;
      RECT  1193.12 4.0975 1195.565 4.5125 ;
      RECT  1195.98 4.0975 1198.425 4.5125 ;
      RECT  1198.84 4.0975 1201.285 4.5125 ;
      RECT  1201.7 4.0975 1204.145 4.5125 ;
      RECT  1204.56 4.0975 1207.005 4.5125 ;
      RECT  1207.42 4.0975 1209.865 4.5125 ;
      RECT  1210.28 4.0975 1212.725 4.5125 ;
      RECT  1213.14 4.0975 1215.585 4.5125 ;
      RECT  1216.0 4.0975 1218.445 4.5125 ;
      RECT  1218.86 4.0975 1221.305 4.5125 ;
      RECT  1221.72 4.0975 1224.165 4.5125 ;
      RECT  1224.58 4.0975 1227.025 4.5125 ;
      RECT  1227.44 4.0975 1229.885 4.5125 ;
      RECT  1230.3 4.0975 1232.745 4.5125 ;
      RECT  1233.16 4.0975 1235.605 4.5125 ;
      RECT  1236.02 4.0975 1238.465 4.5125 ;
      RECT  1238.88 4.0975 1241.325 4.5125 ;
      RECT  1241.74 4.0975 1244.185 4.5125 ;
      RECT  1244.6 4.0975 1247.045 4.5125 ;
      RECT  1247.46 4.0975 1249.905 4.5125 ;
      RECT  1250.32 4.0975 1252.765 4.5125 ;
      RECT  1253.18 4.0975 1255.625 4.5125 ;
      RECT  1256.04 4.0975 1258.485 4.5125 ;
      RECT  1258.9 4.0975 1261.345 4.5125 ;
      RECT  1261.76 4.0975 1264.205 4.5125 ;
      RECT  1264.62 4.0975 1267.065 4.5125 ;
      RECT  1267.48 4.0975 1269.925 4.5125 ;
      RECT  1270.34 4.0975 1272.785 4.5125 ;
      RECT  1273.2 4.0975 1275.645 4.5125 ;
      RECT  1276.06 4.0975 1278.505 4.5125 ;
      RECT  1278.92 4.0975 1281.365 4.5125 ;
      RECT  1281.78 4.0975 1284.225 4.5125 ;
      RECT  1284.64 4.0975 1287.085 4.5125 ;
      RECT  1287.5 4.0975 1289.945 4.5125 ;
      RECT  1290.36 4.0975 1292.805 4.5125 ;
      RECT  1293.22 4.0975 1295.665 4.5125 ;
      RECT  1296.08 4.0975 1298.525 4.5125 ;
      RECT  1298.94 4.0975 1301.385 4.5125 ;
      RECT  1301.8 4.0975 1304.245 4.5125 ;
      RECT  1304.66 4.0975 1307.105 4.5125 ;
      RECT  1307.52 4.0975 1309.965 4.5125 ;
      RECT  1310.38 4.0975 1312.825 4.5125 ;
      RECT  1313.24 4.0975 1315.685 4.5125 ;
      RECT  1316.1 4.0975 1318.545 4.5125 ;
      RECT  1318.96 4.0975 1321.405 4.5125 ;
      RECT  1321.82 4.0975 1324.265 4.5125 ;
      RECT  1324.68 4.0975 1327.125 4.5125 ;
      RECT  1327.54 4.0975 1329.985 4.5125 ;
      RECT  1330.4 4.0975 1332.845 4.5125 ;
      RECT  1333.26 4.0975 1335.705 4.5125 ;
      RECT  1336.12 4.0975 1338.565 4.5125 ;
      RECT  1338.98 4.0975 1341.425 4.5125 ;
      RECT  1341.84 4.0975 1344.285 4.5125 ;
      RECT  1344.7 4.0975 1347.145 4.5125 ;
      RECT  1347.56 4.0975 1350.005 4.5125 ;
      RECT  1350.42 4.0975 1352.865 4.5125 ;
      RECT  1353.28 4.0975 1355.725 4.5125 ;
      RECT  1356.14 4.0975 1358.585 4.5125 ;
      RECT  1359.0 4.0975 1361.445 4.5125 ;
      RECT  1361.86 4.0975 1364.305 4.5125 ;
      RECT  1364.72 4.0975 1367.165 4.5125 ;
      RECT  1367.58 4.0975 1370.025 4.5125 ;
      RECT  1370.44 4.0975 1372.885 4.5125 ;
      RECT  1373.3 4.0975 1375.745 4.5125 ;
      RECT  1376.16 4.0975 1378.605 4.5125 ;
      RECT  1379.02 4.0975 1381.465 4.5125 ;
      RECT  1381.88 4.0975 1384.325 4.5125 ;
      RECT  1384.74 4.0975 1387.185 4.5125 ;
      RECT  1387.6 4.0975 1390.045 4.5125 ;
      RECT  1390.46 4.0975 1392.905 4.5125 ;
      RECT  1393.32 4.0975 1395.765 4.5125 ;
      RECT  1396.18 4.0975 1398.625 4.5125 ;
      RECT  1399.04 4.0975 1401.485 4.5125 ;
      RECT  1401.9 4.0975 1404.345 4.5125 ;
      RECT  1404.76 4.0975 1407.205 4.5125 ;
      RECT  1407.62 4.0975 1410.065 4.5125 ;
      RECT  1410.48 4.0975 1412.925 4.5125 ;
      RECT  1413.34 4.0975 1415.785 4.5125 ;
      RECT  1416.2 4.0975 1418.645 4.5125 ;
      RECT  1419.06 4.0975 1421.505 4.5125 ;
      RECT  1421.92 4.0975 1424.365 4.5125 ;
      RECT  1424.78 4.0975 1427.225 4.5125 ;
      RECT  1427.64 4.0975 1430.085 4.5125 ;
      RECT  1430.5 4.0975 1432.945 4.5125 ;
      RECT  1433.36 4.0975 1435.805 4.5125 ;
      RECT  1436.22 4.0975 1438.665 4.5125 ;
      RECT  1439.08 4.0975 1441.525 4.5125 ;
      RECT  1441.94 4.0975 1444.385 4.5125 ;
      RECT  1444.8 4.0975 1447.245 4.5125 ;
      RECT  1447.66 4.0975 1450.105 4.5125 ;
      RECT  1450.52 4.0975 1452.965 4.5125 ;
      RECT  1453.38 4.0975 1455.825 4.5125 ;
      RECT  1456.24 4.0975 1458.685 4.5125 ;
      RECT  1459.1 4.0975 1461.545 4.5125 ;
      RECT  1461.96 4.0975 1464.405 4.5125 ;
      RECT  1464.82 4.0975 1467.265 4.5125 ;
      RECT  1467.68 4.0975 1470.125 4.5125 ;
      RECT  1470.54 4.0975 1472.985 4.5125 ;
      RECT  1473.4 4.0975 1475.845 4.5125 ;
      RECT  1476.26 4.0975 1478.705 4.5125 ;
      RECT  1479.12 4.0975 1481.565 4.5125 ;
      RECT  1481.98 4.0975 1484.425 4.5125 ;
      RECT  1484.84 4.0975 1487.285 4.5125 ;
      RECT  1487.7 4.0975 1490.145 4.5125 ;
      RECT  1490.56 4.0975 1493.005 4.5125 ;
      RECT  1493.42 4.0975 1495.865 4.5125 ;
      RECT  1496.28 4.0975 1498.725 4.5125 ;
      RECT  1499.14 4.0975 1501.585 4.5125 ;
      RECT  1502.0 4.0975 1504.445 4.5125 ;
      RECT  1504.86 4.0975 1507.305 4.5125 ;
      RECT  1507.72 4.0975 1510.165 4.5125 ;
      RECT  1510.58 4.0975 1513.025 4.5125 ;
      RECT  1513.44 4.0975 1515.885 4.5125 ;
      RECT  1516.3 4.0975 1518.745 4.5125 ;
      RECT  1519.16 4.0975 1521.605 4.5125 ;
      RECT  1522.02 4.0975 1524.465 4.5125 ;
      RECT  1524.88 4.0975 1527.325 4.5125 ;
      RECT  1527.74 4.0975 1530.185 4.5125 ;
      RECT  1530.6 4.0975 1533.045 4.5125 ;
      RECT  1533.46 4.0975 1535.905 4.5125 ;
      RECT  1536.32 4.0975 1538.765 4.5125 ;
      RECT  1539.18 4.0975 1541.625 4.5125 ;
      RECT  1542.04 4.0975 1544.485 4.5125 ;
      RECT  1544.9 4.0975 1547.345 4.5125 ;
      RECT  1547.76 4.0975 1550.205 4.5125 ;
      RECT  1550.62 4.0975 1553.065 4.5125 ;
      RECT  1553.48 4.0975 1555.925 4.5125 ;
      RECT  1556.34 4.0975 1558.785 4.5125 ;
      RECT  1559.2 4.0975 1561.645 4.5125 ;
      RECT  1562.06 4.0975 1564.505 4.5125 ;
      RECT  1564.92 4.0975 1567.365 4.5125 ;
      RECT  1567.78 4.0975 1570.225 4.5125 ;
      RECT  1570.64 4.0975 1573.085 4.5125 ;
      RECT  1573.5 4.0975 1575.945 4.5125 ;
      RECT  1576.36 4.0975 1578.805 4.5125 ;
      RECT  1579.22 4.0975 1581.665 4.5125 ;
      RECT  1582.08 4.0975 1584.525 4.5125 ;
      RECT  1584.94 4.0975 1587.385 4.5125 ;
      RECT  1587.8 4.0975 1593.2 4.5125 ;
      RECT  0.14 122.2925 120.205 122.7075 ;
      RECT  120.205 4.5125 120.62 122.2925 ;
      RECT  120.62 4.5125 125.925 122.2925 ;
      RECT  120.62 122.2925 125.925 122.7075 ;
      RECT  120.205 122.7075 120.62 125.0225 ;
      RECT  120.205 125.4375 120.62 127.2325 ;
      RECT  120.205 127.6475 120.62 129.9625 ;
      RECT  120.205 130.3775 120.62 132.1725 ;
      RECT  120.205 132.5875 120.62 134.9025 ;
      RECT  126.34 4.5125 801.085 96.1625 ;
      RECT  126.34 96.1625 801.085 96.5775 ;
      RECT  801.5 4.5125 1593.2 96.1625 ;
      RECT  801.5 96.1625 1593.2 96.5775 ;
      RECT  801.085 93.8475 801.5 96.1625 ;
      RECT  801.085 91.6375 801.5 93.4325 ;
      RECT  801.085 88.9075 801.5 91.2225 ;
      RECT  801.085 86.6975 801.5 88.4925 ;
      RECT  801.085 4.5125 801.5 83.5525 ;
      RECT  801.085 83.9675 801.5 86.2825 ;
      RECT  0.14 4.5125 3.245 77.7025 ;
      RECT  0.14 77.7025 3.245 78.1175 ;
      RECT  0.14 78.1175 3.245 122.2925 ;
      RECT  3.245 4.5125 3.66 77.7025 ;
      RECT  3.245 78.1175 3.66 122.2925 ;
      RECT  3.66 4.5125 120.205 77.7025 ;
      RECT  918.185 96.5775 918.6 209.8625 ;
      RECT  918.6 96.5775 1593.2 209.8625 ;
      RECT  918.6 209.8625 1593.2 210.2775 ;
      RECT  3.66 77.7025 9.2075 77.7875 ;
      RECT  3.66 77.7875 9.2075 78.1175 ;
      RECT  9.2075 77.7025 9.6225 77.7875 ;
      RECT  9.6225 77.7025 120.205 77.7875 ;
      RECT  9.6225 77.7875 120.205 78.1175 ;
      RECT  3.66 78.1175 9.2075 78.2025 ;
      RECT  3.66 78.2025 9.2075 122.2925 ;
      RECT  9.2075 78.2025 9.6225 122.2925 ;
      RECT  9.6225 78.1175 120.205 78.2025 ;
      RECT  9.6225 78.2025 120.205 122.2925 ;
      RECT  801.5 96.5775 912.0825 209.7775 ;
      RECT  801.5 209.7775 912.0825 209.8625 ;
      RECT  912.0825 96.5775 912.4975 209.7775 ;
      RECT  912.4975 96.5775 918.185 209.7775 ;
      RECT  912.4975 209.7775 918.185 209.8625 ;
      RECT  801.5 209.8625 912.0825 210.1925 ;
      RECT  801.5 210.1925 912.0825 210.2775 ;
      RECT  912.0825 210.1925 912.4975 210.2775 ;
      RECT  912.4975 209.8625 918.185 210.1925 ;
      RECT  912.4975 210.1925 918.185 210.2775 ;
      RECT  126.34 96.5775 159.7825 203.155 ;
      RECT  126.34 203.155 159.7825 203.57 ;
      RECT  159.7825 96.5775 160.1975 203.155 ;
      RECT  160.1975 96.5775 801.085 203.155 ;
      RECT  160.1975 203.155 160.9575 203.57 ;
      RECT  161.3725 203.155 162.1325 203.57 ;
      RECT  162.5475 203.155 163.3075 203.57 ;
      RECT  163.7225 203.155 164.4825 203.57 ;
      RECT  164.8975 203.155 165.6575 203.57 ;
      RECT  166.0725 203.155 166.8325 203.57 ;
      RECT  167.2475 203.155 168.0075 203.57 ;
      RECT  168.4225 203.155 169.1825 203.57 ;
      RECT  169.5975 203.155 170.3575 203.57 ;
      RECT  170.7725 203.155 171.5325 203.57 ;
      RECT  171.9475 203.155 172.7075 203.57 ;
      RECT  173.1225 203.155 173.8825 203.57 ;
      RECT  174.2975 203.155 175.0575 203.57 ;
      RECT  175.4725 203.155 176.2325 203.57 ;
      RECT  176.6475 203.155 177.4075 203.57 ;
      RECT  177.8225 203.155 178.5825 203.57 ;
      RECT  178.9975 203.155 179.7575 203.57 ;
      RECT  180.1725 203.155 180.9325 203.57 ;
      RECT  181.3475 203.155 182.1075 203.57 ;
      RECT  182.5225 203.155 183.2825 203.57 ;
      RECT  183.6975 203.155 184.4575 203.57 ;
      RECT  184.8725 203.155 185.6325 203.57 ;
      RECT  186.0475 203.155 186.8075 203.57 ;
      RECT  187.2225 203.155 187.9825 203.57 ;
      RECT  188.3975 203.155 189.1575 203.57 ;
      RECT  189.5725 203.155 190.3325 203.57 ;
      RECT  190.7475 203.155 191.5075 203.57 ;
      RECT  191.9225 203.155 192.6825 203.57 ;
      RECT  193.0975 203.155 193.8575 203.57 ;
      RECT  194.2725 203.155 195.0325 203.57 ;
      RECT  195.4475 203.155 196.2075 203.57 ;
      RECT  196.6225 203.155 197.3825 203.57 ;
      RECT  197.7975 203.155 198.5575 203.57 ;
      RECT  198.9725 203.155 199.7325 203.57 ;
      RECT  200.1475 203.155 200.9075 203.57 ;
      RECT  201.3225 203.155 202.0825 203.57 ;
      RECT  202.4975 203.155 203.2575 203.57 ;
      RECT  203.6725 203.155 204.4325 203.57 ;
      RECT  204.8475 203.155 205.6075 203.57 ;
      RECT  206.0225 203.155 206.7825 203.57 ;
      RECT  207.1975 203.155 207.9575 203.57 ;
      RECT  208.3725 203.155 209.1325 203.57 ;
      RECT  209.5475 203.155 210.3075 203.57 ;
      RECT  210.7225 203.155 211.4825 203.57 ;
      RECT  211.8975 203.155 212.6575 203.57 ;
      RECT  213.0725 203.155 213.8325 203.57 ;
      RECT  214.2475 203.155 215.0075 203.57 ;
      RECT  215.4225 203.155 216.1825 203.57 ;
      RECT  216.5975 203.155 217.3575 203.57 ;
      RECT  217.7725 203.155 218.5325 203.57 ;
      RECT  218.9475 203.155 219.7075 203.57 ;
      RECT  220.1225 203.155 220.8825 203.57 ;
      RECT  221.2975 203.155 222.0575 203.57 ;
      RECT  222.4725 203.155 223.2325 203.57 ;
      RECT  223.6475 203.155 224.4075 203.57 ;
      RECT  224.8225 203.155 225.5825 203.57 ;
      RECT  225.9975 203.155 226.7575 203.57 ;
      RECT  227.1725 203.155 227.9325 203.57 ;
      RECT  228.3475 203.155 229.1075 203.57 ;
      RECT  229.5225 203.155 230.2825 203.57 ;
      RECT  230.6975 203.155 231.4575 203.57 ;
      RECT  231.8725 203.155 232.6325 203.57 ;
      RECT  233.0475 203.155 233.8075 203.57 ;
      RECT  234.2225 203.155 234.9825 203.57 ;
      RECT  235.3975 203.155 236.1575 203.57 ;
      RECT  236.5725 203.155 237.3325 203.57 ;
      RECT  237.7475 203.155 238.5075 203.57 ;
      RECT  238.9225 203.155 239.6825 203.57 ;
      RECT  240.0975 203.155 240.8575 203.57 ;
      RECT  241.2725 203.155 242.0325 203.57 ;
      RECT  242.4475 203.155 243.2075 203.57 ;
      RECT  243.6225 203.155 244.3825 203.57 ;
      RECT  244.7975 203.155 245.5575 203.57 ;
      RECT  245.9725 203.155 246.7325 203.57 ;
      RECT  247.1475 203.155 247.9075 203.57 ;
      RECT  248.3225 203.155 249.0825 203.57 ;
      RECT  249.4975 203.155 250.2575 203.57 ;
      RECT  250.6725 203.155 251.4325 203.57 ;
      RECT  251.8475 203.155 252.6075 203.57 ;
      RECT  253.0225 203.155 253.7825 203.57 ;
      RECT  254.1975 203.155 254.9575 203.57 ;
      RECT  255.3725 203.155 256.1325 203.57 ;
      RECT  256.5475 203.155 257.3075 203.57 ;
      RECT  257.7225 203.155 258.4825 203.57 ;
      RECT  258.8975 203.155 259.6575 203.57 ;
      RECT  260.0725 203.155 260.8325 203.57 ;
      RECT  261.2475 203.155 262.0075 203.57 ;
      RECT  262.4225 203.155 263.1825 203.57 ;
      RECT  263.5975 203.155 264.3575 203.57 ;
      RECT  264.7725 203.155 265.5325 203.57 ;
      RECT  265.9475 203.155 266.7075 203.57 ;
      RECT  267.1225 203.155 267.8825 203.57 ;
      RECT  268.2975 203.155 269.0575 203.57 ;
      RECT  269.4725 203.155 270.2325 203.57 ;
      RECT  270.6475 203.155 271.4075 203.57 ;
      RECT  271.8225 203.155 272.5825 203.57 ;
      RECT  272.9975 203.155 273.7575 203.57 ;
      RECT  274.1725 203.155 274.9325 203.57 ;
      RECT  275.3475 203.155 276.1075 203.57 ;
      RECT  276.5225 203.155 277.2825 203.57 ;
      RECT  277.6975 203.155 278.4575 203.57 ;
      RECT  278.8725 203.155 279.6325 203.57 ;
      RECT  280.0475 203.155 280.8075 203.57 ;
      RECT  281.2225 203.155 281.9825 203.57 ;
      RECT  282.3975 203.155 283.1575 203.57 ;
      RECT  283.5725 203.155 284.3325 203.57 ;
      RECT  284.7475 203.155 285.5075 203.57 ;
      RECT  285.9225 203.155 286.6825 203.57 ;
      RECT  287.0975 203.155 287.8575 203.57 ;
      RECT  288.2725 203.155 289.0325 203.57 ;
      RECT  289.4475 203.155 290.2075 203.57 ;
      RECT  290.6225 203.155 291.3825 203.57 ;
      RECT  291.7975 203.155 292.5575 203.57 ;
      RECT  292.9725 203.155 293.7325 203.57 ;
      RECT  294.1475 203.155 294.9075 203.57 ;
      RECT  295.3225 203.155 296.0825 203.57 ;
      RECT  296.4975 203.155 297.2575 203.57 ;
      RECT  297.6725 203.155 298.4325 203.57 ;
      RECT  298.8475 203.155 299.6075 203.57 ;
      RECT  300.0225 203.155 300.7825 203.57 ;
      RECT  301.1975 203.155 301.9575 203.57 ;
      RECT  302.3725 203.155 303.1325 203.57 ;
      RECT  303.5475 203.155 304.3075 203.57 ;
      RECT  304.7225 203.155 305.4825 203.57 ;
      RECT  305.8975 203.155 306.6575 203.57 ;
      RECT  307.0725 203.155 307.8325 203.57 ;
      RECT  308.2475 203.155 309.0075 203.57 ;
      RECT  309.4225 203.155 310.1825 203.57 ;
      RECT  310.5975 203.155 311.3575 203.57 ;
      RECT  311.7725 203.155 312.5325 203.57 ;
      RECT  312.9475 203.155 313.7075 203.57 ;
      RECT  314.1225 203.155 314.8825 203.57 ;
      RECT  315.2975 203.155 316.0575 203.57 ;
      RECT  316.4725 203.155 317.2325 203.57 ;
      RECT  317.6475 203.155 318.4075 203.57 ;
      RECT  318.8225 203.155 319.5825 203.57 ;
      RECT  319.9975 203.155 320.7575 203.57 ;
      RECT  321.1725 203.155 321.9325 203.57 ;
      RECT  322.3475 203.155 323.1075 203.57 ;
      RECT  323.5225 203.155 324.2825 203.57 ;
      RECT  324.6975 203.155 325.4575 203.57 ;
      RECT  325.8725 203.155 326.6325 203.57 ;
      RECT  327.0475 203.155 327.8075 203.57 ;
      RECT  328.2225 203.155 328.9825 203.57 ;
      RECT  329.3975 203.155 330.1575 203.57 ;
      RECT  330.5725 203.155 331.3325 203.57 ;
      RECT  331.7475 203.155 332.5075 203.57 ;
      RECT  332.9225 203.155 333.6825 203.57 ;
      RECT  334.0975 203.155 334.8575 203.57 ;
      RECT  335.2725 203.155 336.0325 203.57 ;
      RECT  336.4475 203.155 337.2075 203.57 ;
      RECT  337.6225 203.155 338.3825 203.57 ;
      RECT  338.7975 203.155 339.5575 203.57 ;
      RECT  339.9725 203.155 340.7325 203.57 ;
      RECT  341.1475 203.155 341.9075 203.57 ;
      RECT  342.3225 203.155 343.0825 203.57 ;
      RECT  343.4975 203.155 344.2575 203.57 ;
      RECT  344.6725 203.155 345.4325 203.57 ;
      RECT  345.8475 203.155 346.6075 203.57 ;
      RECT  347.0225 203.155 347.7825 203.57 ;
      RECT  348.1975 203.155 348.9575 203.57 ;
      RECT  349.3725 203.155 350.1325 203.57 ;
      RECT  350.5475 203.155 351.3075 203.57 ;
      RECT  351.7225 203.155 352.4825 203.57 ;
      RECT  352.8975 203.155 353.6575 203.57 ;
      RECT  354.0725 203.155 354.8325 203.57 ;
      RECT  355.2475 203.155 356.0075 203.57 ;
      RECT  356.4225 203.155 357.1825 203.57 ;
      RECT  357.5975 203.155 358.3575 203.57 ;
      RECT  358.7725 203.155 359.5325 203.57 ;
      RECT  359.9475 203.155 360.7075 203.57 ;
      RECT  361.1225 203.155 361.8825 203.57 ;
      RECT  362.2975 203.155 363.0575 203.57 ;
      RECT  363.4725 203.155 364.2325 203.57 ;
      RECT  364.6475 203.155 365.4075 203.57 ;
      RECT  365.8225 203.155 366.5825 203.57 ;
      RECT  366.9975 203.155 367.7575 203.57 ;
      RECT  368.1725 203.155 368.9325 203.57 ;
      RECT  369.3475 203.155 370.1075 203.57 ;
      RECT  370.5225 203.155 371.2825 203.57 ;
      RECT  371.6975 203.155 372.4575 203.57 ;
      RECT  372.8725 203.155 373.6325 203.57 ;
      RECT  374.0475 203.155 374.8075 203.57 ;
      RECT  375.2225 203.155 375.9825 203.57 ;
      RECT  376.3975 203.155 377.1575 203.57 ;
      RECT  377.5725 203.155 378.3325 203.57 ;
      RECT  378.7475 203.155 379.5075 203.57 ;
      RECT  379.9225 203.155 380.6825 203.57 ;
      RECT  381.0975 203.155 381.8575 203.57 ;
      RECT  382.2725 203.155 383.0325 203.57 ;
      RECT  383.4475 203.155 384.2075 203.57 ;
      RECT  384.6225 203.155 385.3825 203.57 ;
      RECT  385.7975 203.155 386.5575 203.57 ;
      RECT  386.9725 203.155 387.7325 203.57 ;
      RECT  388.1475 203.155 388.9075 203.57 ;
      RECT  389.3225 203.155 390.0825 203.57 ;
      RECT  390.4975 203.155 391.2575 203.57 ;
      RECT  391.6725 203.155 392.4325 203.57 ;
      RECT  392.8475 203.155 393.6075 203.57 ;
      RECT  394.0225 203.155 394.7825 203.57 ;
      RECT  395.1975 203.155 395.9575 203.57 ;
      RECT  396.3725 203.155 397.1325 203.57 ;
      RECT  397.5475 203.155 398.3075 203.57 ;
      RECT  398.7225 203.155 399.4825 203.57 ;
      RECT  399.8975 203.155 400.6575 203.57 ;
      RECT  401.0725 203.155 401.8325 203.57 ;
      RECT  402.2475 203.155 403.0075 203.57 ;
      RECT  403.4225 203.155 404.1825 203.57 ;
      RECT  404.5975 203.155 405.3575 203.57 ;
      RECT  405.7725 203.155 406.5325 203.57 ;
      RECT  406.9475 203.155 407.7075 203.57 ;
      RECT  408.1225 203.155 408.8825 203.57 ;
      RECT  409.2975 203.155 410.0575 203.57 ;
      RECT  410.4725 203.155 411.2325 203.57 ;
      RECT  411.6475 203.155 412.4075 203.57 ;
      RECT  412.8225 203.155 413.5825 203.57 ;
      RECT  413.9975 203.155 414.7575 203.57 ;
      RECT  415.1725 203.155 415.9325 203.57 ;
      RECT  416.3475 203.155 417.1075 203.57 ;
      RECT  417.5225 203.155 418.2825 203.57 ;
      RECT  418.6975 203.155 419.4575 203.57 ;
      RECT  419.8725 203.155 420.6325 203.57 ;
      RECT  421.0475 203.155 421.8075 203.57 ;
      RECT  422.2225 203.155 422.9825 203.57 ;
      RECT  423.3975 203.155 424.1575 203.57 ;
      RECT  424.5725 203.155 425.3325 203.57 ;
      RECT  425.7475 203.155 426.5075 203.57 ;
      RECT  426.9225 203.155 427.6825 203.57 ;
      RECT  428.0975 203.155 428.8575 203.57 ;
      RECT  429.2725 203.155 430.0325 203.57 ;
      RECT  430.4475 203.155 431.2075 203.57 ;
      RECT  431.6225 203.155 432.3825 203.57 ;
      RECT  432.7975 203.155 433.5575 203.57 ;
      RECT  433.9725 203.155 434.7325 203.57 ;
      RECT  435.1475 203.155 435.9075 203.57 ;
      RECT  436.3225 203.155 437.0825 203.57 ;
      RECT  437.4975 203.155 438.2575 203.57 ;
      RECT  438.6725 203.155 439.4325 203.57 ;
      RECT  439.8475 203.155 440.6075 203.57 ;
      RECT  441.0225 203.155 441.7825 203.57 ;
      RECT  442.1975 203.155 442.9575 203.57 ;
      RECT  443.3725 203.155 444.1325 203.57 ;
      RECT  444.5475 203.155 445.3075 203.57 ;
      RECT  445.7225 203.155 446.4825 203.57 ;
      RECT  446.8975 203.155 447.6575 203.57 ;
      RECT  448.0725 203.155 448.8325 203.57 ;
      RECT  449.2475 203.155 450.0075 203.57 ;
      RECT  450.4225 203.155 451.1825 203.57 ;
      RECT  451.5975 203.155 452.3575 203.57 ;
      RECT  452.7725 203.155 453.5325 203.57 ;
      RECT  453.9475 203.155 454.7075 203.57 ;
      RECT  455.1225 203.155 455.8825 203.57 ;
      RECT  456.2975 203.155 457.0575 203.57 ;
      RECT  457.4725 203.155 458.2325 203.57 ;
      RECT  458.6475 203.155 459.4075 203.57 ;
      RECT  459.8225 203.155 460.5825 203.57 ;
      RECT  460.9975 203.155 461.7575 203.57 ;
      RECT  462.1725 203.155 462.9325 203.57 ;
      RECT  463.3475 203.155 464.1075 203.57 ;
      RECT  464.5225 203.155 465.2825 203.57 ;
      RECT  465.6975 203.155 466.4575 203.57 ;
      RECT  466.8725 203.155 467.6325 203.57 ;
      RECT  468.0475 203.155 468.8075 203.57 ;
      RECT  469.2225 203.155 469.9825 203.57 ;
      RECT  470.3975 203.155 471.1575 203.57 ;
      RECT  471.5725 203.155 472.3325 203.57 ;
      RECT  472.7475 203.155 473.5075 203.57 ;
      RECT  473.9225 203.155 474.6825 203.57 ;
      RECT  475.0975 203.155 475.8575 203.57 ;
      RECT  476.2725 203.155 477.0325 203.57 ;
      RECT  477.4475 203.155 478.2075 203.57 ;
      RECT  478.6225 203.155 479.3825 203.57 ;
      RECT  479.7975 203.155 480.5575 203.57 ;
      RECT  480.9725 203.155 481.7325 203.57 ;
      RECT  482.1475 203.155 482.9075 203.57 ;
      RECT  483.3225 203.155 484.0825 203.57 ;
      RECT  484.4975 203.155 485.2575 203.57 ;
      RECT  485.6725 203.155 486.4325 203.57 ;
      RECT  486.8475 203.155 487.6075 203.57 ;
      RECT  488.0225 203.155 488.7825 203.57 ;
      RECT  489.1975 203.155 489.9575 203.57 ;
      RECT  490.3725 203.155 491.1325 203.57 ;
      RECT  491.5475 203.155 492.3075 203.57 ;
      RECT  492.7225 203.155 493.4825 203.57 ;
      RECT  493.8975 203.155 494.6575 203.57 ;
      RECT  495.0725 203.155 495.8325 203.57 ;
      RECT  496.2475 203.155 497.0075 203.57 ;
      RECT  497.4225 203.155 498.1825 203.57 ;
      RECT  498.5975 203.155 499.3575 203.57 ;
      RECT  499.7725 203.155 500.5325 203.57 ;
      RECT  500.9475 203.155 501.7075 203.57 ;
      RECT  502.1225 203.155 502.8825 203.57 ;
      RECT  503.2975 203.155 504.0575 203.57 ;
      RECT  504.4725 203.155 505.2325 203.57 ;
      RECT  505.6475 203.155 506.4075 203.57 ;
      RECT  506.8225 203.155 507.5825 203.57 ;
      RECT  507.9975 203.155 508.7575 203.57 ;
      RECT  509.1725 203.155 509.9325 203.57 ;
      RECT  510.3475 203.155 511.1075 203.57 ;
      RECT  511.5225 203.155 512.2825 203.57 ;
      RECT  512.6975 203.155 513.4575 203.57 ;
      RECT  513.8725 203.155 514.6325 203.57 ;
      RECT  515.0475 203.155 515.8075 203.57 ;
      RECT  516.2225 203.155 516.9825 203.57 ;
      RECT  517.3975 203.155 518.1575 203.57 ;
      RECT  518.5725 203.155 519.3325 203.57 ;
      RECT  519.7475 203.155 520.5075 203.57 ;
      RECT  520.9225 203.155 521.6825 203.57 ;
      RECT  522.0975 203.155 522.8575 203.57 ;
      RECT  523.2725 203.155 524.0325 203.57 ;
      RECT  524.4475 203.155 525.2075 203.57 ;
      RECT  525.6225 203.155 526.3825 203.57 ;
      RECT  526.7975 203.155 527.5575 203.57 ;
      RECT  527.9725 203.155 528.7325 203.57 ;
      RECT  529.1475 203.155 529.9075 203.57 ;
      RECT  530.3225 203.155 531.0825 203.57 ;
      RECT  531.4975 203.155 532.2575 203.57 ;
      RECT  532.6725 203.155 533.4325 203.57 ;
      RECT  533.8475 203.155 534.6075 203.57 ;
      RECT  535.0225 203.155 535.7825 203.57 ;
      RECT  536.1975 203.155 536.9575 203.57 ;
      RECT  537.3725 203.155 538.1325 203.57 ;
      RECT  538.5475 203.155 539.3075 203.57 ;
      RECT  539.7225 203.155 540.4825 203.57 ;
      RECT  540.8975 203.155 541.6575 203.57 ;
      RECT  542.0725 203.155 542.8325 203.57 ;
      RECT  543.2475 203.155 544.0075 203.57 ;
      RECT  544.4225 203.155 545.1825 203.57 ;
      RECT  545.5975 203.155 546.3575 203.57 ;
      RECT  546.7725 203.155 547.5325 203.57 ;
      RECT  547.9475 203.155 548.7075 203.57 ;
      RECT  549.1225 203.155 549.8825 203.57 ;
      RECT  550.2975 203.155 551.0575 203.57 ;
      RECT  551.4725 203.155 552.2325 203.57 ;
      RECT  552.6475 203.155 553.4075 203.57 ;
      RECT  553.8225 203.155 554.5825 203.57 ;
      RECT  554.9975 203.155 555.7575 203.57 ;
      RECT  556.1725 203.155 556.9325 203.57 ;
      RECT  557.3475 203.155 558.1075 203.57 ;
      RECT  558.5225 203.155 559.2825 203.57 ;
      RECT  559.6975 203.155 560.4575 203.57 ;
      RECT  560.8725 203.155 561.6325 203.57 ;
      RECT  562.0475 203.155 562.8075 203.57 ;
      RECT  563.2225 203.155 563.9825 203.57 ;
      RECT  564.3975 203.155 565.1575 203.57 ;
      RECT  565.5725 203.155 566.3325 203.57 ;
      RECT  566.7475 203.155 567.5075 203.57 ;
      RECT  567.9225 203.155 568.6825 203.57 ;
      RECT  569.0975 203.155 569.8575 203.57 ;
      RECT  570.2725 203.155 571.0325 203.57 ;
      RECT  571.4475 203.155 572.2075 203.57 ;
      RECT  572.6225 203.155 573.3825 203.57 ;
      RECT  573.7975 203.155 574.5575 203.57 ;
      RECT  574.9725 203.155 575.7325 203.57 ;
      RECT  576.1475 203.155 576.9075 203.57 ;
      RECT  577.3225 203.155 578.0825 203.57 ;
      RECT  578.4975 203.155 579.2575 203.57 ;
      RECT  579.6725 203.155 580.4325 203.57 ;
      RECT  580.8475 203.155 581.6075 203.57 ;
      RECT  582.0225 203.155 582.7825 203.57 ;
      RECT  583.1975 203.155 583.9575 203.57 ;
      RECT  584.3725 203.155 585.1325 203.57 ;
      RECT  585.5475 203.155 586.3075 203.57 ;
      RECT  586.7225 203.155 587.4825 203.57 ;
      RECT  587.8975 203.155 588.6575 203.57 ;
      RECT  589.0725 203.155 589.8325 203.57 ;
      RECT  590.2475 203.155 591.0075 203.57 ;
      RECT  591.4225 203.155 592.1825 203.57 ;
      RECT  592.5975 203.155 593.3575 203.57 ;
      RECT  593.7725 203.155 594.5325 203.57 ;
      RECT  594.9475 203.155 595.7075 203.57 ;
      RECT  596.1225 203.155 596.8825 203.57 ;
      RECT  597.2975 203.155 598.0575 203.57 ;
      RECT  598.4725 203.155 599.2325 203.57 ;
      RECT  599.6475 203.155 600.4075 203.57 ;
      RECT  600.8225 203.155 601.5825 203.57 ;
      RECT  601.9975 203.155 602.7575 203.57 ;
      RECT  603.1725 203.155 603.9325 203.57 ;
      RECT  604.3475 203.155 605.1075 203.57 ;
      RECT  605.5225 203.155 606.2825 203.57 ;
      RECT  606.6975 203.155 607.4575 203.57 ;
      RECT  607.8725 203.155 608.6325 203.57 ;
      RECT  609.0475 203.155 609.8075 203.57 ;
      RECT  610.2225 203.155 610.9825 203.57 ;
      RECT  611.3975 203.155 612.1575 203.57 ;
      RECT  612.5725 203.155 613.3325 203.57 ;
      RECT  613.7475 203.155 614.5075 203.57 ;
      RECT  614.9225 203.155 615.6825 203.57 ;
      RECT  616.0975 203.155 616.8575 203.57 ;
      RECT  617.2725 203.155 618.0325 203.57 ;
      RECT  618.4475 203.155 619.2075 203.57 ;
      RECT  619.6225 203.155 620.3825 203.57 ;
      RECT  620.7975 203.155 621.5575 203.57 ;
      RECT  621.9725 203.155 622.7325 203.57 ;
      RECT  623.1475 203.155 623.9075 203.57 ;
      RECT  624.3225 203.155 625.0825 203.57 ;
      RECT  625.4975 203.155 626.2575 203.57 ;
      RECT  626.6725 203.155 627.4325 203.57 ;
      RECT  627.8475 203.155 628.6075 203.57 ;
      RECT  629.0225 203.155 629.7825 203.57 ;
      RECT  630.1975 203.155 630.9575 203.57 ;
      RECT  631.3725 203.155 632.1325 203.57 ;
      RECT  632.5475 203.155 633.3075 203.57 ;
      RECT  633.7225 203.155 634.4825 203.57 ;
      RECT  634.8975 203.155 635.6575 203.57 ;
      RECT  636.0725 203.155 636.8325 203.57 ;
      RECT  637.2475 203.155 638.0075 203.57 ;
      RECT  638.4225 203.155 639.1825 203.57 ;
      RECT  639.5975 203.155 640.3575 203.57 ;
      RECT  640.7725 203.155 641.5325 203.57 ;
      RECT  641.9475 203.155 642.7075 203.57 ;
      RECT  643.1225 203.155 643.8825 203.57 ;
      RECT  644.2975 203.155 645.0575 203.57 ;
      RECT  645.4725 203.155 646.2325 203.57 ;
      RECT  646.6475 203.155 647.4075 203.57 ;
      RECT  647.8225 203.155 648.5825 203.57 ;
      RECT  648.9975 203.155 649.7575 203.57 ;
      RECT  650.1725 203.155 650.9325 203.57 ;
      RECT  651.3475 203.155 652.1075 203.57 ;
      RECT  652.5225 203.155 653.2825 203.57 ;
      RECT  653.6975 203.155 654.4575 203.57 ;
      RECT  654.8725 203.155 655.6325 203.57 ;
      RECT  656.0475 203.155 656.8075 203.57 ;
      RECT  657.2225 203.155 657.9825 203.57 ;
      RECT  658.3975 203.155 659.1575 203.57 ;
      RECT  659.5725 203.155 660.3325 203.57 ;
      RECT  660.7475 203.155 661.5075 203.57 ;
      RECT  661.9225 203.155 662.6825 203.57 ;
      RECT  663.0975 203.155 663.8575 203.57 ;
      RECT  664.2725 203.155 665.0325 203.57 ;
      RECT  665.4475 203.155 666.2075 203.57 ;
      RECT  666.6225 203.155 667.3825 203.57 ;
      RECT  667.7975 203.155 668.5575 203.57 ;
      RECT  668.9725 203.155 669.7325 203.57 ;
      RECT  670.1475 203.155 670.9075 203.57 ;
      RECT  671.3225 203.155 672.0825 203.57 ;
      RECT  672.4975 203.155 673.2575 203.57 ;
      RECT  673.6725 203.155 674.4325 203.57 ;
      RECT  674.8475 203.155 675.6075 203.57 ;
      RECT  676.0225 203.155 676.7825 203.57 ;
      RECT  677.1975 203.155 677.9575 203.57 ;
      RECT  678.3725 203.155 679.1325 203.57 ;
      RECT  679.5475 203.155 680.3075 203.57 ;
      RECT  680.7225 203.155 681.4825 203.57 ;
      RECT  681.8975 203.155 682.6575 203.57 ;
      RECT  683.0725 203.155 683.8325 203.57 ;
      RECT  684.2475 203.155 685.0075 203.57 ;
      RECT  685.4225 203.155 686.1825 203.57 ;
      RECT  686.5975 203.155 687.3575 203.57 ;
      RECT  687.7725 203.155 688.5325 203.57 ;
      RECT  688.9475 203.155 689.7075 203.57 ;
      RECT  690.1225 203.155 690.8825 203.57 ;
      RECT  691.2975 203.155 692.0575 203.57 ;
      RECT  692.4725 203.155 693.2325 203.57 ;
      RECT  693.6475 203.155 694.4075 203.57 ;
      RECT  694.8225 203.155 695.5825 203.57 ;
      RECT  695.9975 203.155 696.7575 203.57 ;
      RECT  697.1725 203.155 697.9325 203.57 ;
      RECT  698.3475 203.155 699.1075 203.57 ;
      RECT  699.5225 203.155 700.2825 203.57 ;
      RECT  700.6975 203.155 701.4575 203.57 ;
      RECT  701.8725 203.155 702.6325 203.57 ;
      RECT  703.0475 203.155 703.8075 203.57 ;
      RECT  704.2225 203.155 704.9825 203.57 ;
      RECT  705.3975 203.155 706.1575 203.57 ;
      RECT  706.5725 203.155 707.3325 203.57 ;
      RECT  707.7475 203.155 708.5075 203.57 ;
      RECT  708.9225 203.155 709.6825 203.57 ;
      RECT  710.0975 203.155 710.8575 203.57 ;
      RECT  711.2725 203.155 712.0325 203.57 ;
      RECT  712.4475 203.155 713.2075 203.57 ;
      RECT  713.6225 203.155 714.3825 203.57 ;
      RECT  714.7975 203.155 715.5575 203.57 ;
      RECT  715.9725 203.155 716.7325 203.57 ;
      RECT  717.1475 203.155 717.9075 203.57 ;
      RECT  718.3225 203.155 719.0825 203.57 ;
      RECT  719.4975 203.155 720.2575 203.57 ;
      RECT  720.6725 203.155 721.4325 203.57 ;
      RECT  721.8475 203.155 722.6075 203.57 ;
      RECT  723.0225 203.155 723.7825 203.57 ;
      RECT  724.1975 203.155 724.9575 203.57 ;
      RECT  725.3725 203.155 726.1325 203.57 ;
      RECT  726.5475 203.155 727.3075 203.57 ;
      RECT  727.7225 203.155 728.4825 203.57 ;
      RECT  728.8975 203.155 729.6575 203.57 ;
      RECT  730.0725 203.155 730.8325 203.57 ;
      RECT  731.2475 203.155 732.0075 203.57 ;
      RECT  732.4225 203.155 733.1825 203.57 ;
      RECT  733.5975 203.155 734.3575 203.57 ;
      RECT  734.7725 203.155 735.5325 203.57 ;
      RECT  735.9475 203.155 736.7075 203.57 ;
      RECT  737.1225 203.155 737.8825 203.57 ;
      RECT  738.2975 203.155 739.0575 203.57 ;
      RECT  739.4725 203.155 740.2325 203.57 ;
      RECT  740.6475 203.155 741.4075 203.57 ;
      RECT  741.8225 203.155 742.5825 203.57 ;
      RECT  742.9975 203.155 743.7575 203.57 ;
      RECT  744.1725 203.155 744.9325 203.57 ;
      RECT  745.3475 203.155 746.1075 203.57 ;
      RECT  746.5225 203.155 747.2825 203.57 ;
      RECT  747.6975 203.155 748.4575 203.57 ;
      RECT  748.8725 203.155 749.6325 203.57 ;
      RECT  750.0475 203.155 750.8075 203.57 ;
      RECT  751.2225 203.155 751.9825 203.57 ;
      RECT  752.3975 203.155 753.1575 203.57 ;
      RECT  753.5725 203.155 754.3325 203.57 ;
      RECT  754.7475 203.155 755.5075 203.57 ;
      RECT  755.9225 203.155 756.6825 203.57 ;
      RECT  757.0975 203.155 757.8575 203.57 ;
      RECT  758.2725 203.155 759.0325 203.57 ;
      RECT  759.4475 203.155 760.2075 203.57 ;
      RECT  760.6225 203.155 801.085 203.57 ;
      RECT  0.14 1.26 1.26 2.24 ;
      RECT  0.14 2.24 1.26 4.0975 ;
      RECT  1.26 2.24 125.925 4.0975 ;
      RECT  125.925 2.24 126.34 4.0975 ;
      RECT  126.34 2.24 1592.08 4.0975 ;
      RECT  1592.08 1.26 1593.2 2.24 ;
      RECT  1592.08 2.24 1593.2 4.0975 ;
      RECT  125.925 4.5125 126.34 212.1 ;
      RECT  0.14 122.7075 1.26 212.1 ;
      RECT  0.14 212.1 1.26 213.08 ;
      RECT  1.26 122.7075 120.205 212.1 ;
      RECT  120.62 122.7075 125.925 212.1 ;
      RECT  120.205 135.3175 120.62 212.1 ;
      RECT  801.085 96.5775 801.5 212.1 ;
      RECT  801.5 210.2775 918.185 212.1 ;
      RECT  918.185 210.2775 918.6 212.1 ;
      RECT  918.6 210.2775 1592.08 212.1 ;
      RECT  1592.08 210.2775 1593.2 212.1 ;
      RECT  1592.08 212.1 1593.2 213.08 ;
      RECT  126.34 203.57 159.7825 212.1 ;
      RECT  159.7825 203.57 160.1975 212.1 ;
      RECT  160.1975 203.57 801.085 212.1 ;
      RECT  0.14 0.84 1.26 1.26 ;
      RECT  1.26 0.84 125.925 1.26 ;
      RECT  125.925 0.84 126.34 1.26 ;
      RECT  126.34 0.84 1592.08 1.26 ;
      RECT  1592.08 0.84 1593.2 1.26 ;
      RECT  125.925 213.08 126.34 213.5 ;
      RECT  0.14 213.08 1.26 213.5 ;
      RECT  1.26 213.08 120.205 213.5 ;
      RECT  120.62 213.08 125.925 213.5 ;
      RECT  120.205 213.08 120.62 213.5 ;
      RECT  801.085 213.08 801.5 213.5 ;
      RECT  801.5 213.08 918.185 213.5 ;
      RECT  918.185 213.08 918.6 213.5 ;
      RECT  918.6 213.08 1592.08 213.5 ;
      RECT  1592.08 213.08 1593.2 213.5 ;
      RECT  126.34 213.08 159.7825 213.5 ;
      RECT  159.7825 213.08 160.1975 213.5 ;
      RECT  160.1975 213.08 801.085 213.5 ;
   LAYER  metal4 ;
      RECT  1.12 0.14 2.38 1.12 ;
      RECT  1.12 213.22 2.38 214.2 ;
      RECT  2.38 1.12 1590.96 213.22 ;
      RECT  2.38 0.14 1592.36 1.12 ;
      RECT  2.38 213.22 1592.36 214.2 ;
      RECT  1592.22 1.12 1592.36 213.22 ;
      RECT  0.98 0.14 1.12 1.12 ;
      RECT  0.98 1.12 1.12 213.22 ;
      RECT  0.98 213.22 1.12 214.2 ;
   END
END    freepdk45_sram_1w1r_64x512
END    LIBRARY
