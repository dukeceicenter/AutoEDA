../macros/freepdk45_sram_1w1r_128x124_31/freepdk45_sram_1w1r_128x124_31.lef