../macros/freepdk45_sram_1rw0r_64x44_22/freepdk45_sram_1rw0r_64x44_22.lef