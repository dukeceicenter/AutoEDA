../macros/freepdk45_sram_1rw0r_512x64/freepdk45_sram_1rw0r_512x64.lef