VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_27x96_32
   CLASS BLOCK ;
   SIZE 317.615 BY 89.11 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.27 1.105 43.405 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.13 1.105 46.265 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.99 1.105 49.125 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.85 1.105 51.985 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.71 1.105 54.845 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.57 1.105 57.705 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.43 1.105 60.565 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.29 1.105 63.425 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.15 1.105 66.285 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.01 1.105 69.145 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.87 1.105 72.005 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.73 1.105 74.865 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.59 1.105 77.725 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.45 1.105 80.585 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.31 1.105 83.445 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.17 1.105 86.305 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.03 1.105 89.165 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.89 1.105 92.025 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.75 1.105 94.885 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.61 1.105 97.745 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.47 1.105 100.605 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.33 1.105 103.465 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.19 1.105 106.325 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.05 1.105 109.185 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.91 1.105 112.045 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.77 1.105 114.905 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.63 1.105 117.765 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.49 1.105 120.625 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.35 1.105 123.485 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.21 1.105 126.345 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.07 1.105 129.205 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.93 1.105 132.065 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.79 1.105 134.925 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.65 1.105 137.785 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.51 1.105 140.645 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.37 1.105 143.505 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.23 1.105 146.365 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.09 1.105 149.225 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.95 1.105 152.085 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.81 1.105 154.945 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.67 1.105 157.805 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.53 1.105 160.665 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.39 1.105 163.525 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.25 1.105 166.385 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.11 1.105 169.245 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.97 1.105 172.105 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.83 1.105 174.965 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.69 1.105 177.825 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.55 1.105 180.685 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.41 1.105 183.545 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.27 1.105 186.405 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.13 1.105 189.265 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.99 1.105 192.125 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.85 1.105 194.985 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.71 1.105 197.845 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.57 1.105 200.705 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.43 1.105 203.565 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.29 1.105 206.425 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.15 1.105 209.285 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.01 1.105 212.145 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.87 1.105 215.005 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.73 1.105 217.865 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.59 1.105 220.725 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.45 1.105 223.585 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.31 1.105 226.445 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.17 1.105 229.305 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.03 1.105 232.165 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.89 1.105 235.025 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.75 1.105 237.885 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.61 1.105 240.745 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.47 1.105 243.605 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.33 1.105 246.465 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.19 1.105 249.325 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.05 1.105 252.185 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.91 1.105 255.045 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.77 1.105 257.905 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.63 1.105 260.765 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.49 1.105 263.625 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.35 1.105 266.485 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.21 1.105 269.345 1.24 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.07 1.105 272.205 1.24 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.93 1.105 275.065 1.24 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.79 1.105 277.925 1.24 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.65 1.105 280.785 1.24 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.51 1.105 283.645 1.24 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.37 1.105 286.505 1.24 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.23 1.105 289.365 1.24 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.09 1.105 292.225 1.24 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.95 1.105 295.085 1.24 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.81 1.105 297.945 1.24 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.67 1.105 300.805 1.24 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.53 1.105 303.665 1.24 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.39 1.105 306.525 1.24 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.25 1.105 309.385 1.24 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.11 1.105 312.245 1.24 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.97 1.105 315.105 1.24 ;
      END
   END din0[95]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.97 52.6225 29.105 52.7575 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.97 55.3525 29.105 55.4875 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.97 57.5625 29.105 57.6975 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.97 60.2925 29.105 60.4275 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.97 62.5025 29.105 62.6375 ;
      END
   END addr0[4]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.86 29.4825 185.995 29.6175 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.86 26.7525 185.995 26.8875 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.86 24.5425 185.995 24.6775 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.86 21.8125 185.995 21.9475 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.86 19.6025 185.995 19.7375 ;
      END
   END addr1[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 11.0225 0.42 11.1575 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.685 87.8675 214.82 88.0025 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 11.1075 6.3825 11.2425 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.5825 87.7825 208.7175 87.9175 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.69 1.105 34.825 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.55 1.105 37.685 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.41 1.105 40.545 1.24 ;
      END
   END wmask0[2]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.9525 81.1575 51.0875 81.2925 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.1275 81.1575 52.2625 81.2925 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.3025 81.1575 53.4375 81.2925 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.4775 81.1575 54.6125 81.2925 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.6525 81.1575 55.7875 81.2925 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.8275 81.1575 56.9625 81.2925 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.0025 81.1575 58.1375 81.2925 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.1775 81.1575 59.3125 81.2925 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.3525 81.1575 60.4875 81.2925 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.5275 81.1575 61.6625 81.2925 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.7025 81.1575 62.8375 81.2925 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.8775 81.1575 64.0125 81.2925 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.0525 81.1575 65.1875 81.2925 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.2275 81.1575 66.3625 81.2925 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.4025 81.1575 67.5375 81.2925 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.5775 81.1575 68.7125 81.2925 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.7525 81.1575 69.8875 81.2925 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.9275 81.1575 71.0625 81.2925 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.1025 81.1575 72.2375 81.2925 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.2775 81.1575 73.4125 81.2925 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.4525 81.1575 74.5875 81.2925 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.6275 81.1575 75.7625 81.2925 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.8025 81.1575 76.9375 81.2925 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.9775 81.1575 78.1125 81.2925 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.1525 81.1575 79.2875 81.2925 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.3275 81.1575 80.4625 81.2925 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.5025 81.1575 81.6375 81.2925 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.6775 81.1575 82.8125 81.2925 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.8525 81.1575 83.9875 81.2925 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.0275 81.1575 85.1625 81.2925 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.2025 81.1575 86.3375 81.2925 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.3775 81.1575 87.5125 81.2925 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.5525 81.1575 88.6875 81.2925 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.7275 81.1575 89.8625 81.2925 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.9025 81.1575 91.0375 81.2925 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.0775 81.1575 92.2125 81.2925 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.2525 81.1575 93.3875 81.2925 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.4275 81.1575 94.5625 81.2925 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.6025 81.1575 95.7375 81.2925 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.7775 81.1575 96.9125 81.2925 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.9525 81.1575 98.0875 81.2925 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.1275 81.1575 99.2625 81.2925 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.3025 81.1575 100.4375 81.2925 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.4775 81.1575 101.6125 81.2925 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.6525 81.1575 102.7875 81.2925 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.8275 81.1575 103.9625 81.2925 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.0025 81.1575 105.1375 81.2925 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.1775 81.1575 106.3125 81.2925 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.3525 81.1575 107.4875 81.2925 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.5275 81.1575 108.6625 81.2925 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.7025 81.1575 109.8375 81.2925 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.8775 81.1575 111.0125 81.2925 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.0525 81.1575 112.1875 81.2925 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.2275 81.1575 113.3625 81.2925 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.4025 81.1575 114.5375 81.2925 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.5775 81.1575 115.7125 81.2925 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.7525 81.1575 116.8875 81.2925 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.9275 81.1575 118.0625 81.2925 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.1025 81.1575 119.2375 81.2925 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.2775 81.1575 120.4125 81.2925 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.4525 81.1575 121.5875 81.2925 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.6275 81.1575 122.7625 81.2925 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.8025 81.1575 123.9375 81.2925 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.9775 81.1575 125.1125 81.2925 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.1525 81.1575 126.2875 81.2925 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.3275 81.1575 127.4625 81.2925 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.5025 81.1575 128.6375 81.2925 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.6775 81.1575 129.8125 81.2925 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.8525 81.1575 130.9875 81.2925 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.0275 81.1575 132.1625 81.2925 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.2025 81.1575 133.3375 81.2925 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.3775 81.1575 134.5125 81.2925 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.5525 81.1575 135.6875 81.2925 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.7275 81.1575 136.8625 81.2925 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.9025 81.1575 138.0375 81.2925 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.0775 81.1575 139.2125 81.2925 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.2525 81.1575 140.3875 81.2925 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.4275 81.1575 141.5625 81.2925 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.6025 81.1575 142.7375 81.2925 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.7775 81.1575 143.9125 81.2925 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.9525 81.1575 145.0875 81.2925 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.1275 81.1575 146.2625 81.2925 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.3025 81.1575 147.4375 81.2925 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.4775 81.1575 148.6125 81.2925 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.6525 81.1575 149.7875 81.2925 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.8275 81.1575 150.9625 81.2925 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.0025 81.1575 152.1375 81.2925 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.1775 81.1575 153.3125 81.2925 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.3525 81.1575 154.4875 81.2925 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.5275 81.1575 155.6625 81.2925 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.7025 81.1575 156.8375 81.2925 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.8775 81.1575 158.0125 81.2925 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.0525 81.1575 159.1875 81.2925 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.2275 81.1575 160.3625 81.2925 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.4025 81.1575 161.5375 81.2925 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.5775 81.1575 162.7125 81.2925 ;
      END
   END dout1[95]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  46.62 30.585 46.76 71.1225 ;
         LAYER metal3 ;
         RECT  88.7475 2.47 88.8825 2.605 ;
         LAYER metal3 ;
         RECT  54.4275 2.47 54.5625 2.605 ;
         LAYER metal3 ;
         RECT  163.7175 20.3175 163.8525 20.4525 ;
         LAYER metal4 ;
         RECT  40.62 30.585 40.76 71.16 ;
         LAYER metal3 ;
         RECT  65.8675 2.47 66.0025 2.605 ;
         LAYER metal3 ;
         RECT  47.7675 21.285 163.3825 21.355 ;
         LAYER metal4 ;
         RECT  47.7 27.415 47.84 74.01 ;
         LAYER metal3 ;
         RECT  157.3875 2.47 157.5225 2.605 ;
         LAYER metal4 ;
         RECT  214.2775 56.86 214.4175 79.2625 ;
         LAYER metal3 ;
         RECT  203.1475 2.47 203.2825 2.605 ;
         LAYER metal3 ;
         RECT  260.3475 2.47 260.4825 2.605 ;
         LAYER metal3 ;
         RECT  47.7675 26.72 163.8525 26.79 ;
         LAYER metal3 ;
         RECT  46.6225 29.0925 46.7575 29.2275 ;
         LAYER metal3 ;
         RECT  168.8275 2.47 168.9625 2.605 ;
         LAYER metal3 ;
         RECT  271.7875 2.47 271.9225 2.605 ;
         LAYER metal4 ;
         RECT  183.42 76.62 183.56 86.64 ;
         LAYER metal3 ;
         RECT  41.24 29.88 41.375 30.015 ;
         LAYER metal3 ;
         RECT  47.7675 78.6025 163.3825 78.6725 ;
         LAYER metal3 ;
         RECT  168.0125 72.4475 168.1475 72.5825 ;
         LAYER metal4 ;
         RECT  174.01 30.585 174.15 71.16 ;
         LAYER metal4 ;
         RECT  28.685 51.515 28.825 64.07 ;
         LAYER metal4 ;
         RECT  31.405 12.385 31.545 27.345 ;
         LAYER metal4 ;
         RECT  186.14 18.17 186.28 30.725 ;
         LAYER metal4 ;
         RECT  166.93 27.415 167.07 74.01 ;
         LAYER metal3 ;
         RECT  134.5075 2.47 134.6425 2.605 ;
         LAYER metal3 ;
         RECT  294.6675 2.47 294.8025 2.605 ;
         LAYER metal3 ;
         RECT  100.1875 2.47 100.3225 2.605 ;
         LAYER metal3 ;
         RECT  35.0675 44.0425 35.2025 44.1775 ;
         LAYER metal3 ;
         RECT  111.6275 2.47 111.7625 2.605 ;
         LAYER metal3 ;
         RECT  42.9875 2.47 43.1225 2.605 ;
         LAYER metal4 ;
         RECT  168.01 30.585 168.15 71.1225 ;
         LAYER metal3 ;
         RECT  2.425 12.3875 2.56 12.5225 ;
         LAYER metal4 ;
         RECT  0.6875 19.7625 0.8275 42.165 ;
         LAYER metal3 ;
         RECT  35.0675 41.0525 35.2025 41.1875 ;
         LAYER metal3 ;
         RECT  35.0675 50.0225 35.2025 50.1575 ;
         LAYER metal3 ;
         RECT  191.7075 2.47 191.8425 2.605 ;
         LAYER metal3 ;
         RECT  179.2225 35.0725 179.3575 35.2075 ;
         LAYER metal3 ;
         RECT  283.2275 2.47 283.3625 2.605 ;
         LAYER metal3 ;
         RECT  212.545 86.5025 212.68 86.6375 ;
         LAYER metal3 ;
         RECT  173.395 71.66 173.53 71.795 ;
         LAYER metal3 ;
         RECT  237.4675 2.47 237.6025 2.605 ;
         LAYER metal3 ;
         RECT  226.0275 2.47 226.1625 2.605 ;
         LAYER metal3 ;
         RECT  145.9475 2.47 146.0825 2.605 ;
         LAYER metal3 ;
         RECT  180.2675 2.47 180.4025 2.605 ;
         LAYER metal3 ;
         RECT  35.4125 32.0825 35.5475 32.2175 ;
         LAYER metal3 ;
         RECT  123.0675 2.47 123.2025 2.605 ;
         LAYER metal3 ;
         RECT  47.6325 20.3175 47.7675 20.4525 ;
         LAYER metal3 ;
         RECT  35.4125 35.0725 35.5475 35.2075 ;
         LAYER metal3 ;
         RECT  306.1075 2.47 306.2425 2.605 ;
         LAYER metal3 ;
         RECT  35.0675 47.0325 35.2025 47.1675 ;
         LAYER metal3 ;
         RECT  34.4075 2.47 34.5425 2.605 ;
         LAYER metal3 ;
         RECT  179.2225 32.0825 179.3575 32.2175 ;
         LAYER metal3 ;
         RECT  214.5875 2.47 214.7225 2.605 ;
         LAYER metal3 ;
         RECT  77.3075 2.47 77.4425 2.605 ;
         LAYER metal3 ;
         RECT  248.9075 2.47 249.0425 2.605 ;
         LAYER metal3 ;
         RECT  179.5675 50.0225 179.7025 50.1575 ;
         LAYER metal3 ;
         RECT  179.5675 41.0525 179.7025 41.1875 ;
         LAYER metal3 ;
         RECT  179.5675 44.0425 179.7025 44.1775 ;
         LAYER metal3 ;
         RECT  179.5675 47.0325 179.7025 47.1675 ;
         LAYER metal3 ;
         RECT  47.7675 74.705 165.0275 74.775 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  212.215 56.8275 212.355 79.23 ;
         LAYER metal3 ;
         RECT  68.7275 0.0 68.8625 0.135 ;
         LAYER metal4 ;
         RECT  173.45 30.5525 173.59 71.09 ;
         LAYER metal3 ;
         RECT  181.375 48.5275 181.51 48.6625 ;
         LAYER metal3 ;
         RECT  308.9675 0.0 309.1025 0.135 ;
         LAYER metal3 ;
         RECT  194.5675 0.0 194.7025 0.135 ;
         LAYER metal3 ;
         RECT  57.2875 0.0 57.4225 0.135 ;
         LAYER metal3 ;
         RECT  163.7175 18.4975 163.8525 18.6325 ;
         LAYER metal3 ;
         RECT  212.545 88.9725 212.68 89.1075 ;
         LAYER metal3 ;
         RECT  206.0075 0.0 206.1425 0.135 ;
         LAYER metal3 ;
         RECT  33.885 36.5675 34.02 36.7025 ;
         LAYER metal3 ;
         RECT  228.8875 0.0 229.0225 0.135 ;
         LAYER metal3 ;
         RECT  91.6075 0.0 91.7425 0.135 ;
         LAYER metal3 ;
         RECT  2.425 9.9175 2.56 10.0525 ;
         LAYER metal4 ;
         RECT  208.72 74.15 208.86 89.11 ;
         LAYER metal3 ;
         RECT  33.26 51.5175 33.395 51.6525 ;
         LAYER metal3 ;
         RECT  180.75 33.5775 180.885 33.7125 ;
         LAYER metal3 ;
         RECT  114.4875 0.0 114.6225 0.135 ;
         LAYER metal4 ;
         RECT  166.47 27.415 166.61 74.01 ;
         LAYER metal4 ;
         RECT  41.18 30.5525 41.32 71.09 ;
         LAYER metal3 ;
         RECT  181.375 39.5575 181.51 39.6925 ;
         LAYER metal3 ;
         RECT  47.7675 76.71 163.4175 76.78 ;
         LAYER metal3 ;
         RECT  148.8075 0.0 148.9425 0.135 ;
         LAYER metal4 ;
         RECT  31.545 51.45 31.685 64.005 ;
         LAYER metal3 ;
         RECT  125.9275 0.0 126.0625 0.135 ;
         LAYER metal3 ;
         RECT  297.5275 0.0 297.6625 0.135 ;
         LAYER metal4 ;
         RECT  48.16 27.415 48.3 74.01 ;
         LAYER metal3 ;
         RECT  274.6475 0.0 274.7825 0.135 ;
         LAYER metal3 ;
         RECT  137.3675 0.0 137.5025 0.135 ;
         LAYER metal4 ;
         RECT  2.75 19.795 2.89 42.1975 ;
         LAYER metal3 ;
         RECT  286.0875 0.0 286.2225 0.135 ;
         LAYER metal3 ;
         RECT  33.26 39.5575 33.395 39.6925 ;
         LAYER metal4 ;
         RECT  39.03 30.5525 39.17 71.16 ;
         LAYER metal4 ;
         RECT  6.105 9.915 6.245 24.875 ;
         LAYER metal3 ;
         RECT  33.26 42.5475 33.395 42.6825 ;
         LAYER metal3 ;
         RECT  183.1275 0.0 183.2625 0.135 ;
         LAYER metal3 ;
         RECT  33.885 33.5775 34.02 33.7125 ;
         LAYER metal3 ;
         RECT  180.75 30.5875 180.885 30.7225 ;
         LAYER metal3 ;
         RECT  263.2075 0.0 263.3425 0.135 ;
         LAYER metal3 ;
         RECT  103.0475 0.0 103.1825 0.135 ;
         LAYER metal3 ;
         RECT  181.375 51.5175 181.51 51.6525 ;
         LAYER metal3 ;
         RECT  80.1675 0.0 80.3025 0.135 ;
         LAYER metal3 ;
         RECT  33.26 48.5275 33.395 48.6625 ;
         LAYER metal3 ;
         RECT  180.75 36.5675 180.885 36.7025 ;
         LAYER metal3 ;
         RECT  181.375 45.5375 181.51 45.6725 ;
         LAYER metal4 ;
         RECT  183.28 18.235 183.42 30.79 ;
         LAYER metal3 ;
         RECT  181.375 42.5475 181.51 42.6825 ;
         LAYER metal3 ;
         RECT  45.8475 0.0 45.9825 0.135 ;
         LAYER metal3 ;
         RECT  251.7675 0.0 251.9025 0.135 ;
         LAYER metal3 ;
         RECT  240.3275 0.0 240.4625 0.135 ;
         LAYER metal3 ;
         RECT  171.6875 0.0 171.8225 0.135 ;
         LAYER metal3 ;
         RECT  160.2475 0.0 160.3825 0.135 ;
         LAYER metal4 ;
         RECT  175.6 30.5525 175.74 71.16 ;
         LAYER metal3 ;
         RECT  33.26 45.5375 33.395 45.6725 ;
         LAYER metal3 ;
         RECT  33.885 30.5875 34.02 30.7225 ;
         LAYER metal3 ;
         RECT  217.4475 0.0 217.5825 0.135 ;
         LAYER metal3 ;
         RECT  47.7675 23.335 163.3825 23.405 ;
         LAYER metal3 ;
         RECT  47.6325 18.4975 47.7675 18.6325 ;
         LAYER metal3 ;
         RECT  37.2675 0.0 37.4025 0.135 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 317.475 88.97 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 317.475 88.97 ;
   LAYER  metal3 ;
      RECT  43.13 0.14 43.545 0.965 ;
      RECT  43.545 0.965 45.99 1.38 ;
      RECT  46.405 0.965 48.85 1.38 ;
      RECT  49.265 0.965 51.71 1.38 ;
      RECT  52.125 0.965 54.57 1.38 ;
      RECT  54.985 0.965 57.43 1.38 ;
      RECT  57.845 0.965 60.29 1.38 ;
      RECT  60.705 0.965 63.15 1.38 ;
      RECT  63.565 0.965 66.01 1.38 ;
      RECT  66.425 0.965 68.87 1.38 ;
      RECT  69.285 0.965 71.73 1.38 ;
      RECT  72.145 0.965 74.59 1.38 ;
      RECT  75.005 0.965 77.45 1.38 ;
      RECT  77.865 0.965 80.31 1.38 ;
      RECT  80.725 0.965 83.17 1.38 ;
      RECT  83.585 0.965 86.03 1.38 ;
      RECT  86.445 0.965 88.89 1.38 ;
      RECT  89.305 0.965 91.75 1.38 ;
      RECT  92.165 0.965 94.61 1.38 ;
      RECT  95.025 0.965 97.47 1.38 ;
      RECT  97.885 0.965 100.33 1.38 ;
      RECT  100.745 0.965 103.19 1.38 ;
      RECT  103.605 0.965 106.05 1.38 ;
      RECT  106.465 0.965 108.91 1.38 ;
      RECT  109.325 0.965 111.77 1.38 ;
      RECT  112.185 0.965 114.63 1.38 ;
      RECT  115.045 0.965 117.49 1.38 ;
      RECT  117.905 0.965 120.35 1.38 ;
      RECT  120.765 0.965 123.21 1.38 ;
      RECT  123.625 0.965 126.07 1.38 ;
      RECT  126.485 0.965 128.93 1.38 ;
      RECT  129.345 0.965 131.79 1.38 ;
      RECT  132.205 0.965 134.65 1.38 ;
      RECT  135.065 0.965 137.51 1.38 ;
      RECT  137.925 0.965 140.37 1.38 ;
      RECT  140.785 0.965 143.23 1.38 ;
      RECT  143.645 0.965 146.09 1.38 ;
      RECT  146.505 0.965 148.95 1.38 ;
      RECT  149.365 0.965 151.81 1.38 ;
      RECT  152.225 0.965 154.67 1.38 ;
      RECT  155.085 0.965 157.53 1.38 ;
      RECT  157.945 0.965 160.39 1.38 ;
      RECT  160.805 0.965 163.25 1.38 ;
      RECT  163.665 0.965 166.11 1.38 ;
      RECT  166.525 0.965 168.97 1.38 ;
      RECT  169.385 0.965 171.83 1.38 ;
      RECT  172.245 0.965 174.69 1.38 ;
      RECT  175.105 0.965 177.55 1.38 ;
      RECT  177.965 0.965 180.41 1.38 ;
      RECT  180.825 0.965 183.27 1.38 ;
      RECT  183.685 0.965 186.13 1.38 ;
      RECT  186.545 0.965 188.99 1.38 ;
      RECT  189.405 0.965 191.85 1.38 ;
      RECT  192.265 0.965 194.71 1.38 ;
      RECT  195.125 0.965 197.57 1.38 ;
      RECT  197.985 0.965 200.43 1.38 ;
      RECT  200.845 0.965 203.29 1.38 ;
      RECT  203.705 0.965 206.15 1.38 ;
      RECT  206.565 0.965 209.01 1.38 ;
      RECT  209.425 0.965 211.87 1.38 ;
      RECT  212.285 0.965 214.73 1.38 ;
      RECT  215.145 0.965 217.59 1.38 ;
      RECT  218.005 0.965 220.45 1.38 ;
      RECT  220.865 0.965 223.31 1.38 ;
      RECT  223.725 0.965 226.17 1.38 ;
      RECT  226.585 0.965 229.03 1.38 ;
      RECT  229.445 0.965 231.89 1.38 ;
      RECT  232.305 0.965 234.75 1.38 ;
      RECT  235.165 0.965 237.61 1.38 ;
      RECT  238.025 0.965 240.47 1.38 ;
      RECT  240.885 0.965 243.33 1.38 ;
      RECT  243.745 0.965 246.19 1.38 ;
      RECT  246.605 0.965 249.05 1.38 ;
      RECT  249.465 0.965 251.91 1.38 ;
      RECT  252.325 0.965 254.77 1.38 ;
      RECT  255.185 0.965 257.63 1.38 ;
      RECT  258.045 0.965 260.49 1.38 ;
      RECT  260.905 0.965 263.35 1.38 ;
      RECT  263.765 0.965 266.21 1.38 ;
      RECT  266.625 0.965 269.07 1.38 ;
      RECT  269.485 0.965 271.93 1.38 ;
      RECT  272.345 0.965 274.79 1.38 ;
      RECT  275.205 0.965 277.65 1.38 ;
      RECT  278.065 0.965 280.51 1.38 ;
      RECT  280.925 0.965 283.37 1.38 ;
      RECT  283.785 0.965 286.23 1.38 ;
      RECT  286.645 0.965 289.09 1.38 ;
      RECT  289.505 0.965 291.95 1.38 ;
      RECT  292.365 0.965 294.81 1.38 ;
      RECT  295.225 0.965 297.67 1.38 ;
      RECT  298.085 0.965 300.53 1.38 ;
      RECT  300.945 0.965 303.39 1.38 ;
      RECT  303.805 0.965 306.25 1.38 ;
      RECT  306.665 0.965 309.11 1.38 ;
      RECT  309.525 0.965 311.97 1.38 ;
      RECT  312.385 0.965 314.83 1.38 ;
      RECT  315.245 0.965 317.475 1.38 ;
      RECT  0.14 52.4825 28.83 52.8975 ;
      RECT  0.14 52.8975 28.83 88.97 ;
      RECT  28.83 1.38 29.245 52.4825 ;
      RECT  29.245 52.4825 43.13 52.8975 ;
      RECT  29.245 52.8975 43.13 88.97 ;
      RECT  28.83 52.8975 29.245 55.2125 ;
      RECT  28.83 55.6275 29.245 57.4225 ;
      RECT  28.83 57.8375 29.245 60.1525 ;
      RECT  28.83 60.5675 29.245 62.3625 ;
      RECT  28.83 62.7775 29.245 88.97 ;
      RECT  185.72 29.7575 186.135 88.97 ;
      RECT  186.135 29.3425 317.475 29.7575 ;
      RECT  185.72 27.0275 186.135 29.3425 ;
      RECT  185.72 24.8175 186.135 26.6125 ;
      RECT  185.72 22.0875 186.135 24.4025 ;
      RECT  185.72 1.38 186.135 19.4625 ;
      RECT  185.72 19.8775 186.135 21.6725 ;
      RECT  0.14 1.38 0.145 10.8825 ;
      RECT  0.14 10.8825 0.145 11.2975 ;
      RECT  0.14 11.2975 0.145 52.4825 ;
      RECT  0.145 1.38 0.56 10.8825 ;
      RECT  0.145 11.2975 0.56 52.4825 ;
      RECT  214.545 29.7575 214.96 87.7275 ;
      RECT  214.545 88.1425 214.96 88.97 ;
      RECT  214.96 29.7575 317.475 87.7275 ;
      RECT  214.96 87.7275 317.475 88.1425 ;
      RECT  214.96 88.1425 317.475 88.97 ;
      RECT  0.56 10.8825 6.1075 10.9675 ;
      RECT  0.56 10.9675 6.1075 11.2975 ;
      RECT  6.1075 10.8825 6.5225 10.9675 ;
      RECT  6.5225 10.8825 28.83 10.9675 ;
      RECT  6.5225 10.9675 28.83 11.2975 ;
      RECT  0.56 11.2975 6.1075 11.3825 ;
      RECT  6.1075 11.3825 6.5225 52.4825 ;
      RECT  6.5225 11.2975 28.83 11.3825 ;
      RECT  6.5225 11.3825 28.83 52.4825 ;
      RECT  186.135 29.7575 208.4425 87.6425 ;
      RECT  186.135 87.6425 208.4425 87.7275 ;
      RECT  208.4425 29.7575 208.8575 87.6425 ;
      RECT  208.8575 87.6425 214.545 87.7275 ;
      RECT  186.135 87.7275 208.4425 88.0575 ;
      RECT  186.135 88.0575 208.4425 88.1425 ;
      RECT  208.4425 88.0575 208.8575 88.1425 ;
      RECT  208.8575 87.7275 214.545 88.0575 ;
      RECT  208.8575 88.0575 214.545 88.1425 ;
      RECT  0.14 0.965 34.55 1.38 ;
      RECT  34.965 0.965 37.41 1.38 ;
      RECT  37.825 0.965 40.27 1.38 ;
      RECT  40.685 0.965 43.13 1.38 ;
      RECT  43.545 81.0175 50.8125 81.4325 ;
      RECT  43.545 81.4325 50.8125 88.97 ;
      RECT  50.8125 81.4325 51.2275 88.97 ;
      RECT  51.2275 81.4325 185.72 88.97 ;
      RECT  51.2275 81.0175 51.9875 81.4325 ;
      RECT  52.4025 81.0175 53.1625 81.4325 ;
      RECT  53.5775 81.0175 54.3375 81.4325 ;
      RECT  54.7525 81.0175 55.5125 81.4325 ;
      RECT  55.9275 81.0175 56.6875 81.4325 ;
      RECT  57.1025 81.0175 57.8625 81.4325 ;
      RECT  58.2775 81.0175 59.0375 81.4325 ;
      RECT  59.4525 81.0175 60.2125 81.4325 ;
      RECT  60.6275 81.0175 61.3875 81.4325 ;
      RECT  61.8025 81.0175 62.5625 81.4325 ;
      RECT  62.9775 81.0175 63.7375 81.4325 ;
      RECT  64.1525 81.0175 64.9125 81.4325 ;
      RECT  65.3275 81.0175 66.0875 81.4325 ;
      RECT  66.5025 81.0175 67.2625 81.4325 ;
      RECT  67.6775 81.0175 68.4375 81.4325 ;
      RECT  68.8525 81.0175 69.6125 81.4325 ;
      RECT  70.0275 81.0175 70.7875 81.4325 ;
      RECT  71.2025 81.0175 71.9625 81.4325 ;
      RECT  72.3775 81.0175 73.1375 81.4325 ;
      RECT  73.5525 81.0175 74.3125 81.4325 ;
      RECT  74.7275 81.0175 75.4875 81.4325 ;
      RECT  75.9025 81.0175 76.6625 81.4325 ;
      RECT  77.0775 81.0175 77.8375 81.4325 ;
      RECT  78.2525 81.0175 79.0125 81.4325 ;
      RECT  79.4275 81.0175 80.1875 81.4325 ;
      RECT  80.6025 81.0175 81.3625 81.4325 ;
      RECT  81.7775 81.0175 82.5375 81.4325 ;
      RECT  82.9525 81.0175 83.7125 81.4325 ;
      RECT  84.1275 81.0175 84.8875 81.4325 ;
      RECT  85.3025 81.0175 86.0625 81.4325 ;
      RECT  86.4775 81.0175 87.2375 81.4325 ;
      RECT  87.6525 81.0175 88.4125 81.4325 ;
      RECT  88.8275 81.0175 89.5875 81.4325 ;
      RECT  90.0025 81.0175 90.7625 81.4325 ;
      RECT  91.1775 81.0175 91.9375 81.4325 ;
      RECT  92.3525 81.0175 93.1125 81.4325 ;
      RECT  93.5275 81.0175 94.2875 81.4325 ;
      RECT  94.7025 81.0175 95.4625 81.4325 ;
      RECT  95.8775 81.0175 96.6375 81.4325 ;
      RECT  97.0525 81.0175 97.8125 81.4325 ;
      RECT  98.2275 81.0175 98.9875 81.4325 ;
      RECT  99.4025 81.0175 100.1625 81.4325 ;
      RECT  100.5775 81.0175 101.3375 81.4325 ;
      RECT  101.7525 81.0175 102.5125 81.4325 ;
      RECT  102.9275 81.0175 103.6875 81.4325 ;
      RECT  104.1025 81.0175 104.8625 81.4325 ;
      RECT  105.2775 81.0175 106.0375 81.4325 ;
      RECT  106.4525 81.0175 107.2125 81.4325 ;
      RECT  107.6275 81.0175 108.3875 81.4325 ;
      RECT  108.8025 81.0175 109.5625 81.4325 ;
      RECT  109.9775 81.0175 110.7375 81.4325 ;
      RECT  111.1525 81.0175 111.9125 81.4325 ;
      RECT  112.3275 81.0175 113.0875 81.4325 ;
      RECT  113.5025 81.0175 114.2625 81.4325 ;
      RECT  114.6775 81.0175 115.4375 81.4325 ;
      RECT  115.8525 81.0175 116.6125 81.4325 ;
      RECT  117.0275 81.0175 117.7875 81.4325 ;
      RECT  118.2025 81.0175 118.9625 81.4325 ;
      RECT  119.3775 81.0175 120.1375 81.4325 ;
      RECT  120.5525 81.0175 121.3125 81.4325 ;
      RECT  121.7275 81.0175 122.4875 81.4325 ;
      RECT  122.9025 81.0175 123.6625 81.4325 ;
      RECT  124.0775 81.0175 124.8375 81.4325 ;
      RECT  125.2525 81.0175 126.0125 81.4325 ;
      RECT  126.4275 81.0175 127.1875 81.4325 ;
      RECT  127.6025 81.0175 128.3625 81.4325 ;
      RECT  128.7775 81.0175 129.5375 81.4325 ;
      RECT  129.9525 81.0175 130.7125 81.4325 ;
      RECT  131.1275 81.0175 131.8875 81.4325 ;
      RECT  132.3025 81.0175 133.0625 81.4325 ;
      RECT  133.4775 81.0175 134.2375 81.4325 ;
      RECT  134.6525 81.0175 135.4125 81.4325 ;
      RECT  135.8275 81.0175 136.5875 81.4325 ;
      RECT  137.0025 81.0175 137.7625 81.4325 ;
      RECT  138.1775 81.0175 138.9375 81.4325 ;
      RECT  139.3525 81.0175 140.1125 81.4325 ;
      RECT  140.5275 81.0175 141.2875 81.4325 ;
      RECT  141.7025 81.0175 142.4625 81.4325 ;
      RECT  142.8775 81.0175 143.6375 81.4325 ;
      RECT  144.0525 81.0175 144.8125 81.4325 ;
      RECT  145.2275 81.0175 145.9875 81.4325 ;
      RECT  146.4025 81.0175 147.1625 81.4325 ;
      RECT  147.5775 81.0175 148.3375 81.4325 ;
      RECT  148.7525 81.0175 149.5125 81.4325 ;
      RECT  149.9275 81.0175 150.6875 81.4325 ;
      RECT  151.1025 81.0175 151.8625 81.4325 ;
      RECT  152.2775 81.0175 153.0375 81.4325 ;
      RECT  153.4525 81.0175 154.2125 81.4325 ;
      RECT  154.6275 81.0175 155.3875 81.4325 ;
      RECT  155.8025 81.0175 156.5625 81.4325 ;
      RECT  156.9775 81.0175 157.7375 81.4325 ;
      RECT  158.1525 81.0175 158.9125 81.4325 ;
      RECT  159.3275 81.0175 160.0875 81.4325 ;
      RECT  160.5025 81.0175 161.2625 81.4325 ;
      RECT  161.6775 81.0175 162.4375 81.4325 ;
      RECT  162.8525 81.0175 185.72 81.4325 ;
      RECT  43.545 1.38 88.6075 2.33 ;
      RECT  88.6075 1.38 89.0225 2.33 ;
      RECT  89.0225 1.38 185.72 2.33 ;
      RECT  43.545 2.33 54.2875 2.745 ;
      RECT  89.0225 2.745 163.5775 20.1775 ;
      RECT  89.0225 20.1775 163.5775 20.5925 ;
      RECT  163.9925 2.745 185.72 20.1775 ;
      RECT  163.9925 20.1775 185.72 20.5925 ;
      RECT  163.9925 20.5925 185.72 29.3425 ;
      RECT  54.7025 2.33 65.7275 2.745 ;
      RECT  43.545 21.145 47.6275 21.495 ;
      RECT  88.6075 2.745 89.0225 21.145 ;
      RECT  89.0225 20.5925 163.5225 21.145 ;
      RECT  163.5225 20.5925 163.5775 21.145 ;
      RECT  163.5225 21.145 163.5775 21.495 ;
      RECT  186.135 1.38 203.0075 2.33 ;
      RECT  186.135 2.745 203.0075 29.3425 ;
      RECT  203.0075 1.38 203.4225 2.33 ;
      RECT  203.0075 2.745 203.4225 29.3425 ;
      RECT  203.4225 1.38 317.475 2.33 ;
      RECT  203.4225 2.745 317.475 29.3425 ;
      RECT  163.5775 20.5925 163.9925 26.58 ;
      RECT  163.5775 26.93 163.9925 29.3425 ;
      RECT  47.6275 26.93 88.6075 29.3425 ;
      RECT  88.6075 26.93 89.0225 29.3425 ;
      RECT  89.0225 26.93 163.5225 29.3425 ;
      RECT  163.5225 21.495 163.5775 26.58 ;
      RECT  163.5225 26.93 163.5775 29.3425 ;
      RECT  43.545 29.3425 46.4825 29.3675 ;
      RECT  43.545 29.3675 46.4825 29.7575 ;
      RECT  46.4825 29.3675 46.8975 29.7575 ;
      RECT  46.8975 29.3425 185.72 29.3675 ;
      RECT  46.8975 29.3675 185.72 29.7575 ;
      RECT  43.545 21.495 46.4825 28.9525 ;
      RECT  43.545 28.9525 46.4825 29.3425 ;
      RECT  46.4825 21.495 46.8975 28.9525 ;
      RECT  46.8975 21.495 47.6275 28.9525 ;
      RECT  46.8975 28.9525 47.6275 29.3425 ;
      RECT  157.6625 2.33 168.6875 2.745 ;
      RECT  260.6225 2.33 271.6475 2.745 ;
      RECT  29.245 29.74 41.1 30.155 ;
      RECT  41.1 1.38 41.515 29.74 ;
      RECT  41.1 30.155 41.515 52.4825 ;
      RECT  41.515 29.74 43.13 30.155 ;
      RECT  41.515 30.155 43.13 52.4825 ;
      RECT  43.545 29.7575 47.6275 78.4625 ;
      RECT  43.545 78.4625 47.6275 78.8125 ;
      RECT  43.545 78.8125 47.6275 81.0175 ;
      RECT  47.6275 78.8125 50.8125 81.0175 ;
      RECT  50.8125 78.8125 51.2275 81.0175 ;
      RECT  51.2275 78.8125 163.5225 81.0175 ;
      RECT  163.5225 78.4625 185.72 78.8125 ;
      RECT  163.5225 78.8125 185.72 81.0175 ;
      RECT  163.5225 29.7575 167.8725 72.3075 ;
      RECT  163.5225 72.3075 167.8725 72.7225 ;
      RECT  167.8725 29.7575 168.2875 72.3075 ;
      RECT  167.8725 72.7225 168.2875 78.4625 ;
      RECT  168.2875 72.3075 185.72 72.7225 ;
      RECT  168.2875 72.7225 185.72 78.4625 ;
      RECT  89.0225 2.33 100.0475 2.745 ;
      RECT  29.245 43.9025 34.9275 44.3175 ;
      RECT  35.3425 43.9025 41.1 44.3175 ;
      RECT  35.3425 44.3175 41.1 52.4825 ;
      RECT  100.4625 2.33 111.4875 2.745 ;
      RECT  43.13 1.38 43.2625 2.33 ;
      RECT  43.13 2.745 43.2625 88.97 ;
      RECT  43.2625 1.38 43.545 2.33 ;
      RECT  43.2625 2.33 43.545 2.745 ;
      RECT  43.2625 2.745 43.545 88.97 ;
      RECT  41.515 1.38 42.8475 2.33 ;
      RECT  41.515 2.33 42.8475 2.745 ;
      RECT  41.515 2.745 42.8475 29.74 ;
      RECT  42.8475 1.38 43.13 2.33 ;
      RECT  42.8475 2.745 43.13 29.74 ;
      RECT  0.56 11.3825 2.285 12.2475 ;
      RECT  0.56 12.2475 2.285 12.6625 ;
      RECT  0.56 12.6625 2.285 52.4825 ;
      RECT  2.285 11.3825 2.7 12.2475 ;
      RECT  2.285 12.6625 2.7 52.4825 ;
      RECT  2.7 11.3825 6.1075 12.2475 ;
      RECT  2.7 12.2475 6.1075 12.6625 ;
      RECT  2.7 12.6625 6.1075 52.4825 ;
      RECT  34.9275 41.3275 35.3425 43.9025 ;
      RECT  34.9275 50.2975 35.3425 52.4825 ;
      RECT  186.135 2.33 191.5675 2.745 ;
      RECT  191.9825 2.33 203.0075 2.745 ;
      RECT  168.2875 29.7575 179.0825 34.9325 ;
      RECT  168.2875 34.9325 179.0825 35.3475 ;
      RECT  179.4975 34.9325 185.72 35.3475 ;
      RECT  272.0625 2.33 283.0875 2.745 ;
      RECT  283.5025 2.33 294.5275 2.745 ;
      RECT  208.8575 29.7575 212.405 86.3625 ;
      RECT  208.8575 86.3625 212.405 86.7775 ;
      RECT  208.8575 86.7775 212.405 87.6425 ;
      RECT  212.405 29.7575 212.82 86.3625 ;
      RECT  212.405 86.7775 212.82 87.6425 ;
      RECT  212.82 29.7575 214.545 86.3625 ;
      RECT  212.82 86.3625 214.545 86.7775 ;
      RECT  212.82 86.7775 214.545 87.6425 ;
      RECT  168.2875 35.3475 173.255 71.52 ;
      RECT  168.2875 71.52 173.255 71.935 ;
      RECT  168.2875 71.935 173.255 72.3075 ;
      RECT  173.255 35.3475 173.67 71.52 ;
      RECT  173.255 71.935 173.67 72.3075 ;
      RECT  173.67 35.3475 179.0825 71.52 ;
      RECT  173.67 71.52 179.0825 71.935 ;
      RECT  173.67 71.935 179.0825 72.3075 ;
      RECT  226.3025 2.33 237.3275 2.745 ;
      RECT  134.7825 2.33 145.8075 2.745 ;
      RECT  146.2225 2.33 157.2475 2.745 ;
      RECT  169.1025 2.33 180.1275 2.745 ;
      RECT  180.5425 2.33 185.72 2.745 ;
      RECT  35.3425 30.155 35.6875 31.9425 ;
      RECT  35.6875 30.155 41.1 31.9425 ;
      RECT  35.6875 31.9425 41.1 32.3575 ;
      RECT  35.6875 32.3575 41.1 43.9025 ;
      RECT  34.9275 30.155 35.2725 31.9425 ;
      RECT  34.9275 31.9425 35.2725 32.3575 ;
      RECT  34.9275 32.3575 35.2725 40.9125 ;
      RECT  35.2725 30.155 35.3425 31.9425 ;
      RECT  111.9025 2.33 122.9275 2.745 ;
      RECT  123.3425 2.33 134.3675 2.745 ;
      RECT  43.545 2.745 47.4925 20.1775 ;
      RECT  43.545 20.1775 47.4925 20.5925 ;
      RECT  43.545 20.5925 47.4925 21.145 ;
      RECT  47.4925 20.5925 47.6275 21.145 ;
      RECT  47.6275 20.5925 47.9075 21.145 ;
      RECT  47.9075 2.745 88.6075 20.1775 ;
      RECT  47.9075 20.1775 88.6075 20.5925 ;
      RECT  47.9075 20.5925 88.6075 21.145 ;
      RECT  35.3425 32.3575 35.6875 34.9325 ;
      RECT  35.3425 35.3475 35.6875 43.9025 ;
      RECT  35.2725 32.3575 35.3425 34.9325 ;
      RECT  35.2725 35.3475 35.3425 40.9125 ;
      RECT  294.9425 2.33 305.9675 2.745 ;
      RECT  306.3825 2.33 317.475 2.745 ;
      RECT  34.9275 44.3175 35.3425 46.8925 ;
      RECT  34.9275 47.3075 35.3425 49.8825 ;
      RECT  29.245 1.38 34.2675 2.33 ;
      RECT  29.245 2.33 34.2675 2.745 ;
      RECT  29.245 2.745 34.2675 29.74 ;
      RECT  34.2675 1.38 34.6825 2.33 ;
      RECT  34.2675 2.745 34.6825 29.74 ;
      RECT  34.6825 1.38 41.1 2.33 ;
      RECT  34.6825 2.33 41.1 2.745 ;
      RECT  34.6825 2.745 41.1 29.74 ;
      RECT  179.0825 29.7575 179.4975 31.9425 ;
      RECT  179.0825 32.3575 179.4975 34.9325 ;
      RECT  203.4225 2.33 214.4475 2.745 ;
      RECT  214.8625 2.33 225.8875 2.745 ;
      RECT  66.1425 2.33 77.1675 2.745 ;
      RECT  77.5825 2.33 88.6075 2.745 ;
      RECT  237.7425 2.33 248.7675 2.745 ;
      RECT  249.1825 2.33 260.2075 2.745 ;
      RECT  179.0825 35.3475 179.4275 49.8825 ;
      RECT  179.0825 49.8825 179.4275 50.2975 ;
      RECT  179.0825 50.2975 179.4275 72.3075 ;
      RECT  179.4275 50.2975 179.4975 72.3075 ;
      RECT  179.4975 50.2975 179.8425 72.3075 ;
      RECT  179.8425 49.8825 185.72 50.2975 ;
      RECT  179.4275 35.3475 179.4975 40.9125 ;
      RECT  179.4975 35.3475 179.8425 40.9125 ;
      RECT  179.4275 41.3275 179.4975 43.9025 ;
      RECT  179.4975 41.3275 179.8425 43.9025 ;
      RECT  179.4275 44.3175 179.4975 46.8925 ;
      RECT  179.4275 47.3075 179.4975 49.8825 ;
      RECT  179.4975 44.3175 179.8425 46.8925 ;
      RECT  179.4975 47.3075 179.8425 49.8825 ;
      RECT  47.6275 29.7575 50.8125 74.565 ;
      RECT  50.8125 29.7575 51.2275 74.565 ;
      RECT  51.2275 29.7575 163.5225 74.565 ;
      RECT  163.5225 72.7225 165.1675 74.565 ;
      RECT  165.1675 72.7225 167.8725 74.565 ;
      RECT  165.1675 74.565 167.8725 74.915 ;
      RECT  165.1675 74.915 167.8725 78.4625 ;
      RECT  43.545 0.275 68.5875 0.965 ;
      RECT  68.5875 0.275 69.0025 0.965 ;
      RECT  69.0025 0.275 317.475 0.965 ;
      RECT  179.8425 48.3875 181.235 48.8025 ;
      RECT  179.8425 48.8025 181.235 49.8825 ;
      RECT  181.235 48.8025 181.65 49.8825 ;
      RECT  181.65 35.3475 185.72 48.3875 ;
      RECT  181.65 48.3875 185.72 48.8025 ;
      RECT  181.65 48.8025 185.72 49.8825 ;
      RECT  309.2425 0.14 317.475 0.275 ;
      RECT  57.5625 0.14 68.5875 0.275 ;
      RECT  163.5775 2.745 163.9925 18.3575 ;
      RECT  163.5775 18.7725 163.9925 20.1775 ;
      RECT  186.135 88.1425 212.405 88.8325 ;
      RECT  186.135 88.8325 212.405 88.97 ;
      RECT  212.405 88.1425 212.82 88.8325 ;
      RECT  212.82 88.1425 214.545 88.8325 ;
      RECT  212.82 88.8325 214.545 88.97 ;
      RECT  194.8425 0.14 205.8675 0.275 ;
      RECT  29.245 30.155 33.745 36.4275 ;
      RECT  29.245 36.4275 33.745 36.8425 ;
      RECT  33.745 36.8425 34.16 43.9025 ;
      RECT  34.16 30.155 34.9275 36.4275 ;
      RECT  34.16 36.4275 34.9275 36.8425 ;
      RECT  34.16 36.8425 34.9275 43.9025 ;
      RECT  0.56 1.38 2.285 9.7775 ;
      RECT  0.56 9.7775 2.285 10.1925 ;
      RECT  0.56 10.1925 2.285 10.8825 ;
      RECT  2.285 1.38 2.7 9.7775 ;
      RECT  2.285 10.1925 2.7 10.8825 ;
      RECT  2.7 1.38 28.83 9.7775 ;
      RECT  2.7 9.7775 28.83 10.1925 ;
      RECT  2.7 10.1925 28.83 10.8825 ;
      RECT  29.245 44.3175 33.12 51.3775 ;
      RECT  29.245 51.3775 33.12 51.7925 ;
      RECT  29.245 51.7925 33.12 52.4825 ;
      RECT  33.12 51.7925 33.535 52.4825 ;
      RECT  33.535 44.3175 34.9275 51.3775 ;
      RECT  33.535 51.3775 34.9275 51.7925 ;
      RECT  33.535 51.7925 34.9275 52.4825 ;
      RECT  179.4975 29.7575 180.61 33.4375 ;
      RECT  179.4975 33.4375 180.61 33.8525 ;
      RECT  179.4975 33.8525 180.61 34.9325 ;
      RECT  180.61 33.8525 181.025 34.9325 ;
      RECT  181.025 29.7575 185.72 33.4375 ;
      RECT  181.025 33.4375 185.72 33.8525 ;
      RECT  181.025 33.8525 185.72 34.9325 ;
      RECT  181.235 35.3475 181.65 39.4175 ;
      RECT  47.6275 74.915 50.8125 76.57 ;
      RECT  47.6275 76.92 50.8125 78.4625 ;
      RECT  50.8125 74.915 51.2275 76.57 ;
      RECT  50.8125 76.92 51.2275 78.4625 ;
      RECT  51.2275 74.915 163.5225 76.57 ;
      RECT  51.2275 76.92 163.5225 78.4625 ;
      RECT  163.5225 74.915 163.5575 76.57 ;
      RECT  163.5225 76.92 163.5575 78.4625 ;
      RECT  163.5575 74.915 165.1675 76.57 ;
      RECT  163.5575 76.57 165.1675 76.92 ;
      RECT  163.5575 76.92 165.1675 78.4625 ;
      RECT  114.7625 0.14 125.7875 0.275 ;
      RECT  297.8025 0.14 308.8275 0.275 ;
      RECT  126.2025 0.14 137.2275 0.275 ;
      RECT  137.6425 0.14 148.6675 0.275 ;
      RECT  274.9225 0.14 285.9475 0.275 ;
      RECT  286.3625 0.14 297.3875 0.275 ;
      RECT  29.245 36.8425 33.12 39.4175 ;
      RECT  29.245 39.4175 33.12 39.8325 ;
      RECT  29.245 39.8325 33.12 43.9025 ;
      RECT  33.12 36.8425 33.535 39.4175 ;
      RECT  33.535 36.8425 33.745 39.4175 ;
      RECT  33.535 39.4175 33.745 39.8325 ;
      RECT  33.535 39.8325 33.745 43.9025 ;
      RECT  33.12 39.8325 33.535 42.4075 ;
      RECT  33.12 42.8225 33.535 43.9025 ;
      RECT  183.4025 0.14 194.4275 0.275 ;
      RECT  33.745 33.8525 34.16 36.4275 ;
      RECT  180.61 29.7575 181.025 30.4475 ;
      RECT  180.61 30.8625 181.025 33.4375 ;
      RECT  263.4825 0.14 274.5075 0.275 ;
      RECT  91.8825 0.14 102.9075 0.275 ;
      RECT  103.3225 0.14 114.3475 0.275 ;
      RECT  179.8425 50.2975 181.235 51.3775 ;
      RECT  179.8425 51.3775 181.235 51.7925 ;
      RECT  179.8425 51.7925 181.235 72.3075 ;
      RECT  181.235 50.2975 181.65 51.3775 ;
      RECT  181.235 51.7925 181.65 72.3075 ;
      RECT  181.65 50.2975 185.72 51.3775 ;
      RECT  181.65 51.3775 185.72 51.7925 ;
      RECT  181.65 51.7925 185.72 72.3075 ;
      RECT  69.0025 0.14 80.0275 0.275 ;
      RECT  80.4425 0.14 91.4675 0.275 ;
      RECT  33.12 48.8025 33.535 51.3775 ;
      RECT  179.8425 35.3475 180.61 36.4275 ;
      RECT  179.8425 36.4275 180.61 36.8425 ;
      RECT  179.8425 36.8425 180.61 48.3875 ;
      RECT  180.61 35.3475 181.025 36.4275 ;
      RECT  180.61 36.8425 181.025 48.3875 ;
      RECT  181.025 35.3475 181.235 36.4275 ;
      RECT  181.025 36.4275 181.235 36.8425 ;
      RECT  181.025 36.8425 181.235 48.3875 ;
      RECT  181.235 45.8125 181.65 48.3875 ;
      RECT  181.235 39.8325 181.65 42.4075 ;
      RECT  181.235 42.8225 181.65 45.3975 ;
      RECT  43.545 0.14 45.7075 0.275 ;
      RECT  46.1225 0.14 57.1475 0.275 ;
      RECT  252.0425 0.14 263.0675 0.275 ;
      RECT  229.1625 0.14 240.1875 0.275 ;
      RECT  240.6025 0.14 251.6275 0.275 ;
      RECT  171.9625 0.14 182.9875 0.275 ;
      RECT  149.0825 0.14 160.1075 0.275 ;
      RECT  160.5225 0.14 171.5475 0.275 ;
      RECT  33.12 44.3175 33.535 45.3975 ;
      RECT  33.12 45.8125 33.535 48.3875 ;
      RECT  33.745 30.155 34.16 30.4475 ;
      RECT  33.745 30.8625 34.16 33.4375 ;
      RECT  206.2825 0.14 217.3075 0.275 ;
      RECT  217.7225 0.14 228.7475 0.275 ;
      RECT  47.6275 21.495 88.6075 23.195 ;
      RECT  47.6275 23.545 88.6075 26.58 ;
      RECT  88.6075 21.495 89.0225 23.195 ;
      RECT  88.6075 23.545 89.0225 26.58 ;
      RECT  89.0225 21.495 163.5225 23.195 ;
      RECT  89.0225 23.545 163.5225 26.58 ;
      RECT  47.4925 2.745 47.6275 18.3575 ;
      RECT  47.4925 18.7725 47.6275 20.1775 ;
      RECT  47.6275 2.745 47.9075 18.3575 ;
      RECT  47.6275 18.7725 47.9075 20.1775 ;
      RECT  0.14 0.14 37.1275 0.275 ;
      RECT  0.14 0.275 37.1275 0.965 ;
      RECT  37.1275 0.275 37.5425 0.965 ;
      RECT  37.5425 0.14 43.13 0.275 ;
      RECT  37.5425 0.275 43.13 0.965 ;
   LAYER  metal4 ;
      RECT  46.34 0.14 47.04 30.305 ;
      RECT  46.34 71.4025 47.04 88.97 ;
      RECT  0.14 71.44 40.34 88.97 ;
      RECT  40.34 71.44 41.04 88.97 ;
      RECT  41.04 71.4025 46.34 71.44 ;
      RECT  41.04 71.44 46.34 88.97 ;
      RECT  47.04 0.14 47.42 27.135 ;
      RECT  47.04 27.135 47.42 30.305 ;
      RECT  47.42 0.14 48.12 27.135 ;
      RECT  47.04 30.305 47.42 71.4025 ;
      RECT  47.04 71.4025 47.42 74.29 ;
      RECT  47.04 74.29 47.42 88.97 ;
      RECT  47.42 74.29 48.12 88.97 ;
      RECT  213.9975 30.305 214.6975 56.58 ;
      RECT  214.6975 30.305 317.475 56.58 ;
      RECT  214.6975 56.58 317.475 71.4025 ;
      RECT  214.6975 71.4025 317.475 74.29 ;
      RECT  213.9975 79.5425 214.6975 88.97 ;
      RECT  214.6975 74.29 317.475 79.5425 ;
      RECT  214.6975 79.5425 317.475 88.97 ;
      RECT  48.12 74.29 183.14 76.34 ;
      RECT  48.12 76.34 183.14 79.5425 ;
      RECT  183.14 74.29 183.84 76.34 ;
      RECT  48.12 79.5425 183.14 86.92 ;
      RECT  48.12 86.92 183.14 88.97 ;
      RECT  183.14 86.92 183.84 88.97 ;
      RECT  173.73 71.44 174.43 74.29 ;
      RECT  0.14 51.235 28.405 64.35 ;
      RECT  0.14 64.35 28.405 71.4025 ;
      RECT  28.405 30.305 29.105 51.235 ;
      RECT  28.405 64.35 29.105 71.4025 ;
      RECT  31.125 0.14 31.825 12.105 ;
      RECT  31.125 27.625 31.825 30.305 ;
      RECT  31.825 0.14 46.34 12.105 ;
      RECT  31.825 12.105 46.34 27.625 ;
      RECT  48.12 0.14 185.86 17.89 ;
      RECT  185.86 0.14 186.56 17.89 ;
      RECT  186.56 0.14 317.475 17.89 ;
      RECT  186.56 17.89 317.475 27.135 ;
      RECT  186.56 27.135 317.475 30.305 ;
      RECT  185.86 31.005 186.56 56.58 ;
      RECT  186.56 30.305 213.9975 31.005 ;
      RECT  167.35 71.4025 173.73 71.44 ;
      RECT  167.35 71.44 173.73 74.29 ;
      RECT  167.35 30.305 167.73 56.58 ;
      RECT  167.35 56.58 167.73 71.4025 ;
      RECT  0.14 30.305 0.4075 42.445 ;
      RECT  0.14 42.445 0.4075 51.235 ;
      RECT  0.4075 42.445 1.1075 51.235 ;
      RECT  0.14 12.105 0.4075 19.4825 ;
      RECT  0.14 19.4825 0.4075 27.625 ;
      RECT  0.4075 12.105 1.1075 19.4825 ;
      RECT  0.14 27.625 0.4075 30.305 ;
      RECT  212.635 74.29 213.9975 76.34 ;
      RECT  211.935 79.51 212.635 79.5425 ;
      RECT  212.635 76.34 213.9975 79.51 ;
      RECT  212.635 79.51 213.9975 79.5425 ;
      RECT  212.635 56.58 213.9975 71.4025 ;
      RECT  212.635 71.4025 213.9975 71.44 ;
      RECT  212.635 71.44 213.9975 74.29 ;
      RECT  186.56 31.005 211.935 56.5475 ;
      RECT  186.56 56.5475 211.935 56.58 ;
      RECT  211.935 31.005 212.635 56.5475 ;
      RECT  212.635 31.005 213.9975 56.5475 ;
      RECT  212.635 56.5475 213.9975 56.58 ;
      RECT  167.35 27.135 173.17 30.2725 ;
      RECT  167.35 30.2725 173.17 30.305 ;
      RECT  173.17 27.135 173.87 30.2725 ;
      RECT  168.43 30.305 173.17 56.58 ;
      RECT  168.43 56.58 173.17 71.37 ;
      RECT  168.43 71.37 173.17 71.4025 ;
      RECT  173.17 71.37 173.73 71.4025 ;
      RECT  183.84 79.5425 208.44 86.92 ;
      RECT  209.14 79.5425 213.9975 86.92 ;
      RECT  183.84 86.92 208.44 88.97 ;
      RECT  209.14 86.92 213.9975 88.97 ;
      RECT  183.84 74.29 208.44 76.34 ;
      RECT  209.14 74.29 211.935 76.34 ;
      RECT  183.84 76.34 208.44 79.51 ;
      RECT  209.14 76.34 211.935 79.51 ;
      RECT  183.84 79.51 208.44 79.5425 ;
      RECT  209.14 79.51 211.935 79.5425 ;
      RECT  174.43 71.44 208.44 73.87 ;
      RECT  174.43 73.87 208.44 74.29 ;
      RECT  208.44 71.44 209.14 73.87 ;
      RECT  209.14 71.44 211.935 73.87 ;
      RECT  209.14 73.87 211.935 74.29 ;
      RECT  41.04 71.37 41.6 71.4025 ;
      RECT  41.6 30.305 46.34 71.37 ;
      RECT  41.6 71.37 46.34 71.4025 ;
      RECT  31.825 27.625 40.9 30.2725 ;
      RECT  40.9 27.625 41.6 30.2725 ;
      RECT  41.6 27.625 46.34 30.2725 ;
      RECT  41.6 30.2725 46.34 30.305 ;
      RECT  29.105 30.305 31.265 51.17 ;
      RECT  29.105 51.17 31.265 51.235 ;
      RECT  31.265 30.305 31.965 51.17 ;
      RECT  29.105 51.235 31.265 64.285 ;
      RECT  29.105 64.285 31.265 64.35 ;
      RECT  31.265 64.285 31.965 64.35 ;
      RECT  48.58 30.305 166.19 56.58 ;
      RECT  48.58 56.58 166.19 71.4025 ;
      RECT  48.58 71.4025 166.19 71.44 ;
      RECT  48.58 71.44 166.19 74.29 ;
      RECT  48.58 27.135 166.19 30.305 ;
      RECT  1.1075 30.305 2.47 42.445 ;
      RECT  3.17 30.305 28.405 42.445 ;
      RECT  1.1075 42.445 2.47 42.4775 ;
      RECT  1.1075 42.4775 2.47 51.235 ;
      RECT  2.47 42.4775 3.17 51.235 ;
      RECT  3.17 42.445 28.405 42.4775 ;
      RECT  3.17 42.4775 28.405 51.235 ;
      RECT  1.1075 19.4825 2.47 19.515 ;
      RECT  1.1075 19.515 2.47 27.625 ;
      RECT  2.47 19.4825 3.17 19.515 ;
      RECT  1.1075 27.625 2.47 30.305 ;
      RECT  3.17 27.625 31.125 30.305 ;
      RECT  0.14 71.4025 38.75 71.44 ;
      RECT  39.45 71.4025 40.34 71.44 ;
      RECT  29.105 64.35 38.75 71.4025 ;
      RECT  39.45 64.35 40.34 71.4025 ;
      RECT  31.825 30.2725 38.75 30.305 ;
      RECT  39.45 30.2725 40.9 30.305 ;
      RECT  31.965 30.305 38.75 51.17 ;
      RECT  39.45 30.305 40.34 51.17 ;
      RECT  31.965 51.17 38.75 51.235 ;
      RECT  39.45 51.17 40.34 51.235 ;
      RECT  31.965 51.235 38.75 64.285 ;
      RECT  39.45 51.235 40.34 64.285 ;
      RECT  31.965 64.285 38.75 64.35 ;
      RECT  39.45 64.285 40.34 64.35 ;
      RECT  0.14 0.14 5.825 9.635 ;
      RECT  0.14 9.635 5.825 12.105 ;
      RECT  5.825 0.14 6.525 9.635 ;
      RECT  6.525 0.14 31.125 9.635 ;
      RECT  6.525 9.635 31.125 12.105 ;
      RECT  1.1075 12.105 5.825 19.4825 ;
      RECT  6.525 12.105 31.125 19.4825 ;
      RECT  3.17 19.4825 5.825 19.515 ;
      RECT  6.525 19.4825 31.125 19.515 ;
      RECT  3.17 19.515 5.825 25.155 ;
      RECT  3.17 25.155 5.825 27.625 ;
      RECT  5.825 25.155 6.525 27.625 ;
      RECT  6.525 19.515 31.125 25.155 ;
      RECT  6.525 25.155 31.125 27.625 ;
      RECT  48.12 17.89 183.0 17.955 ;
      RECT  48.12 17.955 183.0 27.135 ;
      RECT  183.0 17.89 183.7 17.955 ;
      RECT  183.7 17.89 185.86 17.955 ;
      RECT  183.7 17.955 185.86 27.135 ;
      RECT  183.7 30.305 185.86 31.005 ;
      RECT  183.0 31.07 183.7 56.58 ;
      RECT  183.7 31.005 185.86 31.07 ;
      RECT  183.7 31.07 185.86 56.58 ;
      RECT  173.87 27.135 183.0 30.2725 ;
      RECT  183.7 27.135 185.86 30.2725 ;
      RECT  183.7 30.2725 185.86 30.305 ;
      RECT  174.43 56.58 175.32 71.4025 ;
      RECT  176.02 56.58 211.935 71.4025 ;
      RECT  174.43 71.4025 175.32 71.44 ;
      RECT  176.02 71.4025 211.935 71.44 ;
      RECT  174.43 30.305 175.32 31.005 ;
      RECT  176.02 30.305 183.0 31.005 ;
      RECT  174.43 31.005 175.32 31.07 ;
      RECT  176.02 31.005 183.0 31.07 ;
      RECT  174.43 31.07 175.32 56.58 ;
      RECT  176.02 31.07 183.0 56.58 ;
      RECT  173.87 30.2725 175.32 30.305 ;
      RECT  176.02 30.2725 183.0 30.305 ;
   END
END    freepdk45_sram_1w1r_27x96_32
END    LIBRARY
