../macros/freepdk45_sram_1w1r_128x40/freepdk45_sram_1w1r_128x40.lef