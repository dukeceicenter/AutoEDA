/home/yl996/proj/mcp-eda-example/libraries/FreePDK45/OpenRAM/macros/freepdk45_sram_1w1r_28x128_32/freepdk45_sram_1w1r_28x128_32.lef