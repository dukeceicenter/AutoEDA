/home/yl996/proj/mcp-eda-example/libraries/FreePDK45/OpenRAM/macros/freepdk45_sram_1w1r_2048x8_2/freepdk45_sram_1w1r_2048x8_2.lef