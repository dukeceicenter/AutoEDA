../macros/freepdk45_sram_1rw0r_64x20_64/freepdk45_sram_1rw0r_64x20_64.lef