/home/yl996/proj/mcp-eda-example/libraries/FreePDK45/OpenRAM/macros/freepdk45_sram_1rw0r_256x64/freepdk45_sram_1rw0r_256x64.lef