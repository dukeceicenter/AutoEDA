../macros/freepdk45_sram_1w1r_128x44_11/freepdk45_sram_1w1r_128x44_11.lef