../macros/freepdk45_sram_1w1r_40x72/freepdk45_sram_1w1r_40x72.lef