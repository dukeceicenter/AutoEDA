../macros/freepdk45_sram_1w1r_256x4_1/freepdk45_sram_1w1r_256x4_1.lef