../macros/freepdk45_sram_1w1r_32x32_32/freepdk45_sram_1w1r_32x32_32.lef