VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1rw0r_64x160_20
   CLASS BLOCK ;
   SIZE 529.81 BY 143.4675 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.425 1.105 72.56 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.285 1.105 75.42 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.145 1.105 78.28 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.005 1.105 81.14 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.865 1.105 84.0 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.725 1.105 86.86 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.585 1.105 89.72 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.445 1.105 92.58 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.305 1.105 95.44 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.165 1.105 98.3 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.025 1.105 101.16 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.885 1.105 104.02 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.745 1.105 106.88 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.605 1.105 109.74 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.465 1.105 112.6 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.325 1.105 115.46 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.185 1.105 118.32 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.045 1.105 121.18 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.905 1.105 124.04 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.765 1.105 126.9 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.625 1.105 129.76 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.485 1.105 132.62 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.345 1.105 135.48 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.205 1.105 138.34 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.065 1.105 141.2 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.925 1.105 144.06 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.785 1.105 146.92 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.645 1.105 149.78 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.505 1.105 152.64 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.365 1.105 155.5 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.225 1.105 158.36 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.085 1.105 161.22 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.945 1.105 164.08 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.805 1.105 166.94 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.665 1.105 169.8 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.525 1.105 172.66 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.385 1.105 175.52 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.245 1.105 178.38 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.105 1.105 181.24 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.965 1.105 184.1 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.825 1.105 186.96 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.685 1.105 189.82 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.545 1.105 192.68 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.405 1.105 195.54 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.265 1.105 198.4 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.125 1.105 201.26 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.985 1.105 204.12 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.845 1.105 206.98 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.705 1.105 209.84 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.565 1.105 212.7 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.425 1.105 215.56 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.285 1.105 218.42 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.145 1.105 221.28 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.005 1.105 224.14 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.865 1.105 227.0 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.725 1.105 229.86 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.585 1.105 232.72 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.445 1.105 235.58 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.305 1.105 238.44 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.165 1.105 241.3 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.025 1.105 244.16 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.885 1.105 247.02 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.745 1.105 249.88 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.605 1.105 252.74 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.465 1.105 255.6 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.325 1.105 258.46 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.185 1.105 261.32 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.045 1.105 264.18 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.905 1.105 267.04 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.765 1.105 269.9 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.625 1.105 272.76 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.485 1.105 275.62 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.345 1.105 278.48 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.205 1.105 281.34 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.065 1.105 284.2 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.925 1.105 287.06 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.785 1.105 289.92 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.645 1.105 292.78 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.505 1.105 295.64 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.365 1.105 298.5 1.24 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.225 1.105 301.36 1.24 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.085 1.105 304.22 1.24 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.945 1.105 307.08 1.24 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.805 1.105 309.94 1.24 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.665 1.105 312.8 1.24 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.525 1.105 315.66 1.24 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.385 1.105 318.52 1.24 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.245 1.105 321.38 1.24 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.105 1.105 324.24 1.24 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.965 1.105 327.1 1.24 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.825 1.105 329.96 1.24 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.685 1.105 332.82 1.24 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.545 1.105 335.68 1.24 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.405 1.105 338.54 1.24 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.265 1.105 341.4 1.24 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.125 1.105 344.26 1.24 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.985 1.105 347.12 1.24 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.845 1.105 349.98 1.24 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.705 1.105 352.84 1.24 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.565 1.105 355.7 1.24 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.425 1.105 358.56 1.24 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.285 1.105 361.42 1.24 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.145 1.105 364.28 1.24 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.005 1.105 367.14 1.24 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.865 1.105 370.0 1.24 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.725 1.105 372.86 1.24 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.585 1.105 375.72 1.24 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.445 1.105 378.58 1.24 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.305 1.105 381.44 1.24 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.165 1.105 384.3 1.24 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  387.025 1.105 387.16 1.24 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.885 1.105 390.02 1.24 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.745 1.105 392.88 1.24 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.605 1.105 395.74 1.24 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.465 1.105 398.6 1.24 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.325 1.105 401.46 1.24 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.185 1.105 404.32 1.24 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.045 1.105 407.18 1.24 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.905 1.105 410.04 1.24 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.765 1.105 412.9 1.24 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.625 1.105 415.76 1.24 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.485 1.105 418.62 1.24 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.345 1.105 421.48 1.24 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.205 1.105 424.34 1.24 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.065 1.105 427.2 1.24 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.925 1.105 430.06 1.24 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.785 1.105 432.92 1.24 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.645 1.105 435.78 1.24 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.505 1.105 438.64 1.24 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.365 1.105 441.5 1.24 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.225 1.105 444.36 1.24 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.085 1.105 447.22 1.24 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.945 1.105 450.08 1.24 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.805 1.105 452.94 1.24 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.665 1.105 455.8 1.24 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.525 1.105 458.66 1.24 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.385 1.105 461.52 1.24 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.245 1.105 464.38 1.24 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.105 1.105 467.24 1.24 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.965 1.105 470.1 1.24 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.825 1.105 472.96 1.24 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.685 1.105 475.82 1.24 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.545 1.105 478.68 1.24 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.405 1.105 481.54 1.24 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.265 1.105 484.4 1.24 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.125 1.105 487.26 1.24 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.985 1.105 490.12 1.24 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.845 1.105 492.98 1.24 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.705 1.105 495.84 1.24 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.565 1.105 498.7 1.24 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.425 1.105 501.56 1.24 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.285 1.105 504.42 1.24 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.145 1.105 507.28 1.24 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.005 1.105 510.14 1.24 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.865 1.105 513.0 1.24 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.725 1.105 515.86 1.24 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.585 1.105 518.72 1.24 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.445 1.105 521.58 1.24 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  524.305 1.105 524.44 1.24 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.165 1.105 527.3 1.24 ;
      END
   END din0[159]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.825 77.4225 43.96 77.5575 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.825 80.1525 43.96 80.2875 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.825 82.3625 43.96 82.4975 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.825 85.0925 43.96 85.2275 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.825 87.3025 43.96 87.4375 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.825 90.0325 43.96 90.1675 ;
      END
   END addr0[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 32.7025 0.42 32.8375 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 35.4325 0.42 35.5675 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 32.7875 6.6625 32.9225 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.545 1.105 49.68 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.405 1.105 52.54 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.265 1.105 55.4 1.24 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.125 1.105 58.26 1.24 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.985 1.105 61.12 1.24 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.845 1.105 63.98 1.24 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.705 1.105 66.84 1.24 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.565 1.105 69.7 1.24 ;
      END
   END wmask0[7]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.7125 44.3525 68.8475 44.4875 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.4175 44.3525 69.5525 44.4875 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.1225 44.3525 70.2575 44.4875 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.8275 44.3525 70.9625 44.4875 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.5325 44.3525 71.6675 44.4875 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.2375 44.3525 72.3725 44.4875 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.9425 44.3525 73.0775 44.4875 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.6475 44.3525 73.7825 44.4875 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.3525 44.3525 74.4875 44.4875 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.0575 44.3525 75.1925 44.4875 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.7625 44.3525 75.8975 44.4875 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.4675 44.3525 76.6025 44.4875 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.1725 44.3525 77.3075 44.4875 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.8775 44.3525 78.0125 44.4875 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.5825 44.3525 78.7175 44.4875 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.2875 44.3525 79.4225 44.4875 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.9925 44.3525 80.1275 44.4875 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.6975 44.3525 80.8325 44.4875 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.4025 44.3525 81.5375 44.4875 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.1075 44.3525 82.2425 44.4875 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.8125 44.3525 82.9475 44.4875 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.5175 44.3525 83.6525 44.4875 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.2225 44.3525 84.3575 44.4875 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.9275 44.3525 85.0625 44.4875 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.6325 44.3525 85.7675 44.4875 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.3375 44.3525 86.4725 44.4875 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.0425 44.3525 87.1775 44.4875 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.7475 44.3525 87.8825 44.4875 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.4525 44.3525 88.5875 44.4875 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.1575 44.3525 89.2925 44.4875 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.8625 44.3525 89.9975 44.4875 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.5675 44.3525 90.7025 44.4875 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.2725 44.3525 91.4075 44.4875 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.9775 44.3525 92.1125 44.4875 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.6825 44.3525 92.8175 44.4875 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.3875 44.3525 93.5225 44.4875 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.0925 44.3525 94.2275 44.4875 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.7975 44.3525 94.9325 44.4875 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.5025 44.3525 95.6375 44.4875 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.2075 44.3525 96.3425 44.4875 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.9125 44.3525 97.0475 44.4875 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.6175 44.3525 97.7525 44.4875 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.3225 44.3525 98.4575 44.4875 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.0275 44.3525 99.1625 44.4875 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.7325 44.3525 99.8675 44.4875 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.4375 44.3525 100.5725 44.4875 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.1425 44.3525 101.2775 44.4875 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.8475 44.3525 101.9825 44.4875 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.5525 44.3525 102.6875 44.4875 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.2575 44.3525 103.3925 44.4875 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.9625 44.3525 104.0975 44.4875 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.6675 44.3525 104.8025 44.4875 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.3725 44.3525 105.5075 44.4875 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.0775 44.3525 106.2125 44.4875 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.7825 44.3525 106.9175 44.4875 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.4875 44.3525 107.6225 44.4875 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.1925 44.3525 108.3275 44.4875 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.8975 44.3525 109.0325 44.4875 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.6025 44.3525 109.7375 44.4875 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.3075 44.3525 110.4425 44.4875 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.0125 44.3525 111.1475 44.4875 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.7175 44.3525 111.8525 44.4875 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.4225 44.3525 112.5575 44.4875 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.1275 44.3525 113.2625 44.4875 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.8325 44.3525 113.9675 44.4875 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.5375 44.3525 114.6725 44.4875 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.2425 44.3525 115.3775 44.4875 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.9475 44.3525 116.0825 44.4875 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.6525 44.3525 116.7875 44.4875 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.3575 44.3525 117.4925 44.4875 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.0625 44.3525 118.1975 44.4875 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.7675 44.3525 118.9025 44.4875 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.4725 44.3525 119.6075 44.4875 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.1775 44.3525 120.3125 44.4875 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.8825 44.3525 121.0175 44.4875 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.5875 44.3525 121.7225 44.4875 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.2925 44.3525 122.4275 44.4875 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.9975 44.3525 123.1325 44.4875 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.7025 44.3525 123.8375 44.4875 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.4075 44.3525 124.5425 44.4875 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.1125 44.3525 125.2475 44.4875 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.8175 44.3525 125.9525 44.4875 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.5225 44.3525 126.6575 44.4875 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.2275 44.3525 127.3625 44.4875 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.9325 44.3525 128.0675 44.4875 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.6375 44.3525 128.7725 44.4875 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.3425 44.3525 129.4775 44.4875 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.0475 44.3525 130.1825 44.4875 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.7525 44.3525 130.8875 44.4875 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.4575 44.3525 131.5925 44.4875 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.1625 44.3525 132.2975 44.4875 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.8675 44.3525 133.0025 44.4875 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.5725 44.3525 133.7075 44.4875 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.2775 44.3525 134.4125 44.4875 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.9825 44.3525 135.1175 44.4875 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.6875 44.3525 135.8225 44.4875 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.3925 44.3525 136.5275 44.4875 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.0975 44.3525 137.2325 44.4875 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.8025 44.3525 137.9375 44.4875 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.5075 44.3525 138.6425 44.4875 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.2125 44.3525 139.3475 44.4875 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.9175 44.3525 140.0525 44.4875 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.6225 44.3525 140.7575 44.4875 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.3275 44.3525 141.4625 44.4875 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.0325 44.3525 142.1675 44.4875 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.7375 44.3525 142.8725 44.4875 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.4425 44.3525 143.5775 44.4875 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.1475 44.3525 144.2825 44.4875 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.8525 44.3525 144.9875 44.4875 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.5575 44.3525 145.6925 44.4875 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.2625 44.3525 146.3975 44.4875 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.9675 44.3525 147.1025 44.4875 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.6725 44.3525 147.8075 44.4875 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.3775 44.3525 148.5125 44.4875 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.0825 44.3525 149.2175 44.4875 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.7875 44.3525 149.9225 44.4875 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.4925 44.3525 150.6275 44.4875 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.1975 44.3525 151.3325 44.4875 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.9025 44.3525 152.0375 44.4875 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.6075 44.3525 152.7425 44.4875 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.3125 44.3525 153.4475 44.4875 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.0175 44.3525 154.1525 44.4875 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.7225 44.3525 154.8575 44.4875 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.4275 44.3525 155.5625 44.4875 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.1325 44.3525 156.2675 44.4875 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.8375 44.3525 156.9725 44.4875 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.5425 44.3525 157.6775 44.4875 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.2475 44.3525 158.3825 44.4875 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.9525 44.3525 159.0875 44.4875 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.6575 44.3525 159.7925 44.4875 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.3625 44.3525 160.4975 44.4875 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.0675 44.3525 161.2025 44.4875 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.7725 44.3525 161.9075 44.4875 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.4775 44.3525 162.6125 44.4875 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.1825 44.3525 163.3175 44.4875 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.8875 44.3525 164.0225 44.4875 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.5925 44.3525 164.7275 44.4875 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.2975 44.3525 165.4325 44.4875 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.0025 44.3525 166.1375 44.4875 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.7075 44.3525 166.8425 44.4875 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.4125 44.3525 167.5475 44.4875 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.1175 44.3525 168.2525 44.4875 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.8225 44.3525 168.9575 44.4875 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.5275 44.3525 169.6625 44.4875 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.2325 44.3525 170.3675 44.4875 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.9375 44.3525 171.0725 44.4875 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.6425 44.3525 171.7775 44.4875 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.3475 44.3525 172.4825 44.4875 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.0525 44.3525 173.1875 44.4875 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.7575 44.3525 173.8925 44.4875 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.4625 44.3525 174.5975 44.4875 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.1675 44.3525 175.3025 44.4875 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.8725 44.3525 176.0075 44.4875 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.5775 44.3525 176.7125 44.4875 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.2825 44.3525 177.4175 44.4875 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.9875 44.3525 178.1225 44.4875 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.6925 44.3525 178.8275 44.4875 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.3975 44.3525 179.5325 44.4875 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.1025 44.3525 180.2375 44.4875 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.8075 44.3525 180.9425 44.4875 ;
      END
   END dout0[159]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  49.2625 2.47 49.3975 2.605 ;
         LAYER metal3 ;
         RECT  66.4675 40.045 181.6125 40.115 ;
         LAYER metal3 ;
         RECT  95.0225 2.47 95.1575 2.605 ;
         LAYER metal3 ;
         RECT  381.0225 2.47 381.1575 2.605 ;
         LAYER metal3 ;
         RECT  495.4225 2.47 495.5575 2.605 ;
         LAYER metal3 ;
         RECT  518.3025 2.47 518.4375 2.605 ;
         LAYER metal3 ;
         RECT  175.1025 2.47 175.2375 2.605 ;
         LAYER metal3 ;
         RECT  66.3325 39.0775 66.4675 39.2125 ;
         LAYER metal3 ;
         RECT  506.8625 2.47 506.9975 2.605 ;
         LAYER metal3 ;
         RECT  266.6225 2.47 266.7575 2.605 ;
         LAYER metal3 ;
         RECT  312.3825 2.47 312.5175 2.605 ;
         LAYER metal3 ;
         RECT  197.9825 2.47 198.1175 2.605 ;
         LAYER metal3 ;
         RECT  472.5425 2.47 472.6775 2.605 ;
         LAYER metal4 ;
         RECT  55.195 54.475 55.335 142.045 ;
         LAYER metal3 ;
         RECT  117.9025 2.47 118.0375 2.605 ;
         LAYER metal3 ;
         RECT  300.9425 2.47 301.0775 2.605 ;
         LAYER metal3 ;
         RECT  186.5425 2.47 186.6775 2.605 ;
         LAYER metal3 ;
         RECT  140.7825 2.47 140.9175 2.605 ;
         LAYER metal3 ;
         RECT  220.8625 2.47 220.9975 2.605 ;
         LAYER metal3 ;
         RECT  65.3225 53.1125 65.4575 53.2475 ;
         LAYER metal3 ;
         RECT  181.4775 39.0775 181.6125 39.2125 ;
         LAYER metal3 ;
         RECT  403.9025 2.47 404.0375 2.605 ;
         LAYER metal4 ;
         RECT  46.26 34.065 46.4 49.025 ;
         LAYER metal3 ;
         RECT  278.0625 2.47 278.1975 2.605 ;
         LAYER metal3 ;
         RECT  209.4225 2.47 209.5575 2.605 ;
         LAYER metal3 ;
         RECT  483.9825 2.47 484.1175 2.605 ;
         LAYER metal3 ;
         RECT  243.7425 2.47 243.8775 2.605 ;
         LAYER metal3 ;
         RECT  49.6425 64.0325 49.7775 64.1675 ;
         LAYER metal3 ;
         RECT  66.4675 50.87 181.6125 50.94 ;
         LAYER metal3 ;
         RECT  49.6425 72.2225 49.7775 72.3575 ;
         LAYER metal3 ;
         RECT  426.7825 2.47 426.9175 2.605 ;
         LAYER metal3 ;
         RECT  55.815 53.77 55.95 53.905 ;
         LAYER metal3 ;
         RECT  323.8225 2.47 323.9575 2.605 ;
         LAYER metal3 ;
         RECT  346.7025 2.47 346.8375 2.605 ;
         LAYER metal3 ;
         RECT  392.4625 2.47 392.5975 2.605 ;
         LAYER metal3 ;
         RECT  438.2225 2.47 438.3575 2.605 ;
         LAYER metal4 ;
         RECT  0.0 31.595 0.14 36.675 ;
         LAYER metal3 ;
         RECT  129.3425 2.47 129.4775 2.605 ;
         LAYER metal3 ;
         RECT  232.3025 2.47 232.4375 2.605 ;
         LAYER metal3 ;
         RECT  369.5825 2.47 369.7175 2.605 ;
         LAYER metal3 ;
         RECT  358.1425 2.47 358.2775 2.605 ;
         LAYER metal3 ;
         RECT  49.6425 74.9525 49.7775 75.0875 ;
         LAYER metal4 ;
         RECT  43.54 76.315 43.68 91.275 ;
         LAYER metal3 ;
         RECT  163.6625 2.47 163.7975 2.605 ;
         LAYER metal3 ;
         RECT  255.1825 2.47 255.3175 2.605 ;
         LAYER metal3 ;
         RECT  289.5025 2.47 289.6375 2.605 ;
         LAYER metal3 ;
         RECT  72.1425 2.47 72.2775 2.605 ;
         LAYER metal3 ;
         RECT  49.6425 58.5725 49.7775 58.7075 ;
         LAYER metal3 ;
         RECT  415.3425 2.47 415.4775 2.605 ;
         LAYER metal4 ;
         RECT  65.32 54.475 65.46 141.975 ;
         LAYER metal3 ;
         RECT  83.5825 2.47 83.7175 2.605 ;
         LAYER metal4 ;
         RECT  183.045 51.565 183.185 143.27 ;
         LAYER metal4 ;
         RECT  66.4 51.565 66.54 143.27 ;
         LAYER metal3 ;
         RECT  49.6425 66.7625 49.7775 66.8975 ;
         LAYER metal3 ;
         RECT  335.2625 2.47 335.3975 2.605 ;
         LAYER metal3 ;
         RECT  461.1025 2.47 461.2375 2.605 ;
         LAYER metal3 ;
         RECT  49.6425 55.8425 49.7775 55.9775 ;
         LAYER metal3 ;
         RECT  66.4675 46.9725 181.6125 47.0425 ;
         LAYER metal3 ;
         RECT  60.7025 2.47 60.8375 2.605 ;
         LAYER metal3 ;
         RECT  449.6625 2.47 449.7975 2.605 ;
         LAYER metal3 ;
         RECT  106.4625 2.47 106.5975 2.605 ;
         LAYER metal3 ;
         RECT  152.2225 2.47 152.3575 2.605 ;
         LAYER metal4 ;
         RECT  0.6875 41.4425 0.8275 63.845 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  181.4775 37.2575 181.6125 37.3925 ;
         LAYER metal3 ;
         RECT  452.5225 0.0 452.6575 0.135 ;
         LAYER metal3 ;
         RECT  66.4675 42.095 181.6125 42.165 ;
         LAYER metal3 ;
         RECT  269.4825 0.0 269.6175 0.135 ;
         LAYER metal3 ;
         RECT  441.0825 0.0 441.2175 0.135 ;
         LAYER metal3 ;
         RECT  48.115 68.1275 48.25 68.2625 ;
         LAYER metal3 ;
         RECT  521.1625 0.0 521.2975 0.135 ;
         LAYER metal3 ;
         RECT  48.115 62.6675 48.25 62.8025 ;
         LAYER metal3 ;
         RECT  155.0825 0.0 155.2175 0.135 ;
         LAYER metal3 ;
         RECT  48.115 57.2075 48.25 57.3425 ;
         LAYER metal3 ;
         RECT  338.1225 0.0 338.2575 0.135 ;
         LAYER metal3 ;
         RECT  143.6425 0.0 143.7775 0.135 ;
         LAYER metal3 ;
         RECT  48.115 65.3975 48.25 65.5325 ;
         LAYER metal3 ;
         RECT  212.2825 0.0 212.4175 0.135 ;
         LAYER metal3 ;
         RECT  372.4425 0.0 372.5775 0.135 ;
         LAYER metal4 ;
         RECT  4.845 31.53 4.985 36.74 ;
         LAYER metal3 ;
         RECT  132.2025 0.0 132.3375 0.135 ;
         LAYER metal3 ;
         RECT  509.7225 0.0 509.8575 0.135 ;
         LAYER metal4 ;
         RECT  55.755 54.4425 55.895 142.0075 ;
         LAYER metal3 ;
         RECT  86.4425 0.0 86.5775 0.135 ;
         LAYER metal3 ;
         RECT  75.0025 0.0 75.1375 0.135 ;
         LAYER metal3 ;
         RECT  486.8425 0.0 486.9775 0.135 ;
         LAYER metal3 ;
         RECT  48.115 73.5875 48.25 73.7225 ;
         LAYER metal3 ;
         RECT  292.3625 0.0 292.4975 0.135 ;
         LAYER metal3 ;
         RECT  361.0025 0.0 361.1375 0.135 ;
         LAYER metal3 ;
         RECT  315.2425 0.0 315.3775 0.135 ;
         LAYER metal3 ;
         RECT  418.2025 0.0 418.3375 0.135 ;
         LAYER metal3 ;
         RECT  200.8425 0.0 200.9775 0.135 ;
         LAYER metal4 ;
         RECT  46.4 76.25 46.54 91.34 ;
         LAYER metal3 ;
         RECT  223.7225 0.0 223.8575 0.135 ;
         LAYER metal4 ;
         RECT  2.75 41.475 2.89 63.8775 ;
         LAYER metal3 ;
         RECT  52.1225 0.0 52.2575 0.135 ;
         LAYER metal3 ;
         RECT  349.5625 0.0 349.6975 0.135 ;
         LAYER metal3 ;
         RECT  166.5225 0.0 166.6575 0.135 ;
         LAYER metal3 ;
         RECT  429.6425 0.0 429.7775 0.135 ;
         LAYER metal3 ;
         RECT  120.7625 0.0 120.8975 0.135 ;
         LAYER metal4 ;
         RECT  182.585 51.565 182.725 143.27 ;
         LAYER metal3 ;
         RECT  63.5625 0.0 63.6975 0.135 ;
         LAYER metal3 ;
         RECT  177.9625 0.0 178.0975 0.135 ;
         LAYER metal3 ;
         RECT  235.1625 0.0 235.2975 0.135 ;
         LAYER metal3 ;
         RECT  48.115 59.9375 48.25 60.0725 ;
         LAYER metal3 ;
         RECT  395.3225 0.0 395.4575 0.135 ;
         LAYER metal3 ;
         RECT  189.4025 0.0 189.5375 0.135 ;
         LAYER metal3 ;
         RECT  66.4675 48.865 181.6475 48.935 ;
         LAYER metal3 ;
         RECT  406.7625 0.0 406.8975 0.135 ;
         LAYER metal3 ;
         RECT  66.3325 37.2575 66.4675 37.3925 ;
         LAYER metal3 ;
         RECT  498.2825 0.0 498.4175 0.135 ;
         LAYER metal3 ;
         RECT  326.6825 0.0 326.8175 0.135 ;
         LAYER metal3 ;
         RECT  280.9225 0.0 281.0575 0.135 ;
         LAYER metal3 ;
         RECT  463.9625 0.0 464.0975 0.135 ;
         LAYER metal3 ;
         RECT  383.8825 0.0 384.0175 0.135 ;
         LAYER metal3 ;
         RECT  48.115 54.4775 48.25 54.6125 ;
         LAYER metal4 ;
         RECT  66.86 51.565 67.0 143.27 ;
         LAYER metal4 ;
         RECT  53.26 54.4425 53.4 142.045 ;
         LAYER metal3 ;
         RECT  48.115 70.8575 48.25 70.9925 ;
         LAYER metal3 ;
         RECT  97.8825 0.0 98.0175 0.135 ;
         LAYER metal3 ;
         RECT  48.115 76.3175 48.25 76.4525 ;
         LAYER metal3 ;
         RECT  258.0425 0.0 258.1775 0.135 ;
         LAYER metal3 ;
         RECT  109.3225 0.0 109.4575 0.135 ;
         LAYER metal3 ;
         RECT  246.6025 0.0 246.7375 0.135 ;
         LAYER metal3 ;
         RECT  303.8025 0.0 303.9375 0.135 ;
         LAYER metal4 ;
         RECT  6.385 31.595 6.525 51.495 ;
         LAYER metal3 ;
         RECT  475.4025 0.0 475.5375 0.135 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 529.67 143.3275 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 529.67 143.3275 ;
   LAYER  metal3 ;
      RECT  72.285 0.14 72.7 0.965 ;
      RECT  72.7 0.965 75.145 1.38 ;
      RECT  75.56 0.965 78.005 1.38 ;
      RECT  78.42 0.965 80.865 1.38 ;
      RECT  81.28 0.965 83.725 1.38 ;
      RECT  84.14 0.965 86.585 1.38 ;
      RECT  87.0 0.965 89.445 1.38 ;
      RECT  89.86 0.965 92.305 1.38 ;
      RECT  92.72 0.965 95.165 1.38 ;
      RECT  95.58 0.965 98.025 1.38 ;
      RECT  98.44 0.965 100.885 1.38 ;
      RECT  101.3 0.965 103.745 1.38 ;
      RECT  104.16 0.965 106.605 1.38 ;
      RECT  107.02 0.965 109.465 1.38 ;
      RECT  109.88 0.965 112.325 1.38 ;
      RECT  112.74 0.965 115.185 1.38 ;
      RECT  115.6 0.965 118.045 1.38 ;
      RECT  118.46 0.965 120.905 1.38 ;
      RECT  121.32 0.965 123.765 1.38 ;
      RECT  124.18 0.965 126.625 1.38 ;
      RECT  127.04 0.965 129.485 1.38 ;
      RECT  129.9 0.965 132.345 1.38 ;
      RECT  132.76 0.965 135.205 1.38 ;
      RECT  135.62 0.965 138.065 1.38 ;
      RECT  138.48 0.965 140.925 1.38 ;
      RECT  141.34 0.965 143.785 1.38 ;
      RECT  144.2 0.965 146.645 1.38 ;
      RECT  147.06 0.965 149.505 1.38 ;
      RECT  149.92 0.965 152.365 1.38 ;
      RECT  152.78 0.965 155.225 1.38 ;
      RECT  155.64 0.965 158.085 1.38 ;
      RECT  158.5 0.965 160.945 1.38 ;
      RECT  161.36 0.965 163.805 1.38 ;
      RECT  164.22 0.965 166.665 1.38 ;
      RECT  167.08 0.965 169.525 1.38 ;
      RECT  169.94 0.965 172.385 1.38 ;
      RECT  172.8 0.965 175.245 1.38 ;
      RECT  175.66 0.965 178.105 1.38 ;
      RECT  178.52 0.965 180.965 1.38 ;
      RECT  181.38 0.965 183.825 1.38 ;
      RECT  184.24 0.965 186.685 1.38 ;
      RECT  187.1 0.965 189.545 1.38 ;
      RECT  189.96 0.965 192.405 1.38 ;
      RECT  192.82 0.965 195.265 1.38 ;
      RECT  195.68 0.965 198.125 1.38 ;
      RECT  198.54 0.965 200.985 1.38 ;
      RECT  201.4 0.965 203.845 1.38 ;
      RECT  204.26 0.965 206.705 1.38 ;
      RECT  207.12 0.965 209.565 1.38 ;
      RECT  209.98 0.965 212.425 1.38 ;
      RECT  212.84 0.965 215.285 1.38 ;
      RECT  215.7 0.965 218.145 1.38 ;
      RECT  218.56 0.965 221.005 1.38 ;
      RECT  221.42 0.965 223.865 1.38 ;
      RECT  224.28 0.965 226.725 1.38 ;
      RECT  227.14 0.965 229.585 1.38 ;
      RECT  230.0 0.965 232.445 1.38 ;
      RECT  232.86 0.965 235.305 1.38 ;
      RECT  235.72 0.965 238.165 1.38 ;
      RECT  238.58 0.965 241.025 1.38 ;
      RECT  241.44 0.965 243.885 1.38 ;
      RECT  244.3 0.965 246.745 1.38 ;
      RECT  247.16 0.965 249.605 1.38 ;
      RECT  250.02 0.965 252.465 1.38 ;
      RECT  252.88 0.965 255.325 1.38 ;
      RECT  255.74 0.965 258.185 1.38 ;
      RECT  258.6 0.965 261.045 1.38 ;
      RECT  261.46 0.965 263.905 1.38 ;
      RECT  264.32 0.965 266.765 1.38 ;
      RECT  267.18 0.965 269.625 1.38 ;
      RECT  270.04 0.965 272.485 1.38 ;
      RECT  272.9 0.965 275.345 1.38 ;
      RECT  275.76 0.965 278.205 1.38 ;
      RECT  278.62 0.965 281.065 1.38 ;
      RECT  281.48 0.965 283.925 1.38 ;
      RECT  284.34 0.965 286.785 1.38 ;
      RECT  287.2 0.965 289.645 1.38 ;
      RECT  290.06 0.965 292.505 1.38 ;
      RECT  292.92 0.965 295.365 1.38 ;
      RECT  295.78 0.965 298.225 1.38 ;
      RECT  298.64 0.965 301.085 1.38 ;
      RECT  301.5 0.965 303.945 1.38 ;
      RECT  304.36 0.965 306.805 1.38 ;
      RECT  307.22 0.965 309.665 1.38 ;
      RECT  310.08 0.965 312.525 1.38 ;
      RECT  312.94 0.965 315.385 1.38 ;
      RECT  315.8 0.965 318.245 1.38 ;
      RECT  318.66 0.965 321.105 1.38 ;
      RECT  321.52 0.965 323.965 1.38 ;
      RECT  324.38 0.965 326.825 1.38 ;
      RECT  327.24 0.965 329.685 1.38 ;
      RECT  330.1 0.965 332.545 1.38 ;
      RECT  332.96 0.965 335.405 1.38 ;
      RECT  335.82 0.965 338.265 1.38 ;
      RECT  338.68 0.965 341.125 1.38 ;
      RECT  341.54 0.965 343.985 1.38 ;
      RECT  344.4 0.965 346.845 1.38 ;
      RECT  347.26 0.965 349.705 1.38 ;
      RECT  350.12 0.965 352.565 1.38 ;
      RECT  352.98 0.965 355.425 1.38 ;
      RECT  355.84 0.965 358.285 1.38 ;
      RECT  358.7 0.965 361.145 1.38 ;
      RECT  361.56 0.965 364.005 1.38 ;
      RECT  364.42 0.965 366.865 1.38 ;
      RECT  367.28 0.965 369.725 1.38 ;
      RECT  370.14 0.965 372.585 1.38 ;
      RECT  373.0 0.965 375.445 1.38 ;
      RECT  375.86 0.965 378.305 1.38 ;
      RECT  378.72 0.965 381.165 1.38 ;
      RECT  381.58 0.965 384.025 1.38 ;
      RECT  384.44 0.965 386.885 1.38 ;
      RECT  387.3 0.965 389.745 1.38 ;
      RECT  390.16 0.965 392.605 1.38 ;
      RECT  393.02 0.965 395.465 1.38 ;
      RECT  395.88 0.965 398.325 1.38 ;
      RECT  398.74 0.965 401.185 1.38 ;
      RECT  401.6 0.965 404.045 1.38 ;
      RECT  404.46 0.965 406.905 1.38 ;
      RECT  407.32 0.965 409.765 1.38 ;
      RECT  410.18 0.965 412.625 1.38 ;
      RECT  413.04 0.965 415.485 1.38 ;
      RECT  415.9 0.965 418.345 1.38 ;
      RECT  418.76 0.965 421.205 1.38 ;
      RECT  421.62 0.965 424.065 1.38 ;
      RECT  424.48 0.965 426.925 1.38 ;
      RECT  427.34 0.965 429.785 1.38 ;
      RECT  430.2 0.965 432.645 1.38 ;
      RECT  433.06 0.965 435.505 1.38 ;
      RECT  435.92 0.965 438.365 1.38 ;
      RECT  438.78 0.965 441.225 1.38 ;
      RECT  441.64 0.965 444.085 1.38 ;
      RECT  444.5 0.965 446.945 1.38 ;
      RECT  447.36 0.965 449.805 1.38 ;
      RECT  450.22 0.965 452.665 1.38 ;
      RECT  453.08 0.965 455.525 1.38 ;
      RECT  455.94 0.965 458.385 1.38 ;
      RECT  458.8 0.965 461.245 1.38 ;
      RECT  461.66 0.965 464.105 1.38 ;
      RECT  464.52 0.965 466.965 1.38 ;
      RECT  467.38 0.965 469.825 1.38 ;
      RECT  470.24 0.965 472.685 1.38 ;
      RECT  473.1 0.965 475.545 1.38 ;
      RECT  475.96 0.965 478.405 1.38 ;
      RECT  478.82 0.965 481.265 1.38 ;
      RECT  481.68 0.965 484.125 1.38 ;
      RECT  484.54 0.965 486.985 1.38 ;
      RECT  487.4 0.965 489.845 1.38 ;
      RECT  490.26 0.965 492.705 1.38 ;
      RECT  493.12 0.965 495.565 1.38 ;
      RECT  495.98 0.965 498.425 1.38 ;
      RECT  498.84 0.965 501.285 1.38 ;
      RECT  501.7 0.965 504.145 1.38 ;
      RECT  504.56 0.965 507.005 1.38 ;
      RECT  507.42 0.965 509.865 1.38 ;
      RECT  510.28 0.965 512.725 1.38 ;
      RECT  513.14 0.965 515.585 1.38 ;
      RECT  516.0 0.965 518.445 1.38 ;
      RECT  518.86 0.965 521.305 1.38 ;
      RECT  521.72 0.965 524.165 1.38 ;
      RECT  524.58 0.965 527.025 1.38 ;
      RECT  527.44 0.965 529.67 1.38 ;
      RECT  0.14 77.2825 43.685 77.6975 ;
      RECT  0.14 77.6975 43.685 143.3275 ;
      RECT  43.685 1.38 44.1 77.2825 ;
      RECT  44.1 77.2825 72.285 77.6975 ;
      RECT  44.1 77.6975 72.285 143.3275 ;
      RECT  43.685 77.6975 44.1 80.0125 ;
      RECT  43.685 80.4275 44.1 82.2225 ;
      RECT  43.685 82.6375 44.1 84.9525 ;
      RECT  43.685 85.3675 44.1 87.1625 ;
      RECT  43.685 87.5775 44.1 89.8925 ;
      RECT  43.685 90.3075 44.1 143.3275 ;
      RECT  0.14 1.38 0.145 32.5625 ;
      RECT  0.14 32.5625 0.145 32.9775 ;
      RECT  0.14 32.9775 0.145 77.2825 ;
      RECT  0.145 1.38 0.56 32.5625 ;
      RECT  0.56 1.38 43.685 32.5625 ;
      RECT  0.145 32.9775 0.56 35.2925 ;
      RECT  0.145 35.7075 0.56 77.2825 ;
      RECT  0.56 32.5625 6.3875 32.6475 ;
      RECT  0.56 32.6475 6.3875 32.9775 ;
      RECT  6.3875 32.5625 6.8025 32.6475 ;
      RECT  6.8025 32.5625 43.685 32.6475 ;
      RECT  6.8025 32.6475 43.685 32.9775 ;
      RECT  0.56 32.9775 6.3875 33.0625 ;
      RECT  0.56 33.0625 6.3875 77.2825 ;
      RECT  6.3875 33.0625 6.8025 77.2825 ;
      RECT  6.8025 32.9775 43.685 33.0625 ;
      RECT  6.8025 33.0625 43.685 77.2825 ;
      RECT  0.14 0.965 49.405 1.38 ;
      RECT  49.82 0.965 52.265 1.38 ;
      RECT  52.68 0.965 55.125 1.38 ;
      RECT  55.54 0.965 57.985 1.38 ;
      RECT  58.4 0.965 60.845 1.38 ;
      RECT  61.26 0.965 63.705 1.38 ;
      RECT  64.12 0.965 66.565 1.38 ;
      RECT  66.98 0.965 69.425 1.38 ;
      RECT  69.84 0.965 72.285 1.38 ;
      RECT  44.1 44.2125 68.5725 44.6275 ;
      RECT  68.9875 44.2125 69.2775 44.6275 ;
      RECT  69.6925 44.2125 69.9825 44.6275 ;
      RECT  70.3975 44.2125 70.6875 44.6275 ;
      RECT  71.1025 44.2125 71.3925 44.6275 ;
      RECT  72.5125 44.2125 72.7 44.6275 ;
      RECT  71.8075 44.2125 72.0975 44.6275 ;
      RECT  72.7 44.2125 72.8025 44.6275 ;
      RECT  73.2175 44.2125 73.5075 44.6275 ;
      RECT  73.9225 44.2125 74.2125 44.6275 ;
      RECT  74.6275 44.2125 74.9175 44.6275 ;
      RECT  75.3325 44.2125 75.6225 44.6275 ;
      RECT  76.0375 44.2125 76.3275 44.6275 ;
      RECT  76.7425 44.2125 77.0325 44.6275 ;
      RECT  77.4475 44.2125 77.7375 44.6275 ;
      RECT  78.1525 44.2125 78.4425 44.6275 ;
      RECT  78.8575 44.2125 79.1475 44.6275 ;
      RECT  79.5625 44.2125 79.8525 44.6275 ;
      RECT  80.2675 44.2125 80.5575 44.6275 ;
      RECT  80.9725 44.2125 81.2625 44.6275 ;
      RECT  81.6775 44.2125 81.9675 44.6275 ;
      RECT  82.3825 44.2125 82.6725 44.6275 ;
      RECT  83.0875 44.2125 83.3775 44.6275 ;
      RECT  83.7925 44.2125 84.0825 44.6275 ;
      RECT  84.4975 44.2125 84.7875 44.6275 ;
      RECT  85.2025 44.2125 85.4925 44.6275 ;
      RECT  85.9075 44.2125 86.1975 44.6275 ;
      RECT  86.6125 44.2125 86.9025 44.6275 ;
      RECT  87.3175 44.2125 87.6075 44.6275 ;
      RECT  88.0225 44.2125 88.3125 44.6275 ;
      RECT  88.7275 44.2125 89.0175 44.6275 ;
      RECT  89.4325 44.2125 89.7225 44.6275 ;
      RECT  90.1375 44.2125 90.4275 44.6275 ;
      RECT  90.8425 44.2125 91.1325 44.6275 ;
      RECT  91.5475 44.2125 91.8375 44.6275 ;
      RECT  92.2525 44.2125 92.5425 44.6275 ;
      RECT  92.9575 44.2125 93.2475 44.6275 ;
      RECT  93.6625 44.2125 93.9525 44.6275 ;
      RECT  94.3675 44.2125 94.6575 44.6275 ;
      RECT  95.0725 44.2125 95.3625 44.6275 ;
      RECT  95.7775 44.2125 96.0675 44.6275 ;
      RECT  96.4825 44.2125 96.7725 44.6275 ;
      RECT  97.1875 44.2125 97.4775 44.6275 ;
      RECT  97.8925 44.2125 98.1825 44.6275 ;
      RECT  98.5975 44.2125 98.8875 44.6275 ;
      RECT  99.3025 44.2125 99.5925 44.6275 ;
      RECT  100.0075 44.2125 100.2975 44.6275 ;
      RECT  100.7125 44.2125 101.0025 44.6275 ;
      RECT  101.4175 44.2125 101.7075 44.6275 ;
      RECT  102.1225 44.2125 102.4125 44.6275 ;
      RECT  102.8275 44.2125 103.1175 44.6275 ;
      RECT  103.5325 44.2125 103.8225 44.6275 ;
      RECT  104.2375 44.2125 104.5275 44.6275 ;
      RECT  104.9425 44.2125 105.2325 44.6275 ;
      RECT  105.6475 44.2125 105.9375 44.6275 ;
      RECT  106.3525 44.2125 106.6425 44.6275 ;
      RECT  107.0575 44.2125 107.3475 44.6275 ;
      RECT  107.7625 44.2125 108.0525 44.6275 ;
      RECT  108.4675 44.2125 108.7575 44.6275 ;
      RECT  109.1725 44.2125 109.4625 44.6275 ;
      RECT  109.8775 44.2125 110.1675 44.6275 ;
      RECT  110.5825 44.2125 110.8725 44.6275 ;
      RECT  111.2875 44.2125 111.5775 44.6275 ;
      RECT  111.9925 44.2125 112.2825 44.6275 ;
      RECT  112.6975 44.2125 112.9875 44.6275 ;
      RECT  113.4025 44.2125 113.6925 44.6275 ;
      RECT  114.1075 44.2125 114.3975 44.6275 ;
      RECT  114.8125 44.2125 115.1025 44.6275 ;
      RECT  115.5175 44.2125 115.8075 44.6275 ;
      RECT  116.2225 44.2125 116.5125 44.6275 ;
      RECT  116.9275 44.2125 117.2175 44.6275 ;
      RECT  117.6325 44.2125 117.9225 44.6275 ;
      RECT  118.3375 44.2125 118.6275 44.6275 ;
      RECT  119.0425 44.2125 119.3325 44.6275 ;
      RECT  119.7475 44.2125 120.0375 44.6275 ;
      RECT  120.4525 44.2125 120.7425 44.6275 ;
      RECT  121.1575 44.2125 121.4475 44.6275 ;
      RECT  121.8625 44.2125 122.1525 44.6275 ;
      RECT  122.5675 44.2125 122.8575 44.6275 ;
      RECT  123.2725 44.2125 123.5625 44.6275 ;
      RECT  123.9775 44.2125 124.2675 44.6275 ;
      RECT  124.6825 44.2125 124.9725 44.6275 ;
      RECT  125.3875 44.2125 125.6775 44.6275 ;
      RECT  126.0925 44.2125 126.3825 44.6275 ;
      RECT  126.7975 44.2125 127.0875 44.6275 ;
      RECT  127.5025 44.2125 127.7925 44.6275 ;
      RECT  128.2075 44.2125 128.4975 44.6275 ;
      RECT  128.9125 44.2125 129.2025 44.6275 ;
      RECT  129.6175 44.2125 129.9075 44.6275 ;
      RECT  130.3225 44.2125 130.6125 44.6275 ;
      RECT  131.0275 44.2125 131.3175 44.6275 ;
      RECT  131.7325 44.2125 132.0225 44.6275 ;
      RECT  132.4375 44.2125 132.7275 44.6275 ;
      RECT  133.1425 44.2125 133.4325 44.6275 ;
      RECT  133.8475 44.2125 134.1375 44.6275 ;
      RECT  134.5525 44.2125 134.8425 44.6275 ;
      RECT  135.2575 44.2125 135.5475 44.6275 ;
      RECT  135.9625 44.2125 136.2525 44.6275 ;
      RECT  136.6675 44.2125 136.9575 44.6275 ;
      RECT  137.3725 44.2125 137.6625 44.6275 ;
      RECT  138.0775 44.2125 138.3675 44.6275 ;
      RECT  138.7825 44.2125 139.0725 44.6275 ;
      RECT  139.4875 44.2125 139.7775 44.6275 ;
      RECT  140.1925 44.2125 140.4825 44.6275 ;
      RECT  140.8975 44.2125 141.1875 44.6275 ;
      RECT  141.6025 44.2125 141.8925 44.6275 ;
      RECT  142.3075 44.2125 142.5975 44.6275 ;
      RECT  143.0125 44.2125 143.3025 44.6275 ;
      RECT  143.7175 44.2125 144.0075 44.6275 ;
      RECT  144.4225 44.2125 144.7125 44.6275 ;
      RECT  145.1275 44.2125 145.4175 44.6275 ;
      RECT  145.8325 44.2125 146.1225 44.6275 ;
      RECT  146.5375 44.2125 146.8275 44.6275 ;
      RECT  147.2425 44.2125 147.5325 44.6275 ;
      RECT  147.9475 44.2125 148.2375 44.6275 ;
      RECT  148.6525 44.2125 148.9425 44.6275 ;
      RECT  149.3575 44.2125 149.6475 44.6275 ;
      RECT  150.0625 44.2125 150.3525 44.6275 ;
      RECT  150.7675 44.2125 151.0575 44.6275 ;
      RECT  151.4725 44.2125 151.7625 44.6275 ;
      RECT  152.1775 44.2125 152.4675 44.6275 ;
      RECT  152.8825 44.2125 153.1725 44.6275 ;
      RECT  153.5875 44.2125 153.8775 44.6275 ;
      RECT  154.2925 44.2125 154.5825 44.6275 ;
      RECT  154.9975 44.2125 155.2875 44.6275 ;
      RECT  155.7025 44.2125 155.9925 44.6275 ;
      RECT  156.4075 44.2125 156.6975 44.6275 ;
      RECT  157.1125 44.2125 157.4025 44.6275 ;
      RECT  157.8175 44.2125 158.1075 44.6275 ;
      RECT  158.5225 44.2125 158.8125 44.6275 ;
      RECT  159.2275 44.2125 159.5175 44.6275 ;
      RECT  159.9325 44.2125 160.2225 44.6275 ;
      RECT  160.6375 44.2125 160.9275 44.6275 ;
      RECT  161.3425 44.2125 161.6325 44.6275 ;
      RECT  162.0475 44.2125 162.3375 44.6275 ;
      RECT  162.7525 44.2125 163.0425 44.6275 ;
      RECT  163.4575 44.2125 163.7475 44.6275 ;
      RECT  164.1625 44.2125 164.4525 44.6275 ;
      RECT  164.8675 44.2125 165.1575 44.6275 ;
      RECT  165.5725 44.2125 165.8625 44.6275 ;
      RECT  166.2775 44.2125 166.5675 44.6275 ;
      RECT  166.9825 44.2125 167.2725 44.6275 ;
      RECT  167.6875 44.2125 167.9775 44.6275 ;
      RECT  168.3925 44.2125 168.6825 44.6275 ;
      RECT  169.0975 44.2125 169.3875 44.6275 ;
      RECT  169.8025 44.2125 170.0925 44.6275 ;
      RECT  170.5075 44.2125 170.7975 44.6275 ;
      RECT  171.2125 44.2125 171.5025 44.6275 ;
      RECT  171.9175 44.2125 172.2075 44.6275 ;
      RECT  172.6225 44.2125 172.9125 44.6275 ;
      RECT  173.3275 44.2125 173.6175 44.6275 ;
      RECT  174.0325 44.2125 174.3225 44.6275 ;
      RECT  174.7375 44.2125 175.0275 44.6275 ;
      RECT  175.4425 44.2125 175.7325 44.6275 ;
      RECT  176.1475 44.2125 176.4375 44.6275 ;
      RECT  176.8525 44.2125 177.1425 44.6275 ;
      RECT  177.5575 44.2125 177.8475 44.6275 ;
      RECT  178.2625 44.2125 178.5525 44.6275 ;
      RECT  178.9675 44.2125 179.2575 44.6275 ;
      RECT  179.6725 44.2125 179.9625 44.6275 ;
      RECT  180.3775 44.2125 180.6675 44.6275 ;
      RECT  181.0825 44.2125 529.67 44.6275 ;
      RECT  44.1 1.38 49.1225 2.33 ;
      RECT  44.1 2.33 49.1225 2.745 ;
      RECT  44.1 2.745 49.1225 44.2125 ;
      RECT  49.1225 1.38 49.5375 2.33 ;
      RECT  49.1225 2.745 49.5375 44.2125 ;
      RECT  49.5375 1.38 68.5725 2.33 ;
      RECT  68.5725 1.38 68.9875 39.905 ;
      RECT  72.5125 1.38 72.7 39.905 ;
      RECT  72.7 1.38 72.8025 39.905 ;
      RECT  72.8025 1.38 73.2175 39.905 ;
      RECT  181.7525 39.905 529.67 40.255 ;
      RECT  181.7525 40.255 529.67 44.2125 ;
      RECT  49.5375 39.905 66.3275 40.255 ;
      RECT  49.5375 40.255 66.3275 44.2125 ;
      RECT  73.2175 1.38 94.8825 2.33 ;
      RECT  73.2175 2.745 94.8825 39.905 ;
      RECT  94.8825 1.38 95.2975 2.33 ;
      RECT  94.8825 2.745 95.2975 39.905 ;
      RECT  95.2975 1.38 181.7525 2.33 ;
      RECT  181.7525 1.38 380.8825 2.33 ;
      RECT  181.7525 2.745 380.8825 39.905 ;
      RECT  380.8825 1.38 381.2975 2.33 ;
      RECT  380.8825 2.745 381.2975 39.905 ;
      RECT  381.2975 1.38 529.67 2.33 ;
      RECT  381.2975 2.745 529.67 39.905 ;
      RECT  518.5775 2.33 529.67 2.745 ;
      RECT  175.3775 2.33 181.7525 2.745 ;
      RECT  49.5375 2.745 66.1925 38.9375 ;
      RECT  49.5375 38.9375 66.1925 39.3525 ;
      RECT  49.5375 39.3525 66.1925 39.905 ;
      RECT  66.1925 39.3525 66.3275 39.905 ;
      RECT  66.3275 39.3525 66.6075 39.905 ;
      RECT  66.6075 2.745 68.5725 38.9375 ;
      RECT  66.6075 38.9375 68.5725 39.3525 ;
      RECT  66.6075 39.3525 68.5725 39.905 ;
      RECT  495.6975 2.33 506.7225 2.745 ;
      RECT  507.1375 2.33 518.1625 2.745 ;
      RECT  301.2175 2.33 312.2425 2.745 ;
      RECT  181.7525 2.33 186.4025 2.745 ;
      RECT  186.8175 2.33 197.8425 2.745 ;
      RECT  44.1 44.6275 65.1825 52.9725 ;
      RECT  44.1 52.9725 65.1825 53.3875 ;
      RECT  65.1825 44.6275 65.5975 52.9725 ;
      RECT  65.1825 53.3875 65.5975 77.2825 ;
      RECT  65.5975 52.9725 68.5725 53.3875 ;
      RECT  65.5975 53.3875 68.5725 77.2825 ;
      RECT  95.2975 2.745 181.3375 38.9375 ;
      RECT  95.2975 38.9375 181.3375 39.3525 ;
      RECT  95.2975 39.3525 181.3375 39.905 ;
      RECT  181.3375 39.3525 181.7525 39.905 ;
      RECT  266.8975 2.33 277.9225 2.745 ;
      RECT  198.2575 2.33 209.2825 2.745 ;
      RECT  209.6975 2.33 220.7225 2.745 ;
      RECT  472.8175 2.33 483.8425 2.745 ;
      RECT  484.2575 2.33 495.2825 2.745 ;
      RECT  44.1 63.8925 49.5025 64.3075 ;
      RECT  49.9175 63.8925 65.1825 64.3075 ;
      RECT  49.9175 64.3075 65.1825 77.2825 ;
      RECT  68.5725 51.08 68.9875 77.2825 ;
      RECT  68.9875 51.08 72.285 77.2825 ;
      RECT  72.285 51.08 72.5125 143.3275 ;
      RECT  72.5125 51.08 72.7 143.3275 ;
      RECT  72.7 51.08 72.8025 143.3275 ;
      RECT  72.8025 51.08 73.2175 143.3275 ;
      RECT  73.2175 51.08 181.7525 143.3275 ;
      RECT  181.7525 50.73 529.67 51.08 ;
      RECT  181.7525 51.08 529.67 143.3275 ;
      RECT  65.5975 44.6275 66.3275 50.73 ;
      RECT  65.5975 50.73 66.3275 51.08 ;
      RECT  65.5975 51.08 66.3275 52.9725 ;
      RECT  66.3275 51.08 68.5725 52.9725 ;
      RECT  49.9175 53.3875 55.675 53.63 ;
      RECT  49.9175 53.63 55.675 54.045 ;
      RECT  49.9175 54.045 55.675 63.8925 ;
      RECT  55.675 53.3875 56.09 53.63 ;
      RECT  55.675 54.045 56.09 63.8925 ;
      RECT  56.09 53.3875 65.1825 53.63 ;
      RECT  56.09 53.63 65.1825 54.045 ;
      RECT  56.09 54.045 65.1825 63.8925 ;
      RECT  312.6575 2.33 323.6825 2.745 ;
      RECT  381.2975 2.33 392.3225 2.745 ;
      RECT  392.7375 2.33 403.7625 2.745 ;
      RECT  427.0575 2.33 438.0825 2.745 ;
      RECT  118.1775 2.33 129.2025 2.745 ;
      RECT  129.6175 2.33 140.6425 2.745 ;
      RECT  221.1375 2.33 232.1625 2.745 ;
      RECT  232.5775 2.33 243.6025 2.745 ;
      RECT  369.8575 2.33 380.8825 2.745 ;
      RECT  346.9775 2.33 358.0025 2.745 ;
      RECT  358.4175 2.33 369.4425 2.745 ;
      RECT  49.5025 72.4975 49.9175 74.8125 ;
      RECT  49.5025 75.2275 49.9175 77.2825 ;
      RECT  163.9375 2.33 174.9625 2.745 ;
      RECT  244.0175 2.33 255.0425 2.745 ;
      RECT  255.4575 2.33 266.4825 2.745 ;
      RECT  278.3375 2.33 289.3625 2.745 ;
      RECT  289.7775 2.33 300.8025 2.745 ;
      RECT  68.9875 1.38 72.0025 2.33 ;
      RECT  68.9875 2.33 72.0025 2.745 ;
      RECT  68.9875 2.745 72.0025 39.905 ;
      RECT  72.0025 1.38 72.285 2.33 ;
      RECT  72.0025 2.745 72.285 39.905 ;
      RECT  72.285 1.38 72.4175 2.33 ;
      RECT  72.285 2.745 72.4175 39.905 ;
      RECT  72.4175 1.38 72.5125 2.33 ;
      RECT  72.4175 2.33 72.5125 2.745 ;
      RECT  72.4175 2.745 72.5125 39.905 ;
      RECT  49.5025 58.8475 49.9175 63.8925 ;
      RECT  404.1775 2.33 415.2025 2.745 ;
      RECT  415.6175 2.33 426.6425 2.745 ;
      RECT  73.2175 2.33 83.4425 2.745 ;
      RECT  83.8575 2.33 94.8825 2.745 ;
      RECT  49.5025 64.3075 49.9175 66.6225 ;
      RECT  49.5025 67.0375 49.9175 72.0825 ;
      RECT  324.0975 2.33 335.1225 2.745 ;
      RECT  335.5375 2.33 346.5625 2.745 ;
      RECT  461.3775 2.33 472.4025 2.745 ;
      RECT  49.5025 53.3875 49.9175 55.7025 ;
      RECT  49.5025 56.1175 49.9175 58.4325 ;
      RECT  68.5725 44.6275 68.9875 46.8325 ;
      RECT  68.9875 44.6275 72.285 46.8325 ;
      RECT  72.285 44.6275 72.5125 46.8325 ;
      RECT  72.5125 44.6275 72.7 46.8325 ;
      RECT  72.7 44.6275 72.8025 46.8325 ;
      RECT  72.8025 44.6275 73.2175 46.8325 ;
      RECT  73.2175 44.6275 181.7525 46.8325 ;
      RECT  66.3275 44.6275 68.5725 46.8325 ;
      RECT  49.5375 2.33 60.5625 2.745 ;
      RECT  60.9775 2.33 68.5725 2.745 ;
      RECT  438.4975 2.33 449.5225 2.745 ;
      RECT  449.9375 2.33 460.9625 2.745 ;
      RECT  95.2975 2.33 106.3225 2.745 ;
      RECT  106.7375 2.33 117.7625 2.745 ;
      RECT  141.0575 2.33 152.0825 2.745 ;
      RECT  152.4975 2.33 163.5225 2.745 ;
      RECT  181.3375 2.745 181.7525 37.1175 ;
      RECT  181.3375 37.5325 181.7525 38.9375 ;
      RECT  72.7 0.275 452.3825 0.965 ;
      RECT  452.3825 0.275 452.7975 0.965 ;
      RECT  452.7975 0.275 529.67 0.965 ;
      RECT  68.5725 40.255 68.9875 41.955 ;
      RECT  68.5725 42.305 68.9875 44.2125 ;
      RECT  68.9875 40.255 72.285 41.955 ;
      RECT  68.9875 42.305 72.285 44.2125 ;
      RECT  72.285 40.255 72.5125 41.955 ;
      RECT  72.285 42.305 72.5125 44.2125 ;
      RECT  72.5125 40.255 72.7 41.955 ;
      RECT  72.5125 42.305 72.7 44.2125 ;
      RECT  72.7 40.255 72.8025 41.955 ;
      RECT  72.7 42.305 72.8025 44.2125 ;
      RECT  72.8025 40.255 73.2175 41.955 ;
      RECT  72.8025 42.305 73.2175 44.2125 ;
      RECT  73.2175 40.255 181.7525 41.955 ;
      RECT  73.2175 42.305 181.7525 44.2125 ;
      RECT  66.3275 40.255 68.5725 41.955 ;
      RECT  66.3275 42.305 68.5725 44.2125 ;
      RECT  441.3575 0.14 452.3825 0.275 ;
      RECT  44.1 64.3075 47.975 67.9875 ;
      RECT  44.1 67.9875 47.975 68.4025 ;
      RECT  44.1 68.4025 47.975 77.2825 ;
      RECT  48.39 64.3075 49.5025 67.9875 ;
      RECT  48.39 67.9875 49.5025 68.4025 ;
      RECT  48.39 68.4025 49.5025 77.2825 ;
      RECT  521.4375 0.14 529.67 0.275 ;
      RECT  44.1 53.3875 47.975 62.5275 ;
      RECT  44.1 62.5275 47.975 62.9425 ;
      RECT  44.1 62.9425 47.975 63.8925 ;
      RECT  47.975 62.9425 48.39 63.8925 ;
      RECT  48.39 53.3875 49.5025 62.5275 ;
      RECT  48.39 62.5275 49.5025 62.9425 ;
      RECT  48.39 62.9425 49.5025 63.8925 ;
      RECT  143.9175 0.14 154.9425 0.275 ;
      RECT  47.975 64.3075 48.39 65.2575 ;
      RECT  47.975 65.6725 48.39 67.9875 ;
      RECT  132.4775 0.14 143.5025 0.275 ;
      RECT  509.9975 0.14 521.0225 0.275 ;
      RECT  72.7 0.14 74.8625 0.275 ;
      RECT  75.2775 0.14 86.3025 0.275 ;
      RECT  361.2775 0.14 372.3025 0.275 ;
      RECT  201.1175 0.14 212.1425 0.275 ;
      RECT  212.5575 0.14 223.5825 0.275 ;
      RECT  0.14 0.14 51.9825 0.275 ;
      RECT  0.14 0.275 51.9825 0.965 ;
      RECT  51.9825 0.275 52.3975 0.965 ;
      RECT  52.3975 0.275 72.285 0.965 ;
      RECT  338.3975 0.14 349.4225 0.275 ;
      RECT  349.8375 0.14 360.8625 0.275 ;
      RECT  155.3575 0.14 166.3825 0.275 ;
      RECT  418.4775 0.14 429.5025 0.275 ;
      RECT  429.9175 0.14 440.9425 0.275 ;
      RECT  121.0375 0.14 132.0625 0.275 ;
      RECT  52.3975 0.14 63.4225 0.275 ;
      RECT  63.8375 0.14 72.285 0.275 ;
      RECT  166.7975 0.14 177.8225 0.275 ;
      RECT  223.9975 0.14 235.0225 0.275 ;
      RECT  47.975 57.4825 48.39 59.7975 ;
      RECT  47.975 60.2125 48.39 62.5275 ;
      RECT  178.2375 0.14 189.2625 0.275 ;
      RECT  189.6775 0.14 200.7025 0.275 ;
      RECT  181.7525 44.6275 181.7875 48.725 ;
      RECT  181.7525 49.075 181.7875 50.73 ;
      RECT  181.7875 44.6275 529.67 48.725 ;
      RECT  181.7875 48.725 529.67 49.075 ;
      RECT  181.7875 49.075 529.67 50.73 ;
      RECT  68.5725 47.1825 68.9875 48.725 ;
      RECT  68.5725 49.075 68.9875 50.73 ;
      RECT  68.9875 47.1825 72.285 48.725 ;
      RECT  68.9875 49.075 72.285 50.73 ;
      RECT  72.285 47.1825 72.5125 48.725 ;
      RECT  72.285 49.075 72.5125 50.73 ;
      RECT  72.5125 47.1825 72.7 48.725 ;
      RECT  72.5125 49.075 72.7 50.73 ;
      RECT  72.7 47.1825 72.8025 48.725 ;
      RECT  72.7 49.075 72.8025 50.73 ;
      RECT  72.8025 47.1825 73.2175 48.725 ;
      RECT  72.8025 49.075 73.2175 50.73 ;
      RECT  73.2175 47.1825 181.7525 48.725 ;
      RECT  73.2175 49.075 181.7525 50.73 ;
      RECT  66.3275 47.1825 68.5725 48.725 ;
      RECT  66.3275 49.075 68.5725 50.73 ;
      RECT  395.5975 0.14 406.6225 0.275 ;
      RECT  407.0375 0.14 418.0625 0.275 ;
      RECT  66.1925 2.745 66.3275 37.1175 ;
      RECT  66.1925 37.5325 66.3275 38.9375 ;
      RECT  66.3275 2.745 66.6075 37.1175 ;
      RECT  66.3275 37.5325 66.6075 38.9375 ;
      RECT  487.1175 0.14 498.1425 0.275 ;
      RECT  498.5575 0.14 509.5825 0.275 ;
      RECT  315.5175 0.14 326.5425 0.275 ;
      RECT  326.9575 0.14 337.9825 0.275 ;
      RECT  269.7575 0.14 280.7825 0.275 ;
      RECT  281.1975 0.14 292.2225 0.275 ;
      RECT  452.7975 0.14 463.8225 0.275 ;
      RECT  372.7175 0.14 383.7425 0.275 ;
      RECT  384.1575 0.14 395.1825 0.275 ;
      RECT  47.975 53.3875 48.39 54.3375 ;
      RECT  47.975 54.7525 48.39 57.0675 ;
      RECT  47.975 68.4025 48.39 70.7175 ;
      RECT  47.975 71.1325 48.39 73.4475 ;
      RECT  86.7175 0.14 97.7425 0.275 ;
      RECT  47.975 73.8625 48.39 76.1775 ;
      RECT  47.975 76.5925 48.39 77.2825 ;
      RECT  258.3175 0.14 269.3425 0.275 ;
      RECT  98.1575 0.14 109.1825 0.275 ;
      RECT  109.5975 0.14 120.6225 0.275 ;
      RECT  235.4375 0.14 246.4625 0.275 ;
      RECT  246.8775 0.14 257.9025 0.275 ;
      RECT  292.6375 0.14 303.6625 0.275 ;
      RECT  304.0775 0.14 315.1025 0.275 ;
      RECT  464.2375 0.14 475.2625 0.275 ;
      RECT  475.6775 0.14 486.7025 0.275 ;
   LAYER  metal4 ;
      RECT  0.14 142.325 54.915 143.3275 ;
      RECT  54.915 142.325 55.615 143.3275 ;
      RECT  45.98 0.14 46.68 33.785 ;
      RECT  45.98 49.305 46.68 54.195 ;
      RECT  46.68 0.14 54.915 33.785 ;
      RECT  46.68 33.785 54.915 49.305 ;
      RECT  0.14 0.14 0.42 31.315 ;
      RECT  0.14 76.035 43.26 91.555 ;
      RECT  0.14 91.555 43.26 142.325 ;
      RECT  43.26 54.195 43.96 76.035 ;
      RECT  43.26 91.555 43.96 142.325 ;
      RECT  65.04 142.255 65.74 142.325 ;
      RECT  55.615 0.14 182.765 51.285 ;
      RECT  182.765 0.14 183.465 51.285 ;
      RECT  183.465 0.14 529.67 51.285 ;
      RECT  183.465 51.285 529.67 54.195 ;
      RECT  183.465 142.325 529.67 143.3275 ;
      RECT  183.465 54.195 529.67 142.255 ;
      RECT  183.465 142.255 529.67 142.325 ;
      RECT  55.615 142.325 66.12 143.3275 ;
      RECT  65.74 54.195 66.12 142.255 ;
      RECT  65.74 142.255 66.12 142.325 ;
      RECT  0.14 49.305 0.4075 54.195 ;
      RECT  0.14 36.955 0.4075 41.1625 ;
      RECT  0.14 41.1625 0.4075 49.305 ;
      RECT  0.4075 36.955 0.42 41.1625 ;
      RECT  0.42 36.955 1.1075 41.1625 ;
      RECT  0.14 54.195 0.4075 64.125 ;
      RECT  0.14 64.125 0.4075 76.035 ;
      RECT  0.4075 64.125 1.1075 76.035 ;
      RECT  0.42 0.14 4.565 31.25 ;
      RECT  0.42 31.25 4.565 31.315 ;
      RECT  4.565 0.14 5.265 31.25 ;
      RECT  5.265 0.14 45.98 31.25 ;
      RECT  5.265 31.25 45.98 31.315 ;
      RECT  0.42 31.315 4.565 33.785 ;
      RECT  0.42 33.785 4.565 36.955 ;
      RECT  1.1075 36.955 4.565 37.02 ;
      RECT  1.1075 37.02 4.565 41.1625 ;
      RECT  4.565 37.02 5.265 41.1625 ;
      RECT  54.915 0.14 55.475 54.1625 ;
      RECT  54.915 54.1625 55.475 54.195 ;
      RECT  55.475 0.14 55.615 54.1625 ;
      RECT  56.175 54.195 65.04 142.255 ;
      RECT  55.615 142.2875 56.175 142.325 ;
      RECT  56.175 142.255 65.04 142.2875 ;
      RECT  56.175 142.2875 65.04 142.325 ;
      RECT  55.615 51.285 56.175 54.1625 ;
      RECT  56.175 51.285 66.12 54.1625 ;
      RECT  56.175 54.1625 66.12 54.195 ;
      RECT  43.96 54.195 46.12 75.97 ;
      RECT  43.96 75.97 46.12 76.035 ;
      RECT  46.12 54.195 46.82 75.97 ;
      RECT  43.96 76.035 46.12 91.555 ;
      RECT  43.96 91.555 46.12 91.62 ;
      RECT  43.96 91.62 46.12 142.325 ;
      RECT  46.12 91.62 46.82 142.325 ;
      RECT  1.1075 49.305 2.47 54.195 ;
      RECT  1.1075 41.1625 2.47 41.195 ;
      RECT  1.1075 41.195 2.47 49.305 ;
      RECT  2.47 41.1625 3.17 41.195 ;
      RECT  1.1075 54.195 2.47 64.125 ;
      RECT  3.17 54.195 43.26 64.125 ;
      RECT  1.1075 64.125 2.47 64.1575 ;
      RECT  1.1075 64.1575 2.47 76.035 ;
      RECT  2.47 64.1575 3.17 76.035 ;
      RECT  3.17 64.125 43.26 64.1575 ;
      RECT  3.17 64.1575 43.26 76.035 ;
      RECT  67.28 51.285 182.305 54.195 ;
      RECT  67.28 142.325 182.305 143.3275 ;
      RECT  67.28 54.195 182.305 142.255 ;
      RECT  67.28 142.255 182.305 142.325 ;
      RECT  46.68 49.305 52.98 54.1625 ;
      RECT  46.68 54.1625 52.98 54.195 ;
      RECT  52.98 49.305 53.68 54.1625 ;
      RECT  53.68 49.305 54.915 54.1625 ;
      RECT  53.68 54.1625 54.915 54.195 ;
      RECT  46.82 54.195 52.98 75.97 ;
      RECT  53.68 54.195 54.915 75.97 ;
      RECT  46.82 75.97 52.98 76.035 ;
      RECT  53.68 75.97 54.915 76.035 ;
      RECT  46.82 76.035 52.98 91.555 ;
      RECT  53.68 76.035 54.915 91.555 ;
      RECT  46.82 91.555 52.98 91.62 ;
      RECT  53.68 91.555 54.915 91.62 ;
      RECT  46.82 91.62 52.98 142.325 ;
      RECT  53.68 91.62 54.915 142.325 ;
      RECT  5.265 31.315 6.105 33.785 ;
      RECT  6.805 31.315 45.98 33.785 ;
      RECT  5.265 33.785 6.105 36.955 ;
      RECT  6.805 33.785 45.98 36.955 ;
      RECT  5.265 36.955 6.105 37.02 ;
      RECT  6.805 36.955 45.98 37.02 ;
      RECT  5.265 37.02 6.105 41.1625 ;
      RECT  6.805 37.02 45.98 41.1625 ;
      RECT  3.17 49.305 6.105 51.775 ;
      RECT  3.17 51.775 6.105 54.195 ;
      RECT  6.105 51.775 6.805 54.195 ;
      RECT  6.805 49.305 45.98 51.775 ;
      RECT  6.805 51.775 45.98 54.195 ;
      RECT  3.17 41.1625 6.105 41.195 ;
      RECT  6.805 41.1625 45.98 41.195 ;
      RECT  3.17 41.195 6.105 49.305 ;
      RECT  6.805 41.195 45.98 49.305 ;
   END
END    freepdk45_sram_1rw0r_64x160_20
END    LIBRARY
