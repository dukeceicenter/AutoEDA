../macros/freepdk45_sram_1rw0r_45x512/freepdk45_sram_1rw0r_45x512.lef