VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_2048x8_2
   CLASS BLOCK ;
   SIZE 226.63 BY 292.065 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.9725 1.105 42.1075 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.8325 1.105 44.9675 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.6925 1.105 47.8275 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.5525 1.105 50.6875 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.4125 1.105 53.5475 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.2725 1.105 56.4075 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.1325 1.105 59.2675 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.9925 1.105 62.1275 1.24 ;
      END
   END din0[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  19.0925 1.105 19.2275 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.9525 1.105 22.0875 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.8125 1.105 24.9475 1.24 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.6725 1.105 27.8075 1.24 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3725 82.54 13.5075 82.675 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3725 85.27 13.5075 85.405 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3725 87.48 13.5075 87.615 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3725 90.21 13.5075 90.345 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3725 92.42 13.5075 92.555 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3725 95.15 13.5075 95.285 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3725 97.36 13.5075 97.495 ;
      END
   END addr0[10]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.4025 290.825 204.5375 290.96 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.5425 290.825 201.6775 290.96 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.6825 290.825 198.8175 290.96 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.8225 290.825 195.9575 290.96 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.9825 50.43 213.1175 50.565 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.9825 47.7 213.1175 47.835 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.9825 45.49 213.1175 45.625 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.9825 42.76 213.1175 42.895 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.9825 40.55 213.1175 40.685 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.9825 37.82 213.1175 37.955 ;
      END
   END addr1[9]
   PIN addr1[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.9825 35.61 213.1175 35.745 ;
      END
   END addr1[10]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.2875 31.97 0.4225 32.105 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.2075 259.81 226.3425 259.945 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 32.055 6.3825 32.19 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.1075 259.725 220.2425 259.86 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.5325 1.105 30.6675 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.3925 1.105 33.5275 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.2525 1.105 36.3875 1.24 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.1125 1.105 39.2475 1.24 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.915 257.8775 38.05 258.0125 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.715 257.8775 56.85 258.0125 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.515 257.8775 75.65 258.0125 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.315 257.8775 94.45 258.0125 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.115 257.8775 113.25 258.0125 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.915 257.8775 132.05 258.0125 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.715 257.8775 150.85 258.0125 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.515 257.8775 169.65 258.0125 ;
      END
   END dout1[7]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  34.73 37.4575 170.32 37.5275 ;
         LAYER metal3 ;
         RECT  26.8275 50.8275 26.9625 50.9625 ;
         LAYER metal3 ;
         RECT  206.065 64.99 206.2 65.125 ;
         LAYER metal4 ;
         RECT  199.9475 51.5325 200.0875 243.1025 ;
         LAYER metal3 ;
         RECT  20.095 56.02 20.23 56.155 ;
         LAYER metal3 ;
         RECT  34.73 47.6675 188.415 47.7375 ;
         LAYER metal4 ;
         RECT  0.6875 40.71 0.8275 63.1125 ;
         LAYER metal3 ;
         RECT  20.095 62.0 20.23 62.135 ;
         LAYER metal4 ;
         RECT  13.0875 81.4325 13.2275 98.9275 ;
         LAYER metal3 ;
         RECT  19.75 73.96 19.885 74.095 ;
         LAYER metal3 ;
         RECT  30.25 2.47 30.385 2.605 ;
         LAYER metal3 ;
         RECT  206.41 70.97 206.545 71.105 ;
         LAYER metal4 ;
         RECT  34.6625 48.3625 34.8025 245.9525 ;
         LAYER metal4 ;
         RECT  192.5725 51.5325 192.7125 243.0325 ;
         LAYER metal3 ;
         RECT  206.41 79.94 206.545 80.075 ;
         LAYER metal3 ;
         RECT  206.41 76.95 206.545 77.085 ;
         LAYER metal3 ;
         RECT  53.13 2.47 53.265 2.605 ;
         LAYER metal3 ;
         RECT  206.41 73.96 206.545 74.095 ;
         LAYER metal4 ;
         RECT  26.2075 51.5325 26.3475 243.1025 ;
         LAYER metal4 ;
         RECT  15.8075 33.3325 15.9475 48.2925 ;
         LAYER metal3 ;
         RECT  2.425 33.335 2.56 33.47 ;
         LAYER metal3 ;
         RECT  34.73 255.32 170.32 255.39 ;
         LAYER metal4 ;
         RECT  33.5825 51.5325 33.7225 243.0325 ;
         LAYER metal3 ;
         RECT  33.585 50.04 33.72 50.175 ;
         LAYER metal3 ;
         RECT  20.095 64.99 20.23 65.125 ;
         LAYER metal3 ;
         RECT  20.095 53.03 20.23 53.165 ;
         LAYER metal3 ;
         RECT  224.07 258.445 224.205 258.58 ;
         LAYER metal3 ;
         RECT  41.69 2.47 41.825 2.605 ;
         LAYER metal3 ;
         RECT  206.065 53.03 206.2 53.165 ;
         LAYER metal3 ;
         RECT  34.73 246.6475 189.59 246.7175 ;
         LAYER metal3 ;
         RECT  19.75 79.94 19.885 80.075 ;
         LAYER metal3 ;
         RECT  19.75 70.97 19.885 71.105 ;
         LAYER metal4 ;
         RECT  22.2525 5.685 22.3925 45.345 ;
         LAYER metal3 ;
         RECT  192.575 244.39 192.71 244.525 ;
         LAYER metal4 ;
         RECT  225.8025 228.8025 225.9425 251.205 ;
         LAYER metal4 ;
         RECT  213.2625 34.1775 213.4025 51.6725 ;
         LAYER metal3 ;
         RECT  199.3325 243.6025 199.4675 243.7375 ;
         LAYER metal3 ;
         RECT  204.685 289.46 204.82 289.595 ;
         LAYER metal3 ;
         RECT  188.28 36.49 188.415 36.625 ;
         LAYER metal3 ;
         RECT  19.75 76.95 19.885 77.085 ;
         LAYER metal3 ;
         RECT  206.065 56.02 206.2 56.155 ;
         LAYER metal4 ;
         RECT  191.4925 48.3625 191.6325 245.9525 ;
         LAYER metal3 ;
         RECT  18.81 2.47 18.945 2.605 ;
         LAYER metal3 ;
         RECT  34.595 36.49 34.73 36.625 ;
         LAYER metal4 ;
         RECT  203.9025 249.04 204.0425 288.7 ;
         LAYER metal3 ;
         RECT  206.065 62.0 206.2 62.135 ;
         LAYER metal4 ;
         RECT  210.5425 248.5625 210.6825 258.5825 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  34.595 34.67 34.73 34.805 ;
         LAYER metal3 ;
         RECT  207.5925 51.535 207.7275 51.67 ;
         LAYER metal4 ;
         RECT  6.105 30.8625 6.245 45.8225 ;
         LAYER metal3 ;
         RECT  44.55 0.0 44.685 0.135 ;
         LAYER metal3 ;
         RECT  17.9425 75.455 18.0775 75.59 ;
         LAYER metal4 ;
         RECT  191.0325 48.3625 191.1725 245.9525 ;
         LAYER metal3 ;
         RECT  188.28 34.67 188.415 34.805 ;
         LAYER metal3 ;
         RECT  207.5925 63.495 207.7275 63.63 ;
         LAYER metal3 ;
         RECT  21.67 0.0 21.805 0.135 ;
         LAYER metal3 ;
         RECT  201.825 291.93 201.96 292.065 ;
         LAYER metal4 ;
         RECT  24.2725 51.5 24.4125 243.1025 ;
         LAYER metal3 ;
         RECT  208.2175 69.475 208.3525 69.61 ;
         LAYER metal3 ;
         RECT  18.5675 51.535 18.7025 51.67 ;
         LAYER metal3 ;
         RECT  208.2175 78.445 208.3525 78.58 ;
         LAYER metal3 ;
         RECT  34.73 45.0475 188.4475 45.1175 ;
         LAYER metal3 ;
         RECT  17.9425 78.445 18.0775 78.58 ;
         LAYER metal3 ;
         RECT  207.5925 66.485 207.7275 66.62 ;
         LAYER metal3 ;
         RECT  34.73 253.4275 170.355 253.4975 ;
         LAYER metal3 ;
         RECT  207.5925 54.525 207.7275 54.66 ;
         LAYER metal3 ;
         RECT  34.73 249.2675 188.4475 249.3375 ;
         LAYER metal4 ;
         RECT  26.7675 51.5 26.9075 243.065 ;
         LAYER metal4 ;
         RECT  35.1225 48.3625 35.2625 245.9525 ;
         LAYER metal4 ;
         RECT  220.245 246.0925 220.385 261.0525 ;
         LAYER metal4 ;
         RECT  210.4025 34.2425 210.5425 51.7375 ;
         LAYER metal4 ;
         RECT  199.3875 51.5 199.5275 243.065 ;
         LAYER metal3 ;
         RECT  55.99 0.0 56.125 0.135 ;
         LAYER metal4 ;
         RECT  206.125 248.9725 206.265 288.7675 ;
         LAYER metal3 ;
         RECT  18.5675 60.505 18.7025 60.64 ;
         LAYER metal3 ;
         RECT  17.9425 72.465 18.0775 72.6 ;
         LAYER metal3 ;
         RECT  207.5925 60.505 207.7275 60.64 ;
         LAYER metal3 ;
         RECT  33.11 0.0 33.245 0.135 ;
         LAYER metal3 ;
         RECT  2.425 30.865 2.56 31.0 ;
         LAYER metal3 ;
         RECT  18.5675 66.485 18.7025 66.62 ;
         LAYER metal3 ;
         RECT  208.2175 81.435 208.3525 81.57 ;
         LAYER metal3 ;
         RECT  17.9425 69.475 18.0775 69.61 ;
         LAYER metal3 ;
         RECT  18.5675 63.495 18.7025 63.63 ;
         LAYER metal3 ;
         RECT  18.5675 54.525 18.7025 54.66 ;
         LAYER metal4 ;
         RECT  20.03 5.6175 20.17 45.4125 ;
         LAYER metal4 ;
         RECT  201.8825 51.5 202.0225 243.1025 ;
         LAYER metal3 ;
         RECT  18.5675 57.515 18.7025 57.65 ;
         LAYER metal4 ;
         RECT  15.9475 81.3675 16.0875 98.8625 ;
         LAYER metal3 ;
         RECT  17.9425 81.435 18.0775 81.57 ;
         LAYER metal3 ;
         RECT  224.07 260.915 224.205 261.05 ;
         LAYER metal3 ;
         RECT  207.5925 57.515 207.7275 57.65 ;
         LAYER metal3 ;
         RECT  34.73 39.5075 170.32 39.5775 ;
         LAYER metal4 ;
         RECT  223.74 228.77 223.88 251.1725 ;
         LAYER metal4 ;
         RECT  2.75 40.7425 2.89 63.145 ;
         LAYER metal3 ;
         RECT  208.2175 75.455 208.3525 75.59 ;
         LAYER metal3 ;
         RECT  208.2175 72.465 208.3525 72.6 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 226.49 291.925 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 226.49 291.925 ;
   LAYER  metal3 ;
      RECT  41.8325 0.14 42.2475 0.965 ;
      RECT  42.2475 0.965 44.6925 1.38 ;
      RECT  45.1075 0.965 47.5525 1.38 ;
      RECT  47.9675 0.965 50.4125 1.38 ;
      RECT  50.8275 0.965 53.2725 1.38 ;
      RECT  53.6875 0.965 56.1325 1.38 ;
      RECT  56.5475 0.965 58.9925 1.38 ;
      RECT  59.4075 0.965 61.8525 1.38 ;
      RECT  62.2675 0.965 226.49 1.38 ;
      RECT  0.14 0.965 18.9525 1.38 ;
      RECT  19.3675 0.965 21.8125 1.38 ;
      RECT  22.2275 0.965 24.6725 1.38 ;
      RECT  25.0875 0.965 27.5325 1.38 ;
      RECT  0.14 82.4 13.2325 82.815 ;
      RECT  0.14 82.815 13.2325 291.925 ;
      RECT  13.2325 1.38 13.6475 82.4 ;
      RECT  13.6475 82.4 41.8325 82.815 ;
      RECT  13.2325 82.815 13.6475 85.13 ;
      RECT  13.2325 85.545 13.6475 87.34 ;
      RECT  13.2325 87.755 13.6475 90.07 ;
      RECT  13.2325 90.485 13.6475 92.28 ;
      RECT  13.2325 92.695 13.6475 95.01 ;
      RECT  13.2325 95.425 13.6475 97.22 ;
      RECT  13.2325 97.635 13.6475 291.925 ;
      RECT  204.2625 291.1 204.6775 291.925 ;
      RECT  204.6775 290.685 226.49 291.1 ;
      RECT  204.6775 291.1 226.49 291.925 ;
      RECT  201.8175 290.685 204.2625 291.1 ;
      RECT  198.9575 290.685 201.4025 291.1 ;
      RECT  42.2475 290.685 195.6825 291.1 ;
      RECT  196.0975 290.685 198.5425 291.1 ;
      RECT  204.6775 1.38 212.8425 50.29 ;
      RECT  204.6775 50.29 212.8425 50.705 ;
      RECT  212.8425 50.705 213.2575 290.685 ;
      RECT  213.2575 1.38 226.49 50.29 ;
      RECT  213.2575 50.29 226.49 50.705 ;
      RECT  212.8425 47.975 213.2575 50.29 ;
      RECT  212.8425 45.765 213.2575 47.56 ;
      RECT  212.8425 43.035 213.2575 45.35 ;
      RECT  212.8425 40.825 213.2575 42.62 ;
      RECT  212.8425 38.095 213.2575 40.41 ;
      RECT  212.8425 1.38 213.2575 35.47 ;
      RECT  212.8425 35.885 213.2575 37.68 ;
      RECT  0.14 1.38 0.1475 31.83 ;
      RECT  0.14 31.83 0.1475 32.245 ;
      RECT  0.14 32.245 0.1475 82.4 ;
      RECT  0.1475 1.38 0.5625 31.83 ;
      RECT  0.1475 32.245 0.5625 82.4 ;
      RECT  226.0675 50.705 226.4825 259.67 ;
      RECT  226.0675 260.085 226.4825 290.685 ;
      RECT  226.4825 50.705 226.49 259.67 ;
      RECT  226.4825 259.67 226.49 260.085 ;
      RECT  226.4825 260.085 226.49 290.685 ;
      RECT  0.5625 31.83 6.1075 31.915 ;
      RECT  0.5625 31.915 6.1075 32.245 ;
      RECT  6.1075 31.83 6.5225 31.915 ;
      RECT  6.5225 31.83 13.2325 31.915 ;
      RECT  6.5225 31.915 13.2325 32.245 ;
      RECT  0.5625 32.245 6.1075 32.33 ;
      RECT  6.1075 32.33 6.5225 82.4 ;
      RECT  6.5225 32.245 13.2325 32.33 ;
      RECT  6.5225 32.33 13.2325 82.4 ;
      RECT  213.2575 50.705 219.9675 259.585 ;
      RECT  213.2575 259.585 219.9675 259.67 ;
      RECT  219.9675 50.705 220.3825 259.585 ;
      RECT  220.3825 259.585 226.0675 259.67 ;
      RECT  213.2575 259.67 219.9675 260.0 ;
      RECT  213.2575 260.0 219.9675 260.085 ;
      RECT  219.9675 260.0 220.3825 260.085 ;
      RECT  220.3825 259.67 226.0675 260.0 ;
      RECT  220.3825 260.0 226.0675 260.085 ;
      RECT  27.9475 0.965 30.3925 1.38 ;
      RECT  30.8075 0.965 33.2525 1.38 ;
      RECT  33.6675 0.965 36.1125 1.38 ;
      RECT  36.5275 0.965 38.9725 1.38 ;
      RECT  39.3875 0.965 41.8325 1.38 ;
      RECT  13.6475 257.7375 37.775 258.1525 ;
      RECT  13.6475 258.1525 37.775 291.925 ;
      RECT  37.775 258.1525 38.19 291.925 ;
      RECT  38.19 257.7375 41.8325 258.1525 ;
      RECT  38.19 258.1525 41.8325 291.925 ;
      RECT  42.2475 257.7375 56.575 258.1525 ;
      RECT  42.2475 258.1525 56.575 290.685 ;
      RECT  56.575 258.1525 56.99 290.685 ;
      RECT  56.99 258.1525 204.2625 290.685 ;
      RECT  56.99 257.7375 75.375 258.1525 ;
      RECT  75.79 257.7375 94.175 258.1525 ;
      RECT  94.59 257.7375 112.975 258.1525 ;
      RECT  113.39 257.7375 131.775 258.1525 ;
      RECT  132.19 257.7375 150.575 258.1525 ;
      RECT  150.99 257.7375 169.375 258.1525 ;
      RECT  169.79 257.7375 204.2625 258.1525 ;
      RECT  13.6475 37.3175 34.59 37.6675 ;
      RECT  56.575 1.38 56.99 37.3175 ;
      RECT  56.99 1.38 170.46 37.3175 ;
      RECT  170.46 37.3175 204.2625 37.6675 ;
      RECT  13.6475 37.6675 26.6875 50.6875 ;
      RECT  13.6475 50.6875 26.6875 51.1025 ;
      RECT  26.6875 37.6675 27.1025 50.6875 ;
      RECT  26.6875 51.1025 27.1025 82.4 ;
      RECT  27.1025 50.6875 34.59 51.1025 ;
      RECT  27.1025 51.1025 34.59 82.4 ;
      RECT  204.6775 50.705 205.925 64.85 ;
      RECT  204.6775 64.85 205.925 65.265 ;
      RECT  206.34 64.85 212.8425 65.265 ;
      RECT  13.6475 55.88 19.955 56.295 ;
      RECT  20.37 51.1025 26.6875 55.88 ;
      RECT  20.37 55.88 26.6875 56.295 ;
      RECT  20.37 56.295 26.6875 82.4 ;
      RECT  34.59 47.8775 41.8325 82.4 ;
      RECT  188.555 47.5275 204.2625 47.8775 ;
      RECT  19.955 56.295 20.37 61.86 ;
      RECT  13.6475 73.82 19.61 74.235 ;
      RECT  20.025 73.82 20.37 74.235 ;
      RECT  20.025 74.235 20.37 82.4 ;
      RECT  13.6475 1.38 30.11 2.33 ;
      RECT  13.6475 2.745 30.11 37.3175 ;
      RECT  30.11 1.38 30.525 2.33 ;
      RECT  30.11 2.745 30.525 37.3175 ;
      RECT  30.525 1.38 34.59 2.33 ;
      RECT  30.525 2.33 34.59 2.745 ;
      RECT  205.925 65.265 206.27 70.83 ;
      RECT  205.925 70.83 206.27 71.245 ;
      RECT  205.925 71.245 206.27 290.685 ;
      RECT  206.27 65.265 206.34 70.83 ;
      RECT  206.34 65.265 206.685 70.83 ;
      RECT  206.685 70.83 212.8425 71.245 ;
      RECT  206.27 80.215 206.34 290.685 ;
      RECT  206.34 80.215 206.685 290.685 ;
      RECT  206.27 77.225 206.34 79.8 ;
      RECT  206.34 77.225 206.685 79.8 ;
      RECT  42.2475 1.38 52.99 2.33 ;
      RECT  42.2475 2.33 52.99 2.745 ;
      RECT  42.2475 2.745 52.99 37.3175 ;
      RECT  52.99 1.38 53.405 2.33 ;
      RECT  52.99 2.745 53.405 37.3175 ;
      RECT  53.405 1.38 56.575 2.33 ;
      RECT  53.405 2.33 56.575 2.745 ;
      RECT  53.405 2.745 56.575 37.3175 ;
      RECT  206.27 71.245 206.34 73.82 ;
      RECT  206.27 74.235 206.34 76.81 ;
      RECT  206.34 71.245 206.685 73.82 ;
      RECT  206.34 74.235 206.685 76.81 ;
      RECT  0.5625 32.33 2.285 33.195 ;
      RECT  0.5625 33.195 2.285 33.61 ;
      RECT  0.5625 33.61 2.285 82.4 ;
      RECT  2.285 32.33 2.7 33.195 ;
      RECT  2.285 33.61 2.7 82.4 ;
      RECT  2.7 32.33 6.1075 33.195 ;
      RECT  2.7 33.195 6.1075 33.61 ;
      RECT  2.7 33.61 6.1075 82.4 ;
      RECT  13.6475 82.815 34.59 255.18 ;
      RECT  13.6475 255.18 34.59 255.53 ;
      RECT  13.6475 255.53 34.59 257.7375 ;
      RECT  34.59 255.53 37.775 257.7375 ;
      RECT  37.775 255.53 38.19 257.7375 ;
      RECT  38.19 255.53 41.8325 257.7375 ;
      RECT  41.8325 255.53 42.2475 291.925 ;
      RECT  42.2475 255.53 56.575 257.7375 ;
      RECT  56.575 255.53 56.99 257.7375 ;
      RECT  56.99 255.53 170.46 257.7375 ;
      RECT  27.1025 37.6675 33.445 49.9 ;
      RECT  27.1025 49.9 33.445 50.315 ;
      RECT  27.1025 50.315 33.445 50.6875 ;
      RECT  33.445 37.6675 33.86 49.9 ;
      RECT  33.445 50.315 33.86 50.6875 ;
      RECT  33.86 37.6675 34.59 49.9 ;
      RECT  33.86 49.9 34.59 50.315 ;
      RECT  33.86 50.315 34.59 50.6875 ;
      RECT  19.955 62.275 20.025 64.85 ;
      RECT  20.025 62.275 20.37 64.85 ;
      RECT  20.025 65.265 20.37 73.82 ;
      RECT  19.955 51.1025 20.37 52.89 ;
      RECT  19.955 53.305 20.37 55.88 ;
      RECT  220.3825 50.705 223.93 258.305 ;
      RECT  220.3825 258.305 223.93 258.72 ;
      RECT  220.3825 258.72 223.93 259.585 ;
      RECT  223.93 50.705 224.345 258.305 ;
      RECT  223.93 258.72 224.345 259.585 ;
      RECT  224.345 50.705 226.0675 258.305 ;
      RECT  224.345 258.305 226.0675 258.72 ;
      RECT  224.345 258.72 226.0675 259.585 ;
      RECT  41.8325 1.38 41.965 2.33 ;
      RECT  41.8325 2.745 41.965 37.3175 ;
      RECT  41.965 1.38 42.2475 2.33 ;
      RECT  41.965 2.33 42.2475 2.745 ;
      RECT  41.965 2.745 42.2475 37.3175 ;
      RECT  34.59 1.38 41.55 2.33 ;
      RECT  34.59 2.33 41.55 2.745 ;
      RECT  41.55 1.38 41.8325 2.33 ;
      RECT  41.55 2.745 41.8325 37.3175 ;
      RECT  205.925 50.705 206.34 52.89 ;
      RECT  170.46 47.8775 188.555 246.5075 ;
      RECT  188.555 47.8775 189.73 246.5075 ;
      RECT  189.73 246.5075 204.2625 246.8575 ;
      RECT  189.73 246.8575 204.2625 257.7375 ;
      RECT  34.59 82.815 37.775 246.5075 ;
      RECT  37.775 82.815 38.19 246.5075 ;
      RECT  38.19 82.815 41.8325 246.5075 ;
      RECT  41.8325 47.8775 42.2475 246.5075 ;
      RECT  42.2475 47.8775 56.575 246.5075 ;
      RECT  56.575 47.8775 56.99 246.5075 ;
      RECT  56.99 47.8775 170.46 246.5075 ;
      RECT  19.61 80.215 19.955 82.4 ;
      RECT  19.955 80.215 20.025 82.4 ;
      RECT  19.61 56.295 19.955 70.83 ;
      RECT  19.61 71.245 19.955 73.82 ;
      RECT  19.955 65.265 20.025 70.83 ;
      RECT  19.955 71.245 20.025 73.82 ;
      RECT  189.73 47.8775 192.435 244.25 ;
      RECT  189.73 244.25 192.435 244.665 ;
      RECT  189.73 244.665 192.435 246.5075 ;
      RECT  192.435 47.8775 192.85 244.25 ;
      RECT  192.435 244.665 192.85 246.5075 ;
      RECT  192.85 244.25 204.2625 244.665 ;
      RECT  192.85 244.665 204.2625 246.5075 ;
      RECT  192.85 47.8775 199.1925 243.4625 ;
      RECT  192.85 243.4625 199.1925 243.8775 ;
      RECT  192.85 243.8775 199.1925 244.25 ;
      RECT  199.1925 47.8775 199.6075 243.4625 ;
      RECT  199.1925 243.8775 199.6075 244.25 ;
      RECT  199.6075 47.8775 204.2625 243.4625 ;
      RECT  199.6075 243.4625 204.2625 243.8775 ;
      RECT  199.6075 243.8775 204.2625 244.25 ;
      RECT  204.2625 1.38 204.545 289.32 ;
      RECT  204.2625 289.32 204.545 289.735 ;
      RECT  204.2625 289.735 204.545 290.685 ;
      RECT  204.545 1.38 204.6775 289.32 ;
      RECT  204.545 289.735 204.6775 290.685 ;
      RECT  204.6775 65.265 204.96 289.32 ;
      RECT  204.6775 289.735 204.96 290.685 ;
      RECT  204.96 65.265 205.925 289.32 ;
      RECT  204.96 289.32 205.925 289.735 ;
      RECT  204.96 289.735 205.925 290.685 ;
      RECT  170.46 1.38 188.14 36.35 ;
      RECT  170.46 36.35 188.14 36.765 ;
      RECT  170.46 36.765 188.14 37.3175 ;
      RECT  188.14 36.765 188.555 37.3175 ;
      RECT  188.555 1.38 204.2625 36.35 ;
      RECT  188.555 36.35 204.2625 36.765 ;
      RECT  188.555 36.765 204.2625 37.3175 ;
      RECT  19.61 74.235 19.955 76.81 ;
      RECT  19.61 77.225 19.955 79.8 ;
      RECT  19.955 74.235 20.025 76.81 ;
      RECT  19.955 77.225 20.025 79.8 ;
      RECT  205.925 53.305 206.34 55.88 ;
      RECT  13.6475 2.33 18.67 2.745 ;
      RECT  19.085 2.33 30.11 2.745 ;
      RECT  30.525 2.745 34.455 36.35 ;
      RECT  30.525 36.35 34.455 36.765 ;
      RECT  30.525 36.765 34.455 37.3175 ;
      RECT  34.455 36.765 34.59 37.3175 ;
      RECT  34.59 36.765 34.87 37.3175 ;
      RECT  34.87 2.745 41.55 36.35 ;
      RECT  34.87 36.35 41.55 36.765 ;
      RECT  34.87 36.765 41.55 37.3175 ;
      RECT  205.925 56.295 206.34 61.86 ;
      RECT  205.925 62.275 206.34 64.85 ;
      RECT  34.455 2.745 34.59 34.53 ;
      RECT  34.455 34.945 34.59 36.35 ;
      RECT  34.59 2.745 34.87 34.53 ;
      RECT  34.59 34.945 34.87 36.35 ;
      RECT  206.34 50.705 207.4525 51.395 ;
      RECT  206.34 51.395 207.4525 51.81 ;
      RECT  206.34 51.81 207.4525 64.85 ;
      RECT  207.4525 50.705 207.8675 51.395 ;
      RECT  207.8675 50.705 212.8425 51.395 ;
      RECT  207.8675 51.395 212.8425 51.81 ;
      RECT  207.8675 51.81 212.8425 64.85 ;
      RECT  42.2475 0.14 44.41 0.275 ;
      RECT  42.2475 0.275 44.41 0.965 ;
      RECT  44.41 0.275 44.825 0.965 ;
      RECT  44.825 0.275 226.49 0.965 ;
      RECT  13.6475 74.235 17.8025 75.315 ;
      RECT  13.6475 75.315 17.8025 75.73 ;
      RECT  13.6475 75.73 17.8025 82.4 ;
      RECT  17.8025 74.235 18.2175 75.315 ;
      RECT  18.2175 74.235 19.61 75.315 ;
      RECT  18.2175 75.315 19.61 75.73 ;
      RECT  18.2175 75.73 19.61 82.4 ;
      RECT  188.14 1.38 188.555 34.53 ;
      RECT  188.14 34.945 188.555 36.35 ;
      RECT  207.4525 63.77 207.8675 64.85 ;
      RECT  0.14 0.14 21.53 0.275 ;
      RECT  0.14 0.275 21.53 0.965 ;
      RECT  21.53 0.275 21.945 0.965 ;
      RECT  21.945 0.275 41.8325 0.965 ;
      RECT  42.2475 291.1 201.685 291.79 ;
      RECT  42.2475 291.79 201.685 291.925 ;
      RECT  201.685 291.1 202.1 291.79 ;
      RECT  202.1 291.1 204.2625 291.79 ;
      RECT  202.1 291.79 204.2625 291.925 ;
      RECT  206.685 69.335 208.0775 69.75 ;
      RECT  206.685 69.75 208.0775 70.83 ;
      RECT  208.0775 65.265 208.4925 69.335 ;
      RECT  208.0775 69.75 208.4925 70.83 ;
      RECT  208.4925 65.265 212.8425 69.335 ;
      RECT  208.4925 69.335 212.8425 69.75 ;
      RECT  208.4925 69.75 212.8425 70.83 ;
      RECT  13.6475 51.1025 18.4275 51.395 ;
      RECT  13.6475 51.395 18.4275 51.81 ;
      RECT  13.6475 51.81 18.4275 55.88 ;
      RECT  18.4275 51.1025 18.8425 51.395 ;
      RECT  18.8425 51.1025 19.955 51.395 ;
      RECT  18.8425 51.395 19.955 51.81 ;
      RECT  18.8425 51.81 19.955 55.88 ;
      RECT  206.685 71.245 208.0775 78.305 ;
      RECT  206.685 78.305 208.0775 78.72 ;
      RECT  206.685 78.72 208.0775 290.685 ;
      RECT  208.4925 71.245 212.8425 78.305 ;
      RECT  208.4925 78.305 212.8425 78.72 ;
      RECT  208.4925 78.72 212.8425 290.685 ;
      RECT  41.8325 45.2575 42.2475 47.5275 ;
      RECT  34.59 45.2575 41.8325 47.5275 ;
      RECT  42.2475 45.2575 56.575 47.5275 ;
      RECT  56.575 45.2575 56.99 47.5275 ;
      RECT  56.99 45.2575 170.46 47.5275 ;
      RECT  170.46 37.6675 188.555 44.9075 ;
      RECT  170.46 45.2575 188.555 47.5275 ;
      RECT  188.555 37.6675 188.5875 44.9075 ;
      RECT  188.555 45.2575 188.5875 47.5275 ;
      RECT  188.5875 37.6675 204.2625 44.9075 ;
      RECT  188.5875 44.9075 204.2625 45.2575 ;
      RECT  188.5875 45.2575 204.2625 47.5275 ;
      RECT  17.8025 75.73 18.2175 78.305 ;
      RECT  206.685 65.265 207.4525 66.345 ;
      RECT  206.685 66.345 207.4525 66.76 ;
      RECT  206.685 66.76 207.4525 69.335 ;
      RECT  207.4525 65.265 207.8675 66.345 ;
      RECT  207.4525 66.76 207.8675 69.335 ;
      RECT  207.8675 65.265 208.0775 66.345 ;
      RECT  207.8675 66.345 208.0775 66.76 ;
      RECT  207.8675 66.76 208.0775 69.335 ;
      RECT  170.46 253.6375 170.495 257.7375 ;
      RECT  170.495 253.2875 188.555 253.6375 ;
      RECT  170.495 253.6375 188.555 257.7375 ;
      RECT  34.59 253.6375 37.775 255.18 ;
      RECT  37.775 253.6375 38.19 255.18 ;
      RECT  38.19 253.6375 41.8325 255.18 ;
      RECT  41.8325 253.6375 42.2475 255.18 ;
      RECT  42.2475 253.6375 56.575 255.18 ;
      RECT  56.575 253.6375 56.99 255.18 ;
      RECT  56.99 253.6375 170.46 255.18 ;
      RECT  207.4525 51.81 207.8675 54.385 ;
      RECT  188.555 246.8575 188.5875 249.1275 ;
      RECT  188.555 249.4775 188.5875 257.7375 ;
      RECT  188.5875 246.8575 189.73 249.1275 ;
      RECT  188.5875 249.1275 189.73 249.4775 ;
      RECT  188.5875 249.4775 189.73 257.7375 ;
      RECT  170.46 246.8575 170.495 249.1275 ;
      RECT  170.46 249.4775 170.495 253.2875 ;
      RECT  170.495 246.8575 188.555 249.1275 ;
      RECT  170.495 249.4775 188.555 253.2875 ;
      RECT  34.59 246.8575 37.775 249.1275 ;
      RECT  34.59 249.4775 37.775 253.2875 ;
      RECT  37.775 246.8575 38.19 249.1275 ;
      RECT  37.775 249.4775 38.19 253.2875 ;
      RECT  38.19 246.8575 41.8325 249.1275 ;
      RECT  38.19 249.4775 41.8325 253.2875 ;
      RECT  41.8325 246.8575 42.2475 249.1275 ;
      RECT  41.8325 249.4775 42.2475 253.2875 ;
      RECT  42.2475 246.8575 56.575 249.1275 ;
      RECT  42.2475 249.4775 56.575 253.2875 ;
      RECT  56.575 246.8575 56.99 249.1275 ;
      RECT  56.575 249.4775 56.99 253.2875 ;
      RECT  56.99 246.8575 170.46 249.1275 ;
      RECT  56.99 249.4775 170.46 253.2875 ;
      RECT  44.825 0.14 55.85 0.275 ;
      RECT  56.265 0.14 226.49 0.275 ;
      RECT  13.6475 56.295 18.4275 60.365 ;
      RECT  13.6475 60.365 18.4275 60.78 ;
      RECT  18.8425 56.295 19.61 60.365 ;
      RECT  18.8425 60.365 19.61 60.78 ;
      RECT  18.8425 60.78 19.61 73.82 ;
      RECT  13.6475 60.78 17.8025 72.325 ;
      RECT  13.6475 72.325 17.8025 72.74 ;
      RECT  13.6475 72.74 17.8025 73.82 ;
      RECT  17.8025 72.74 18.2175 73.82 ;
      RECT  18.2175 60.78 18.4275 72.325 ;
      RECT  18.2175 72.325 18.4275 72.74 ;
      RECT  18.2175 72.74 18.4275 73.82 ;
      RECT  207.4525 60.78 207.8675 63.355 ;
      RECT  21.945 0.14 32.97 0.275 ;
      RECT  33.385 0.14 41.8325 0.275 ;
      RECT  0.5625 1.38 2.285 30.725 ;
      RECT  0.5625 30.725 2.285 31.14 ;
      RECT  0.5625 31.14 2.285 31.83 ;
      RECT  2.285 1.38 2.7 30.725 ;
      RECT  2.285 31.14 2.7 31.83 ;
      RECT  2.7 1.38 13.2325 30.725 ;
      RECT  2.7 30.725 13.2325 31.14 ;
      RECT  2.7 31.14 13.2325 31.83 ;
      RECT  18.4275 66.76 18.8425 73.82 ;
      RECT  208.0775 78.72 208.4925 81.295 ;
      RECT  208.0775 81.71 208.4925 290.685 ;
      RECT  17.8025 60.78 18.2175 69.335 ;
      RECT  17.8025 69.75 18.2175 72.325 ;
      RECT  18.4275 60.78 18.8425 63.355 ;
      RECT  18.4275 63.77 18.8425 66.345 ;
      RECT  18.4275 51.81 18.8425 54.385 ;
      RECT  18.4275 54.8 18.8425 55.88 ;
      RECT  18.4275 56.295 18.8425 57.375 ;
      RECT  18.4275 57.79 18.8425 60.365 ;
      RECT  17.8025 78.72 18.2175 81.295 ;
      RECT  17.8025 81.71 18.2175 82.4 ;
      RECT  213.2575 260.085 223.93 260.775 ;
      RECT  213.2575 260.775 223.93 261.19 ;
      RECT  213.2575 261.19 223.93 290.685 ;
      RECT  223.93 260.085 224.345 260.775 ;
      RECT  223.93 261.19 224.345 290.685 ;
      RECT  224.345 260.085 226.0675 260.775 ;
      RECT  224.345 260.775 226.0675 261.19 ;
      RECT  224.345 261.19 226.0675 290.685 ;
      RECT  207.4525 54.8 207.8675 57.375 ;
      RECT  207.4525 57.79 207.8675 60.365 ;
      RECT  41.8325 37.6675 42.2475 39.3675 ;
      RECT  41.8325 39.7175 42.2475 44.9075 ;
      RECT  34.59 37.6675 41.8325 39.3675 ;
      RECT  34.59 39.7175 41.8325 44.9075 ;
      RECT  42.2475 37.6675 56.575 39.3675 ;
      RECT  42.2475 39.7175 56.575 44.9075 ;
      RECT  56.575 37.6675 56.99 39.3675 ;
      RECT  56.575 39.7175 56.99 44.9075 ;
      RECT  56.99 37.6675 170.46 39.3675 ;
      RECT  56.99 39.7175 170.46 44.9075 ;
      RECT  208.0775 75.73 208.4925 78.305 ;
      RECT  208.0775 71.245 208.4925 72.325 ;
      RECT  208.0775 72.74 208.4925 75.315 ;
   LAYER  metal4 ;
      RECT  199.6675 243.3825 200.3675 291.925 ;
      RECT  0.14 0.14 0.4075 40.43 ;
      RECT  0.14 40.43 0.4075 51.2525 ;
      RECT  0.4075 0.14 1.1075 40.43 ;
      RECT  0.14 51.2525 0.4075 63.3925 ;
      RECT  0.14 63.3925 0.4075 243.3825 ;
      RECT  0.4075 63.3925 1.1075 243.3825 ;
      RECT  1.1075 81.1525 12.8075 99.2075 ;
      RECT  1.1075 99.2075 12.8075 243.3825 ;
      RECT  12.8075 63.3925 13.5075 81.1525 ;
      RECT  12.8075 99.2075 13.5075 243.3825 ;
      RECT  0.14 243.3825 34.3825 246.2325 ;
      RECT  0.14 246.2325 34.3825 291.925 ;
      RECT  34.3825 246.2325 35.0825 291.925 ;
      RECT  35.0825 246.2325 199.6675 291.925 ;
      RECT  34.3825 40.43 35.0825 48.0825 ;
      RECT  35.0825 40.43 199.6675 48.0825 ;
      RECT  192.2925 243.3125 192.9925 243.3825 ;
      RECT  15.5275 0.14 16.2275 33.0525 ;
      RECT  15.5275 48.5725 16.2275 51.2525 ;
      RECT  16.2275 48.0825 34.3825 48.5725 ;
      RECT  34.0025 51.2525 34.3825 63.3925 ;
      RECT  34.0025 63.3925 34.3825 81.1525 ;
      RECT  34.0025 81.1525 34.3825 99.2075 ;
      RECT  33.3025 243.3125 34.0025 243.3825 ;
      RECT  34.0025 99.2075 34.3825 243.3125 ;
      RECT  34.0025 243.3125 34.3825 243.3825 ;
      RECT  21.9725 0.14 22.6725 5.405 ;
      RECT  22.6725 0.14 199.6675 5.405 ;
      RECT  22.6725 5.405 199.6675 33.0525 ;
      RECT  22.6725 33.0525 199.6675 40.43 ;
      RECT  21.9725 45.625 22.6725 48.0825 ;
      RECT  22.6725 40.43 34.3825 45.625 ;
      RECT  22.6725 45.625 34.3825 48.0825 ;
      RECT  225.5225 51.2525 226.2225 228.5225 ;
      RECT  226.2225 51.2525 226.49 228.5225 ;
      RECT  226.2225 228.5225 226.49 243.3825 ;
      RECT  225.5225 251.485 226.2225 291.925 ;
      RECT  226.2225 243.3825 226.49 251.485 ;
      RECT  226.2225 251.485 226.49 291.925 ;
      RECT  200.3675 0.14 212.9825 33.8975 ;
      RECT  212.9825 0.14 213.6825 33.8975 ;
      RECT  213.6825 0.14 226.49 33.8975 ;
      RECT  213.6825 33.8975 226.49 51.2525 ;
      RECT  212.9825 51.9525 213.6825 228.5225 ;
      RECT  213.6825 51.2525 225.5225 51.9525 ;
      RECT  191.9125 243.3825 199.6675 246.2325 ;
      RECT  191.9125 51.2525 192.2925 63.3925 ;
      RECT  191.9125 63.3925 192.2925 81.1525 ;
      RECT  191.9125 81.1525 192.2925 99.2075 ;
      RECT  191.9125 99.2075 192.2925 243.3125 ;
      RECT  191.9125 243.3125 192.2925 243.3825 ;
      RECT  200.3675 243.3825 203.6225 248.76 ;
      RECT  200.3675 248.76 203.6225 251.485 ;
      RECT  203.6225 243.3825 204.3225 248.76 ;
      RECT  200.3675 251.485 203.6225 288.98 ;
      RECT  200.3675 288.98 203.6225 291.925 ;
      RECT  203.6225 288.98 204.3225 291.925 ;
      RECT  204.3225 243.3825 210.2625 248.2825 ;
      RECT  210.2625 243.3825 210.9625 248.2825 ;
      RECT  210.2625 258.8625 210.9625 288.98 ;
      RECT  1.1075 0.14 5.825 30.5825 ;
      RECT  1.1075 30.5825 5.825 33.0525 ;
      RECT  5.825 0.14 6.525 30.5825 ;
      RECT  6.525 0.14 15.5275 30.5825 ;
      RECT  6.525 30.5825 15.5275 33.0525 ;
      RECT  1.1075 33.0525 5.825 40.43 ;
      RECT  6.525 33.0525 15.5275 40.43 ;
      RECT  5.825 46.1025 6.525 48.0825 ;
      RECT  6.525 40.43 15.5275 46.1025 ;
      RECT  6.525 46.1025 15.5275 48.0825 ;
      RECT  24.6925 51.2525 25.9275 63.3925 ;
      RECT  24.6925 63.3925 25.9275 81.1525 ;
      RECT  24.6925 81.1525 25.9275 99.2075 ;
      RECT  13.5075 99.2075 23.9925 243.3825 ;
      RECT  24.6925 99.2075 25.9275 243.3825 ;
      RECT  16.2275 48.5725 23.9925 51.22 ;
      RECT  16.2275 51.22 23.9925 51.2525 ;
      RECT  23.9925 48.5725 24.6925 51.22 ;
      RECT  24.6925 48.5725 34.3825 51.22 ;
      RECT  27.1875 51.2525 33.3025 63.3925 ;
      RECT  27.1875 63.3925 33.3025 81.1525 ;
      RECT  27.1875 81.1525 33.3025 99.2075 ;
      RECT  27.1875 99.2075 33.3025 243.3125 ;
      RECT  26.6275 243.345 27.1875 243.3825 ;
      RECT  27.1875 243.3125 33.3025 243.345 ;
      RECT  27.1875 243.345 33.3025 243.3825 ;
      RECT  24.6925 51.22 26.4875 51.2525 ;
      RECT  27.1875 51.22 34.3825 51.2525 ;
      RECT  35.5425 243.3825 190.7525 246.2325 ;
      RECT  35.5425 48.0825 190.7525 51.2525 ;
      RECT  35.5425 51.2525 190.7525 63.3925 ;
      RECT  35.5425 63.3925 190.7525 81.1525 ;
      RECT  35.5425 81.1525 190.7525 99.2075 ;
      RECT  35.5425 99.2075 190.7525 243.3125 ;
      RECT  35.5425 243.3125 190.7525 243.3825 ;
      RECT  210.9625 243.3825 219.965 245.8125 ;
      RECT  210.9625 245.8125 219.965 248.2825 ;
      RECT  219.965 243.3825 220.665 245.8125 ;
      RECT  210.9625 248.2825 219.965 248.76 ;
      RECT  210.9625 248.76 219.965 251.485 ;
      RECT  210.9625 251.485 219.965 258.8625 ;
      RECT  220.665 251.485 225.5225 258.8625 ;
      RECT  210.9625 258.8625 219.965 261.3325 ;
      RECT  210.9625 261.3325 219.965 288.98 ;
      RECT  219.965 261.3325 220.665 288.98 ;
      RECT  220.665 258.8625 225.5225 261.3325 ;
      RECT  220.665 261.3325 225.5225 288.98 ;
      RECT  200.3675 33.8975 210.1225 33.9625 ;
      RECT  210.1225 33.8975 210.8225 33.9625 ;
      RECT  210.8225 33.8975 212.9825 33.9625 ;
      RECT  210.8225 33.9625 212.9825 51.2525 ;
      RECT  210.8225 51.2525 212.9825 51.9525 ;
      RECT  210.1225 52.0175 210.8225 228.5225 ;
      RECT  210.8225 51.9525 212.9825 52.0175 ;
      RECT  210.8225 52.0175 212.9825 228.5225 ;
      RECT  199.6675 0.14 199.8075 51.22 ;
      RECT  199.8075 0.14 200.3675 51.22 ;
      RECT  199.8075 51.22 200.3675 51.2525 ;
      RECT  192.9925 51.2525 199.1075 63.3925 ;
      RECT  192.9925 63.3925 199.1075 81.1525 ;
      RECT  192.9925 81.1525 199.1075 99.2075 ;
      RECT  192.9925 99.2075 199.1075 243.3125 ;
      RECT  192.9925 243.3125 199.1075 243.345 ;
      RECT  192.9925 243.345 199.1075 243.3825 ;
      RECT  199.1075 243.345 199.6675 243.3825 ;
      RECT  191.9125 48.0825 199.1075 51.22 ;
      RECT  191.9125 51.22 199.1075 51.2525 ;
      RECT  199.1075 48.0825 199.6675 51.22 ;
      RECT  204.3225 288.98 205.845 289.0475 ;
      RECT  204.3225 289.0475 205.845 291.925 ;
      RECT  205.845 289.0475 206.545 291.925 ;
      RECT  206.545 288.98 225.5225 289.0475 ;
      RECT  206.545 289.0475 225.5225 291.925 ;
      RECT  204.3225 248.2825 205.845 248.6925 ;
      RECT  204.3225 248.6925 205.845 248.76 ;
      RECT  205.845 248.2825 206.545 248.6925 ;
      RECT  206.545 248.2825 210.2625 248.6925 ;
      RECT  206.545 248.6925 210.2625 248.76 ;
      RECT  204.3225 248.76 205.845 251.485 ;
      RECT  206.545 248.76 210.2625 251.485 ;
      RECT  204.3225 251.485 205.845 258.8625 ;
      RECT  206.545 251.485 210.2625 258.8625 ;
      RECT  204.3225 258.8625 205.845 288.98 ;
      RECT  206.545 258.8625 210.2625 288.98 ;
      RECT  16.2275 0.14 19.75 5.3375 ;
      RECT  16.2275 5.3375 19.75 5.405 ;
      RECT  19.75 0.14 20.45 5.3375 ;
      RECT  20.45 0.14 21.9725 5.3375 ;
      RECT  20.45 5.3375 21.9725 5.405 ;
      RECT  16.2275 5.405 19.75 33.0525 ;
      RECT  20.45 5.405 21.9725 33.0525 ;
      RECT  16.2275 33.0525 19.75 40.43 ;
      RECT  20.45 33.0525 21.9725 40.43 ;
      RECT  16.2275 40.43 19.75 45.625 ;
      RECT  20.45 40.43 21.9725 45.625 ;
      RECT  16.2275 45.625 19.75 45.6925 ;
      RECT  16.2275 45.6925 19.75 48.0825 ;
      RECT  19.75 45.6925 20.45 48.0825 ;
      RECT  20.45 45.625 21.9725 45.6925 ;
      RECT  20.45 45.6925 21.9725 48.0825 ;
      RECT  200.3675 228.5225 201.6025 243.3825 ;
      RECT  200.3675 33.9625 201.6025 51.22 ;
      RECT  200.3675 51.22 201.6025 51.2525 ;
      RECT  201.6025 33.9625 202.3025 51.22 ;
      RECT  202.3025 33.9625 210.1225 51.22 ;
      RECT  202.3025 51.22 210.1225 51.2525 ;
      RECT  200.3675 51.2525 201.6025 51.9525 ;
      RECT  202.3025 51.2525 210.1225 51.9525 ;
      RECT  200.3675 51.9525 201.6025 52.0175 ;
      RECT  202.3025 51.9525 210.1225 52.0175 ;
      RECT  200.3675 52.0175 201.6025 228.5225 ;
      RECT  202.3025 52.0175 210.1225 228.5225 ;
      RECT  13.5075 63.3925 15.6675 81.0875 ;
      RECT  13.5075 81.0875 15.6675 81.1525 ;
      RECT  15.6675 63.3925 16.3675 81.0875 ;
      RECT  16.3675 63.3925 23.9925 81.0875 ;
      RECT  16.3675 81.0875 23.9925 81.1525 ;
      RECT  13.5075 81.1525 15.6675 99.1425 ;
      RECT  13.5075 99.1425 15.6675 99.2075 ;
      RECT  15.6675 99.1425 16.3675 99.2075 ;
      RECT  16.3675 81.1525 23.9925 99.1425 ;
      RECT  16.3675 99.1425 23.9925 99.2075 ;
      RECT  213.6825 51.9525 223.46 228.49 ;
      RECT  213.6825 228.49 223.46 228.5225 ;
      RECT  223.46 51.9525 224.16 228.49 ;
      RECT  224.16 51.9525 225.5225 228.49 ;
      RECT  224.16 228.49 225.5225 228.5225 ;
      RECT  220.665 243.3825 223.46 245.8125 ;
      RECT  224.16 243.3825 225.5225 245.8125 ;
      RECT  220.665 245.8125 223.46 248.2825 ;
      RECT  224.16 245.8125 225.5225 248.2825 ;
      RECT  220.665 248.2825 223.46 248.76 ;
      RECT  224.16 248.2825 225.5225 248.76 ;
      RECT  220.665 248.76 223.46 251.4525 ;
      RECT  220.665 251.4525 223.46 251.485 ;
      RECT  223.46 251.4525 224.16 251.485 ;
      RECT  224.16 248.76 225.5225 251.4525 ;
      RECT  224.16 251.4525 225.5225 251.485 ;
      RECT  202.3025 228.5225 223.46 243.3825 ;
      RECT  224.16 228.5225 225.5225 243.3825 ;
      RECT  1.1075 63.3925 2.47 63.425 ;
      RECT  1.1075 63.425 2.47 81.1525 ;
      RECT  2.47 63.425 3.17 81.1525 ;
      RECT  3.17 63.3925 12.8075 63.425 ;
      RECT  3.17 63.425 12.8075 81.1525 ;
      RECT  1.1075 48.0825 2.47 48.5725 ;
      RECT  3.17 48.0825 15.5275 48.5725 ;
      RECT  1.1075 48.5725 2.47 51.2525 ;
      RECT  3.17 48.5725 15.5275 51.2525 ;
      RECT  1.1075 40.43 2.47 40.4625 ;
      RECT  1.1075 40.4625 2.47 46.1025 ;
      RECT  2.47 40.43 3.17 40.4625 ;
      RECT  3.17 40.43 5.825 40.4625 ;
      RECT  3.17 40.4625 5.825 46.1025 ;
      RECT  1.1075 46.1025 2.47 48.0825 ;
      RECT  3.17 46.1025 5.825 48.0825 ;
      RECT  1.1075 51.2525 2.47 63.3925 ;
      RECT  3.17 51.2525 23.9925 63.3925 ;
   END
END    freepdk45_sram_1w1r_2048x8_2
END    LIBRARY
