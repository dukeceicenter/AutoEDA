../macros/freepdk45_sram_1w1r_128x120_30/freepdk45_sram_1w1r_128x120_30.lef