../macros/freepdk45_sram_1w1r_16x120/freepdk45_sram_1w1r_16x120.lef