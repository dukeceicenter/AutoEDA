VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_96x32_32
   CLASS BLOCK ;
   SIZE 147.245 BY 110.59 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.075 1.1075 24.21 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.935 1.1075 27.07 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.795 1.1075 29.93 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.655 1.1075 32.79 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.515 1.1075 35.65 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.375 1.1075 38.51 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.235 1.1075 41.37 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.095 1.1075 44.23 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.955 1.1075 47.09 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.815 1.1075 49.95 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.675 1.1075 52.81 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.535 1.1075 55.67 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.395 1.1075 58.53 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.255 1.1075 61.39 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.115 1.1075 64.25 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.975 1.1075 67.11 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.835 1.1075 69.97 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.695 1.1075 72.83 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.555 1.1075 75.69 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.415 1.1075 78.55 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.275 1.1075 81.41 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.135 1.1075 84.27 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.995 1.1075 87.13 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.855 1.1075 89.99 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.715 1.1075 92.85 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.575 1.1075 95.71 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.435 1.1075 98.57 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.295 1.1075 101.43 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.155 1.1075 104.29 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.015 1.1075 107.15 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.875 1.1075 110.01 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.735 1.1075 112.87 1.2425 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.215 1.1075 21.35 1.2425 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 45.6975 15.63 45.8325 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 48.4275 15.63 48.5625 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 50.6375 15.63 50.7725 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 53.3675 15.63 53.5025 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 55.5775 15.63 55.7125 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.495 58.3075 15.63 58.4425 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.895 108.0825 123.03 108.2175 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 19.5675 131.61 19.7025 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 16.8375 131.61 16.9725 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 14.6275 131.61 14.7625 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 11.8975 131.61 12.0325 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 9.6875 131.61 9.8225 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.475 6.9575 131.61 7.0925 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.825 109.3475 146.96 109.4825 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.7225 109.2625 140.8575 109.3975 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.8225 105.595 35.9575 105.73 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.1725 105.595 38.3075 105.73 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.5225 105.595 40.6575 105.73 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.8725 105.595 43.0075 105.73 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.2225 105.595 45.3575 105.73 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.5725 105.595 47.7075 105.73 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.9225 105.595 50.0575 105.73 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.2725 105.595 52.4075 105.73 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.6225 105.595 54.7575 105.73 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.9725 105.595 57.1075 105.73 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.3225 105.595 59.4575 105.73 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.6725 105.595 61.8075 105.73 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.0225 105.595 64.1575 105.73 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.3725 105.595 66.5075 105.73 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.7225 105.595 68.8575 105.73 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.0725 105.595 71.2075 105.73 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.4225 105.595 73.5575 105.73 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.7725 105.595 75.9075 105.73 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.1225 105.595 78.2575 105.73 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.4725 105.595 80.6075 105.73 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.8225 105.595 82.9575 105.73 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.1725 105.595 85.3075 105.73 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.5225 105.595 87.6575 105.73 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.8725 105.595 90.0075 105.73 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.2225 105.595 92.3575 105.73 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.5725 105.595 94.7075 105.73 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.9225 105.595 97.0575 105.73 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.2725 105.595 99.4075 105.73 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.6225 105.595 101.7575 105.73 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.9725 105.595 104.1075 105.73 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.3225 105.595 106.4575 105.73 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.6725 105.595 108.8075 105.73 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  26.865 20.67 27.005 92.64 ;
         LAYER metal4 ;
         RECT  129.035 98.1 129.175 108.12 ;
         LAYER metal3 ;
         RECT  125.4625 34.1275 125.5975 34.2625 ;
         LAYER metal3 ;
         RECT  69.5525 2.4725 69.6875 2.6075 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
         LAYER metal3 ;
         RECT  27.485 19.965 27.62 20.1 ;
         LAYER metal3 ;
         RECT  32.6375 96.185 112.2975 96.255 ;
         LAYER metal3 ;
         RECT  125.4625 25.1575 125.5975 25.2925 ;
         LAYER metal3 ;
         RECT  125.4625 22.1675 125.5975 22.3025 ;
         LAYER metal3 ;
         RECT  32.6375 8.415 109.4775 8.485 ;
         LAYER metal4 ;
         RECT  146.4175 78.34 146.5575 100.7425 ;
         LAYER metal3 ;
         RECT  125.4625 31.1375 125.5975 31.2725 ;
         LAYER metal4 ;
         RECT  131.755 5.85 131.895 20.81 ;
         LAYER metal4 ;
         RECT  15.21 44.59 15.35 59.55 ;
         LAYER metal4 ;
         RECT  32.57 17.5 32.71 95.49 ;
         LAYER metal3 ;
         RECT  119.29 93.14 119.425 93.275 ;
         LAYER metal3 ;
         RECT  31.4925 19.1775 31.6275 19.3125 ;
         LAYER metal3 ;
         RECT  103.8725 2.4725 104.0075 2.6075 ;
         LAYER metal3 ;
         RECT  25.575 11.9075 25.71 12.0425 ;
         LAYER metal3 ;
         RECT  58.1125 2.4725 58.2475 2.6075 ;
         LAYER metal4 ;
         RECT  119.905 20.67 120.045 92.64 ;
         LAYER metal3 ;
         RECT  21.3125 34.1275 21.4475 34.2625 ;
         LAYER metal3 ;
         RECT  20.9325 2.4725 21.0675 2.6075 ;
         LAYER metal3 ;
         RECT  21.3125 22.1675 21.4475 22.3025 ;
         LAYER metal3 ;
         RECT  21.3125 25.1575 21.4475 25.2925 ;
         LAYER metal3 ;
         RECT  144.685 107.9825 144.82 108.1175 ;
         LAYER metal3 ;
         RECT  92.4325 2.4725 92.5675 2.6075 ;
         LAYER metal4 ;
         RECT  114.2 17.5 114.34 95.49 ;
         LAYER metal4 ;
         RECT  115.28 20.67 115.42 92.57 ;
         LAYER metal3 ;
         RECT  32.6375 16.805 111.1225 16.875 ;
         LAYER metal3 ;
         RECT  21.3125 31.1375 21.4475 31.2725 ;
         LAYER metal3 ;
         RECT  21.3125 43.0975 21.4475 43.2325 ;
         LAYER metal4 ;
         RECT  31.49 20.67 31.63 92.57 ;
         LAYER metal3 ;
         RECT  123.1775 106.7175 123.3125 106.8525 ;
         LAYER metal4 ;
         RECT  17.93 2.47 18.07 17.43 ;
         LAYER metal3 ;
         RECT  125.4625 43.0975 125.5975 43.2325 ;
         LAYER metal3 ;
         RECT  32.6375 103.0375 109.4775 103.1075 ;
         LAYER metal3 ;
         RECT  23.7925 2.4725 23.9275 2.6075 ;
         LAYER metal3 ;
         RECT  35.2325 2.4725 35.3675 2.6075 ;
         LAYER metal3 ;
         RECT  125.4625 40.1075 125.5975 40.2425 ;
         LAYER metal3 ;
         RECT  121.2 101.0175 121.335 101.1525 ;
         LAYER metal3 ;
         RECT  46.6725 2.4725 46.8075 2.6075 ;
         LAYER metal3 ;
         RECT  80.9925 2.4725 81.1275 2.6075 ;
         LAYER metal3 ;
         RECT  115.2825 93.9275 115.4175 94.0625 ;
         LAYER metal3 ;
         RECT  21.3125 40.1075 21.4475 40.2425 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal3 ;
         RECT  26.6525 0.0025 26.7875 0.1375 ;
         LAYER metal3 ;
         RECT  126.99 41.6025 127.125 41.7375 ;
         LAYER metal4 ;
         RECT  119.345 20.6375 119.485 92.6025 ;
         LAYER metal3 ;
         RECT  19.785 44.5925 19.92 44.7275 ;
         LAYER metal3 ;
         RECT  126.99 38.6125 127.125 38.7475 ;
         LAYER metal3 ;
         RECT  126.99 29.6425 127.125 29.7775 ;
         LAYER metal3 ;
         RECT  32.6375 10.465 109.4775 10.535 ;
         LAYER metal3 ;
         RECT  19.785 20.6725 19.92 20.8075 ;
         LAYER metal3 ;
         RECT  19.785 35.6225 19.92 35.7575 ;
         LAYER metal3 ;
         RECT  19.785 41.6025 19.92 41.7375 ;
         LAYER metal4 ;
         RECT  27.425 20.6375 27.565 92.6025 ;
         LAYER metal3 ;
         RECT  83.8525 0.0025 83.9875 0.1375 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal4 ;
         RECT  24.93 20.6375 25.07 92.64 ;
         LAYER metal3 ;
         RECT  144.685 110.4525 144.82 110.5875 ;
         LAYER metal4 ;
         RECT  140.86 95.63 141.0 110.59 ;
         LAYER metal3 ;
         RECT  95.2925 0.0025 95.4275 0.1375 ;
         LAYER metal3 ;
         RECT  120.3175 109.1875 120.4525 109.3225 ;
         LAYER metal3 ;
         RECT  60.9725 0.0025 61.1075 0.1375 ;
         LAYER metal3 ;
         RECT  72.4125 0.0025 72.5475 0.1375 ;
         LAYER metal4 ;
         RECT  144.355 78.3075 144.495 100.71 ;
         LAYER metal3 ;
         RECT  23.7925 0.0025 23.9275 0.1375 ;
         LAYER metal3 ;
         RECT  121.2 103.4875 121.335 103.6225 ;
         LAYER metal3 ;
         RECT  121.2 98.5475 121.335 98.6825 ;
         LAYER metal3 ;
         RECT  19.785 26.6525 19.92 26.7875 ;
         LAYER metal3 ;
         RECT  25.575 14.3775 25.71 14.5125 ;
         LAYER metal3 ;
         RECT  126.99 26.6525 127.125 26.7875 ;
         LAYER metal3 ;
         RECT  32.6375 98.805 111.155 98.875 ;
         LAYER metal4 ;
         RECT  18.07 44.525 18.21 59.615 ;
         LAYER metal3 ;
         RECT  19.785 29.6425 19.92 29.7775 ;
         LAYER metal3 ;
         RECT  19.785 23.6625 19.92 23.7975 ;
         LAYER metal3 ;
         RECT  32.6375 101.145 109.5125 101.215 ;
         LAYER metal3 ;
         RECT  126.99 35.6225 127.125 35.7575 ;
         LAYER metal3 ;
         RECT  126.99 20.6725 127.125 20.8075 ;
         LAYER metal3 ;
         RECT  126.99 44.5925 127.125 44.7275 ;
         LAYER metal3 ;
         RECT  32.6375 14.185 111.155 14.255 ;
         LAYER metal3 ;
         RECT  126.99 23.6625 127.125 23.7975 ;
         LAYER metal3 ;
         RECT  19.785 32.6325 19.92 32.7675 ;
         LAYER metal4 ;
         RECT  113.74 17.5 113.88 95.49 ;
         LAYER metal3 ;
         RECT  49.5325 0.0025 49.6675 0.1375 ;
         LAYER metal3 ;
         RECT  19.785 38.6125 19.92 38.7475 ;
         LAYER metal3 ;
         RECT  38.0925 0.0025 38.2275 0.1375 ;
         LAYER metal3 ;
         RECT  106.7325 0.0025 106.8675 0.1375 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal3 ;
         RECT  126.99 32.6325 127.125 32.7675 ;
         LAYER metal3 ;
         RECT  25.575 9.4375 25.71 9.5725 ;
         LAYER metal4 ;
         RECT  128.895 5.785 129.035 20.875 ;
         LAYER metal4 ;
         RECT  33.03 17.5 33.17 95.49 ;
         LAYER metal4 ;
         RECT  121.84 20.6375 121.98 92.64 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 147.105 110.45 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 147.105 110.45 ;
   LAYER  metal3 ;
      RECT  24.35 0.9675 26.795 1.3825 ;
      RECT  27.21 0.9675 29.655 1.3825 ;
      RECT  30.07 0.9675 32.515 1.3825 ;
      RECT  32.93 0.9675 35.375 1.3825 ;
      RECT  35.79 0.9675 38.235 1.3825 ;
      RECT  38.65 0.9675 41.095 1.3825 ;
      RECT  41.51 0.9675 43.955 1.3825 ;
      RECT  44.37 0.9675 46.815 1.3825 ;
      RECT  47.23 0.9675 49.675 1.3825 ;
      RECT  50.09 0.9675 52.535 1.3825 ;
      RECT  52.95 0.9675 55.395 1.3825 ;
      RECT  55.81 0.9675 58.255 1.3825 ;
      RECT  58.67 0.9675 61.115 1.3825 ;
      RECT  61.53 0.9675 63.975 1.3825 ;
      RECT  64.39 0.9675 66.835 1.3825 ;
      RECT  67.25 0.9675 69.695 1.3825 ;
      RECT  70.11 0.9675 72.555 1.3825 ;
      RECT  72.97 0.9675 75.415 1.3825 ;
      RECT  75.83 0.9675 78.275 1.3825 ;
      RECT  78.69 0.9675 81.135 1.3825 ;
      RECT  81.55 0.9675 83.995 1.3825 ;
      RECT  84.41 0.9675 86.855 1.3825 ;
      RECT  87.27 0.9675 89.715 1.3825 ;
      RECT  90.13 0.9675 92.575 1.3825 ;
      RECT  92.99 0.9675 95.435 1.3825 ;
      RECT  95.85 0.9675 98.295 1.3825 ;
      RECT  98.71 0.9675 101.155 1.3825 ;
      RECT  101.57 0.9675 104.015 1.3825 ;
      RECT  104.43 0.9675 106.875 1.3825 ;
      RECT  107.29 0.9675 109.735 1.3825 ;
      RECT  110.15 0.9675 112.595 1.3825 ;
      RECT  113.01 0.9675 147.105 1.3825 ;
      RECT  21.49 0.9675 23.935 1.3825 ;
      RECT  0.14 45.5575 15.355 45.9725 ;
      RECT  0.14 45.9725 15.355 110.45 ;
      RECT  15.355 1.3825 15.77 45.5575 ;
      RECT  15.77 45.5575 23.935 45.9725 ;
      RECT  15.77 45.9725 23.935 110.45 ;
      RECT  15.355 45.9725 15.77 48.2875 ;
      RECT  15.355 48.7025 15.77 50.4975 ;
      RECT  15.355 50.9125 15.77 53.2275 ;
      RECT  15.355 53.6425 15.77 55.4375 ;
      RECT  15.355 55.8525 15.77 58.1675 ;
      RECT  15.355 58.5825 15.77 110.45 ;
      RECT  24.35 107.9425 122.755 108.3575 ;
      RECT  122.755 108.3575 123.17 110.45 ;
      RECT  123.17 1.3825 131.335 19.4275 ;
      RECT  123.17 19.4275 131.335 19.8425 ;
      RECT  131.335 19.8425 131.75 107.9425 ;
      RECT  131.75 1.3825 147.105 19.4275 ;
      RECT  131.75 19.4275 147.105 19.8425 ;
      RECT  131.335 17.1125 131.75 19.4275 ;
      RECT  131.335 14.9025 131.75 16.6975 ;
      RECT  131.335 12.1725 131.75 14.4875 ;
      RECT  131.335 9.9625 131.75 11.7575 ;
      RECT  131.335 1.3825 131.75 6.8175 ;
      RECT  131.335 7.2325 131.75 9.5475 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  146.685 108.3575 147.1 109.2075 ;
      RECT  146.685 109.6225 147.1 110.45 ;
      RECT  147.1 108.3575 147.105 109.2075 ;
      RECT  147.1 109.2075 147.105 109.6225 ;
      RECT  147.1 109.6225 147.105 110.45 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 45.5575 ;
      RECT  6.5225 1.3825 15.355 1.4675 ;
      RECT  6.5225 1.4675 15.355 45.5575 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 21.075 1.0525 ;
      RECT  6.5225 1.0525 21.075 1.3825 ;
      RECT  123.17 108.3575 140.5825 109.1225 ;
      RECT  123.17 109.1225 140.5825 109.2075 ;
      RECT  140.5825 108.3575 140.9975 109.1225 ;
      RECT  140.9975 108.3575 146.685 109.1225 ;
      RECT  140.9975 109.1225 146.685 109.2075 ;
      RECT  123.17 109.2075 140.5825 109.5375 ;
      RECT  123.17 109.5375 140.5825 109.6225 ;
      RECT  140.5825 109.5375 140.9975 109.6225 ;
      RECT  140.9975 109.2075 146.685 109.5375 ;
      RECT  140.9975 109.5375 146.685 109.6225 ;
      RECT  24.35 105.455 35.6825 105.87 ;
      RECT  24.35 105.87 35.6825 107.9425 ;
      RECT  35.6825 105.87 36.0975 107.9425 ;
      RECT  36.0975 105.87 122.755 107.9425 ;
      RECT  36.0975 105.455 38.0325 105.87 ;
      RECT  38.4475 105.455 40.3825 105.87 ;
      RECT  40.7975 105.455 42.7325 105.87 ;
      RECT  43.1475 105.455 45.0825 105.87 ;
      RECT  45.4975 105.455 47.4325 105.87 ;
      RECT  47.8475 105.455 49.7825 105.87 ;
      RECT  50.1975 105.455 52.1325 105.87 ;
      RECT  52.5475 105.455 54.4825 105.87 ;
      RECT  54.8975 105.455 56.8325 105.87 ;
      RECT  57.2475 105.455 59.1825 105.87 ;
      RECT  59.5975 105.455 61.5325 105.87 ;
      RECT  61.9475 105.455 63.8825 105.87 ;
      RECT  64.2975 105.455 66.2325 105.87 ;
      RECT  66.6475 105.455 68.5825 105.87 ;
      RECT  68.9975 105.455 70.9325 105.87 ;
      RECT  71.3475 105.455 73.2825 105.87 ;
      RECT  73.6975 105.455 75.6325 105.87 ;
      RECT  76.0475 105.455 77.9825 105.87 ;
      RECT  78.3975 105.455 80.3325 105.87 ;
      RECT  80.7475 105.455 82.6825 105.87 ;
      RECT  83.0975 105.455 85.0325 105.87 ;
      RECT  85.4475 105.455 87.3825 105.87 ;
      RECT  87.7975 105.455 89.7325 105.87 ;
      RECT  90.1475 105.455 92.0825 105.87 ;
      RECT  92.4975 105.455 94.4325 105.87 ;
      RECT  94.8475 105.455 96.7825 105.87 ;
      RECT  97.1975 105.455 99.1325 105.87 ;
      RECT  99.5475 105.455 101.4825 105.87 ;
      RECT  101.8975 105.455 103.8325 105.87 ;
      RECT  104.2475 105.455 106.1825 105.87 ;
      RECT  106.5975 105.455 108.5325 105.87 ;
      RECT  108.9475 105.455 122.755 105.87 ;
      RECT  123.17 19.8425 125.3225 33.9875 ;
      RECT  123.17 33.9875 125.3225 34.4025 ;
      RECT  125.7375 33.9875 131.335 34.4025 ;
      RECT  36.0975 1.3825 69.4125 2.3325 ;
      RECT  69.4125 1.3825 69.8275 2.3325 ;
      RECT  69.8275 1.3825 122.755 2.3325 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 45.5575 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 45.5575 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 45.5575 ;
      RECT  24.35 19.825 27.345 20.24 ;
      RECT  24.35 20.24 27.345 105.455 ;
      RECT  27.345 1.3825 27.76 19.825 ;
      RECT  27.345 20.24 27.76 105.455 ;
      RECT  27.76 19.825 35.6825 20.24 ;
      RECT  112.4375 96.045 122.755 96.395 ;
      RECT  27.76 20.24 32.4975 96.045 ;
      RECT  27.76 96.045 32.4975 96.395 ;
      RECT  27.76 96.395 32.4975 105.455 ;
      RECT  32.4975 20.24 35.6825 96.045 ;
      RECT  125.3225 19.8425 125.7375 22.0275 ;
      RECT  125.3225 22.4425 125.7375 25.0175 ;
      RECT  27.76 1.3825 32.4975 8.275 ;
      RECT  27.76 8.275 32.4975 8.625 ;
      RECT  35.6825 1.3825 36.0975 8.275 ;
      RECT  36.0975 2.7475 69.4125 8.275 ;
      RECT  69.4125 2.7475 69.8275 8.275 ;
      RECT  69.8275 2.7475 109.6175 8.275 ;
      RECT  109.6175 2.7475 112.4375 8.275 ;
      RECT  109.6175 8.275 112.4375 8.625 ;
      RECT  125.3225 25.4325 125.7375 30.9975 ;
      RECT  125.3225 31.4125 125.7375 33.9875 ;
      RECT  112.4375 2.7475 119.15 93.0 ;
      RECT  112.4375 93.0 119.15 93.415 ;
      RECT  119.15 2.7475 119.565 93.0 ;
      RECT  119.15 93.415 119.565 96.045 ;
      RECT  119.565 2.7475 122.755 93.0 ;
      RECT  119.565 93.0 122.755 93.415 ;
      RECT  119.565 93.415 122.755 96.045 ;
      RECT  27.76 8.625 31.3525 19.0375 ;
      RECT  27.76 19.0375 31.3525 19.4525 ;
      RECT  27.76 19.4525 31.3525 19.825 ;
      RECT  31.3525 8.625 31.7675 19.0375 ;
      RECT  31.3525 19.4525 31.7675 19.825 ;
      RECT  31.7675 8.625 32.4975 19.0375 ;
      RECT  31.7675 19.0375 32.4975 19.4525 ;
      RECT  31.7675 19.4525 32.4975 19.825 ;
      RECT  104.1475 2.3325 122.755 2.7475 ;
      RECT  24.35 1.3825 25.435 11.7675 ;
      RECT  24.35 11.7675 25.435 12.1825 ;
      RECT  24.35 12.1825 25.435 19.825 ;
      RECT  25.85 1.3825 27.345 11.7675 ;
      RECT  25.85 11.7675 27.345 12.1825 ;
      RECT  25.85 12.1825 27.345 19.825 ;
      RECT  58.3875 2.3325 69.4125 2.7475 ;
      RECT  15.77 33.9875 21.1725 34.4025 ;
      RECT  21.5875 33.9875 23.935 34.4025 ;
      RECT  21.5875 34.4025 23.935 45.5575 ;
      RECT  15.77 1.3825 20.7925 2.3325 ;
      RECT  15.77 2.3325 20.7925 2.7475 ;
      RECT  20.7925 1.3825 21.1725 2.3325 ;
      RECT  20.7925 2.7475 21.1725 33.9875 ;
      RECT  21.1725 1.3825 21.2075 2.3325 ;
      RECT  21.2075 1.3825 21.5875 2.3325 ;
      RECT  21.2075 2.3325 21.5875 2.7475 ;
      RECT  21.1725 2.7475 21.2075 22.0275 ;
      RECT  21.2075 2.7475 21.5875 22.0275 ;
      RECT  21.1725 22.4425 21.2075 25.0175 ;
      RECT  21.2075 22.4425 21.5875 25.0175 ;
      RECT  123.17 107.9425 144.545 108.2575 ;
      RECT  123.17 108.2575 144.545 108.3575 ;
      RECT  144.545 108.2575 144.96 108.3575 ;
      RECT  144.96 107.9425 147.105 108.2575 ;
      RECT  144.96 108.2575 147.105 108.3575 ;
      RECT  131.75 19.8425 144.545 107.8425 ;
      RECT  131.75 107.8425 144.545 107.9425 ;
      RECT  144.545 19.8425 144.96 107.8425 ;
      RECT  144.96 19.8425 147.105 107.8425 ;
      RECT  144.96 107.8425 147.105 107.9425 ;
      RECT  92.7075 2.3325 103.7325 2.7475 ;
      RECT  32.4975 17.015 35.6825 19.825 ;
      RECT  35.6825 17.015 36.0975 96.045 ;
      RECT  36.0975 17.015 69.4125 96.045 ;
      RECT  69.4125 17.015 69.8275 96.045 ;
      RECT  69.8275 17.015 109.6175 96.045 ;
      RECT  109.6175 17.015 111.2625 96.045 ;
      RECT  111.2625 16.665 112.4375 17.015 ;
      RECT  111.2625 17.015 112.4375 96.045 ;
      RECT  21.1725 25.4325 21.2075 30.9975 ;
      RECT  21.1725 31.4125 21.2075 33.9875 ;
      RECT  21.2075 25.4325 21.5875 30.9975 ;
      RECT  21.2075 31.4125 21.5875 33.9875 ;
      RECT  21.1725 43.3725 21.5875 45.5575 ;
      RECT  122.755 1.3825 123.0375 106.5775 ;
      RECT  122.755 106.5775 123.0375 106.9925 ;
      RECT  122.755 106.9925 123.0375 107.9425 ;
      RECT  123.0375 1.3825 123.17 106.5775 ;
      RECT  123.0375 106.9925 123.17 107.9425 ;
      RECT  123.17 34.4025 123.4525 106.5775 ;
      RECT  123.17 106.9925 123.4525 107.9425 ;
      RECT  123.4525 34.4025 125.3225 106.5775 ;
      RECT  123.4525 106.5775 125.3225 106.9925 ;
      RECT  123.4525 106.9925 125.3225 107.9425 ;
      RECT  125.3225 43.3725 125.7375 107.9425 ;
      RECT  35.6825 103.2475 36.0975 105.455 ;
      RECT  36.0975 103.2475 69.4125 105.455 ;
      RECT  69.4125 103.2475 69.8275 105.455 ;
      RECT  69.8275 103.2475 109.6175 105.455 ;
      RECT  109.6175 102.8975 112.4375 103.2475 ;
      RECT  109.6175 103.2475 112.4375 105.455 ;
      RECT  32.4975 103.2475 35.6825 105.455 ;
      RECT  23.935 1.3825 24.0675 2.3325 ;
      RECT  23.935 2.7475 24.0675 110.45 ;
      RECT  24.0675 1.3825 24.35 2.3325 ;
      RECT  24.0675 2.3325 24.35 2.7475 ;
      RECT  24.0675 2.7475 24.35 110.45 ;
      RECT  21.5875 1.3825 23.6525 2.3325 ;
      RECT  21.5875 2.3325 23.6525 2.7475 ;
      RECT  21.5875 2.7475 23.6525 33.9875 ;
      RECT  23.6525 1.3825 23.935 2.3325 ;
      RECT  23.6525 2.7475 23.935 33.9875 ;
      RECT  32.4975 1.3825 35.0925 2.3325 ;
      RECT  32.4975 2.3325 35.0925 2.7475 ;
      RECT  32.4975 2.7475 35.0925 8.275 ;
      RECT  35.0925 1.3825 35.5075 2.3325 ;
      RECT  35.0925 2.7475 35.5075 8.275 ;
      RECT  35.5075 1.3825 35.6825 2.3325 ;
      RECT  35.5075 2.3325 35.6825 2.7475 ;
      RECT  35.5075 2.7475 35.6825 8.275 ;
      RECT  125.3225 34.4025 125.7375 39.9675 ;
      RECT  125.3225 40.3825 125.7375 42.9575 ;
      RECT  112.4375 96.395 121.06 100.8775 ;
      RECT  112.4375 100.8775 121.06 101.2925 ;
      RECT  112.4375 101.2925 121.06 105.455 ;
      RECT  121.475 96.395 122.755 100.8775 ;
      RECT  121.475 100.8775 122.755 101.2925 ;
      RECT  121.475 101.2925 122.755 105.455 ;
      RECT  36.0975 2.3325 46.5325 2.7475 ;
      RECT  46.9475 2.3325 57.9725 2.7475 ;
      RECT  69.8275 2.3325 80.8525 2.7475 ;
      RECT  81.2675 2.3325 92.2925 2.7475 ;
      RECT  112.4375 93.415 115.1425 93.7875 ;
      RECT  112.4375 93.7875 115.1425 94.2025 ;
      RECT  112.4375 94.2025 115.1425 96.045 ;
      RECT  115.1425 93.415 115.5575 93.7875 ;
      RECT  115.1425 94.2025 115.5575 96.045 ;
      RECT  115.5575 93.415 119.15 93.7875 ;
      RECT  115.5575 93.7875 119.15 94.2025 ;
      RECT  115.5575 94.2025 119.15 96.045 ;
      RECT  21.1725 34.4025 21.5875 39.9675 ;
      RECT  21.1725 40.3825 21.5875 42.9575 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  0.14 0.2775 2.285 0.9675 ;
      RECT  2.285 0.2775 2.7 0.9675 ;
      RECT  2.7 0.2775 23.935 0.9675 ;
      RECT  24.35 0.14 26.5125 0.2775 ;
      RECT  24.35 0.2775 26.5125 0.9675 ;
      RECT  26.5125 0.2775 26.9275 0.9675 ;
      RECT  26.9275 0.2775 147.105 0.9675 ;
      RECT  125.7375 34.4025 126.85 41.4625 ;
      RECT  125.7375 41.4625 126.85 41.8775 ;
      RECT  125.7375 41.8775 126.85 107.9425 ;
      RECT  127.265 34.4025 131.335 41.4625 ;
      RECT  127.265 41.4625 131.335 41.8775 ;
      RECT  127.265 41.8775 131.335 107.9425 ;
      RECT  15.77 34.4025 19.645 44.4525 ;
      RECT  15.77 44.4525 19.645 44.8675 ;
      RECT  15.77 44.8675 19.645 45.5575 ;
      RECT  19.645 44.8675 20.06 45.5575 ;
      RECT  20.06 34.4025 21.1725 44.4525 ;
      RECT  20.06 44.4525 21.1725 44.8675 ;
      RECT  20.06 44.8675 21.1725 45.5575 ;
      RECT  126.85 38.8875 127.265 41.4625 ;
      RECT  125.7375 19.8425 126.85 29.5025 ;
      RECT  125.7375 29.5025 126.85 29.9175 ;
      RECT  125.7375 29.9175 126.85 33.9875 ;
      RECT  127.265 19.8425 131.335 29.5025 ;
      RECT  127.265 29.5025 131.335 29.9175 ;
      RECT  127.265 29.9175 131.335 33.9875 ;
      RECT  32.4975 8.625 35.6825 10.325 ;
      RECT  35.6825 8.625 36.0975 10.325 ;
      RECT  36.0975 8.625 69.4125 10.325 ;
      RECT  69.4125 8.625 69.8275 10.325 ;
      RECT  69.8275 8.625 109.6175 10.325 ;
      RECT  15.77 2.7475 19.645 20.5325 ;
      RECT  15.77 20.5325 19.645 20.9475 ;
      RECT  15.77 20.9475 19.645 33.9875 ;
      RECT  19.645 2.7475 20.06 20.5325 ;
      RECT  20.06 2.7475 20.7925 20.5325 ;
      RECT  20.06 20.5325 20.7925 20.9475 ;
      RECT  20.06 20.9475 20.7925 33.9875 ;
      RECT  19.645 34.4025 20.06 35.4825 ;
      RECT  19.645 41.8775 20.06 44.4525 ;
      RECT  123.17 109.6225 144.545 110.3125 ;
      RECT  123.17 110.3125 144.545 110.45 ;
      RECT  144.545 109.6225 144.96 110.3125 ;
      RECT  144.96 109.6225 146.685 110.3125 ;
      RECT  144.96 110.3125 146.685 110.45 ;
      RECT  84.1275 0.14 95.1525 0.2775 ;
      RECT  24.35 108.3575 120.1775 109.0475 ;
      RECT  24.35 109.0475 120.1775 109.4625 ;
      RECT  24.35 109.4625 120.1775 110.45 ;
      RECT  120.1775 108.3575 120.5925 109.0475 ;
      RECT  120.1775 109.4625 120.5925 110.45 ;
      RECT  120.5925 108.3575 122.755 109.0475 ;
      RECT  120.5925 109.0475 122.755 109.4625 ;
      RECT  120.5925 109.4625 122.755 110.45 ;
      RECT  61.2475 0.14 72.2725 0.2775 ;
      RECT  72.6875 0.14 83.7125 0.2775 ;
      RECT  23.935 0.2775 24.0675 0.9675 ;
      RECT  24.0675 0.14 24.35 0.2775 ;
      RECT  24.0675 0.2775 24.35 0.9675 ;
      RECT  2.7 0.14 23.6525 0.2775 ;
      RECT  121.06 101.2925 121.475 103.3475 ;
      RECT  121.06 103.7625 121.475 105.455 ;
      RECT  121.06 96.395 121.475 98.4075 ;
      RECT  121.06 98.8225 121.475 100.8775 ;
      RECT  25.435 12.1825 25.85 14.2375 ;
      RECT  25.435 14.6525 25.85 19.825 ;
      RECT  126.85 26.9275 127.265 29.5025 ;
      RECT  35.6825 96.395 36.0975 98.665 ;
      RECT  36.0975 96.395 69.4125 98.665 ;
      RECT  69.4125 96.395 69.8275 98.665 ;
      RECT  69.8275 96.395 109.6175 98.665 ;
      RECT  109.6175 96.395 111.295 98.665 ;
      RECT  111.295 96.395 112.4375 98.665 ;
      RECT  111.295 98.665 112.4375 99.015 ;
      RECT  111.295 99.015 112.4375 102.8975 ;
      RECT  32.4975 96.395 35.6825 98.665 ;
      RECT  19.645 26.9275 20.06 29.5025 ;
      RECT  19.645 20.9475 20.06 23.5225 ;
      RECT  19.645 23.9375 20.06 26.5125 ;
      RECT  35.6825 99.015 36.0975 101.005 ;
      RECT  35.6825 101.355 36.0975 102.8975 ;
      RECT  36.0975 99.015 69.4125 101.005 ;
      RECT  36.0975 101.355 69.4125 102.8975 ;
      RECT  69.4125 99.015 69.8275 101.005 ;
      RECT  69.4125 101.355 69.8275 102.8975 ;
      RECT  69.8275 99.015 109.6175 101.005 ;
      RECT  69.8275 101.355 109.6175 102.8975 ;
      RECT  109.6175 99.015 109.6525 101.005 ;
      RECT  109.6175 101.355 109.6525 102.8975 ;
      RECT  109.6525 99.015 111.295 101.005 ;
      RECT  109.6525 101.005 111.295 101.355 ;
      RECT  109.6525 101.355 111.295 102.8975 ;
      RECT  32.4975 99.015 35.6825 101.005 ;
      RECT  32.4975 101.355 35.6825 102.8975 ;
      RECT  126.85 34.4025 127.265 35.4825 ;
      RECT  126.85 35.8975 127.265 38.4725 ;
      RECT  126.85 19.8425 127.265 20.5325 ;
      RECT  126.85 41.8775 127.265 44.4525 ;
      RECT  126.85 44.8675 127.265 107.9425 ;
      RECT  109.6175 8.625 111.2625 14.045 ;
      RECT  109.6175 14.395 111.2625 16.665 ;
      RECT  111.2625 8.625 111.295 14.045 ;
      RECT  111.2625 14.395 111.295 16.665 ;
      RECT  111.295 8.625 112.4375 14.045 ;
      RECT  111.295 14.045 112.4375 14.395 ;
      RECT  111.295 14.395 112.4375 16.665 ;
      RECT  32.4975 10.675 35.6825 14.045 ;
      RECT  32.4975 14.395 35.6825 16.665 ;
      RECT  35.6825 10.675 36.0975 14.045 ;
      RECT  35.6825 14.395 36.0975 16.665 ;
      RECT  36.0975 10.675 69.4125 14.045 ;
      RECT  36.0975 14.395 69.4125 16.665 ;
      RECT  69.4125 10.675 69.8275 14.045 ;
      RECT  69.4125 14.395 69.8275 16.665 ;
      RECT  69.8275 10.675 109.6175 14.045 ;
      RECT  69.8275 14.395 109.6175 16.665 ;
      RECT  126.85 20.9475 127.265 23.5225 ;
      RECT  126.85 23.9375 127.265 26.5125 ;
      RECT  19.645 29.9175 20.06 32.4925 ;
      RECT  19.645 32.9075 20.06 33.9875 ;
      RECT  49.8075 0.14 60.8325 0.2775 ;
      RECT  19.645 35.8975 20.06 38.4725 ;
      RECT  19.645 38.8875 20.06 41.4625 ;
      RECT  26.9275 0.14 37.9525 0.2775 ;
      RECT  38.3675 0.14 49.3925 0.2775 ;
      RECT  95.5675 0.14 106.5925 0.2775 ;
      RECT  107.0075 0.14 147.105 0.2775 ;
      RECT  126.85 29.9175 127.265 32.4925 ;
      RECT  126.85 32.9075 127.265 33.9875 ;
      RECT  25.435 1.3825 25.85 9.2975 ;
      RECT  25.435 9.7125 25.85 11.7675 ;
   LAYER  metal4 ;
      RECT  0.14 92.92 26.585 110.45 ;
      RECT  26.585 92.92 27.285 110.45 ;
      RECT  27.285 97.82 128.755 108.4 ;
      RECT  27.285 108.4 128.755 110.45 ;
      RECT  128.755 92.92 129.455 97.82 ;
      RECT  128.755 108.4 129.455 110.45 ;
      RECT  0.14 0.14 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 20.39 ;
      RECT  0.4075 0.14 1.1075 9.5675 ;
      RECT  0.14 20.39 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 92.92 ;
      RECT  0.4075 32.53 1.1075 92.92 ;
      RECT  146.1375 20.39 146.8375 78.06 ;
      RECT  146.8375 20.39 147.105 78.06 ;
      RECT  146.8375 78.06 147.105 92.92 ;
      RECT  146.8375 92.92 147.105 97.82 ;
      RECT  146.1375 101.0225 146.8375 108.4 ;
      RECT  146.8375 97.82 147.105 101.0225 ;
      RECT  146.8375 101.0225 147.105 108.4 ;
      RECT  131.475 0.14 132.175 5.57 ;
      RECT  132.175 0.14 147.105 5.57 ;
      RECT  132.175 5.57 147.105 20.39 ;
      RECT  131.475 21.09 132.175 78.06 ;
      RECT  132.175 20.39 146.1375 21.09 ;
      RECT  1.1075 44.31 14.93 59.83 ;
      RECT  1.1075 59.83 14.93 92.92 ;
      RECT  14.93 32.53 15.63 44.31 ;
      RECT  14.93 59.83 15.63 92.92 ;
      RECT  27.285 92.92 32.29 95.77 ;
      RECT  27.285 95.77 32.29 97.82 ;
      RECT  32.29 95.77 32.99 97.82 ;
      RECT  32.99 95.77 128.755 97.82 ;
      RECT  27.285 5.57 32.29 17.22 ;
      RECT  32.29 5.57 32.99 17.22 ;
      RECT  114.62 92.92 128.755 95.77 ;
      RECT  114.62 78.06 115.0 92.85 ;
      RECT  114.62 92.85 115.0 92.92 ;
      RECT  115.0 92.85 115.7 92.92 ;
      RECT  114.62 20.39 115.0 21.09 ;
      RECT  114.62 21.09 115.0 78.06 ;
      RECT  31.21 92.85 31.91 92.92 ;
      RECT  31.91 78.06 32.29 92.85 ;
      RECT  31.91 92.85 32.29 92.92 ;
      RECT  31.91 20.39 32.29 21.09 ;
      RECT  31.91 21.09 32.29 78.06 ;
      RECT  17.65 0.14 18.35 2.19 ;
      RECT  18.35 0.14 26.585 2.19 ;
      RECT  18.35 2.19 26.585 9.5675 ;
      RECT  17.65 17.71 18.35 20.39 ;
      RECT  18.35 9.5675 26.585 17.71 ;
      RECT  114.62 17.22 119.065 20.3575 ;
      RECT  114.62 20.3575 119.065 20.39 ;
      RECT  119.065 17.22 119.765 20.3575 ;
      RECT  115.7 78.06 119.065 92.85 ;
      RECT  115.7 92.85 119.065 92.8825 ;
      RECT  115.7 92.8825 119.065 92.92 ;
      RECT  119.065 92.8825 119.625 92.92 ;
      RECT  115.7 20.39 119.065 21.09 ;
      RECT  115.7 21.09 119.065 78.06 ;
      RECT  26.585 0.14 27.145 20.3575 ;
      RECT  26.585 20.3575 27.145 20.39 ;
      RECT  27.145 0.14 27.285 20.3575 ;
      RECT  27.285 17.22 27.845 20.3575 ;
      RECT  27.845 17.22 32.29 20.3575 ;
      RECT  27.845 20.3575 32.29 20.39 ;
      RECT  27.845 78.06 31.21 92.85 ;
      RECT  27.285 92.8825 27.845 92.92 ;
      RECT  27.845 92.85 31.21 92.8825 ;
      RECT  27.845 92.8825 31.21 92.92 ;
      RECT  27.845 20.39 31.21 21.09 ;
      RECT  27.845 21.09 31.21 78.06 ;
      RECT  1.1075 20.39 2.47 32.53 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 44.31 ;
      RECT  2.47 32.5625 3.17 44.31 ;
      RECT  3.17 32.53 14.93 32.5625 ;
      RECT  3.17 32.5625 14.93 44.31 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 17.71 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  1.1075 17.71 2.47 20.39 ;
      RECT  3.17 17.71 17.65 20.39 ;
      RECT  25.35 32.53 26.585 44.31 ;
      RECT  25.35 44.31 26.585 59.83 ;
      RECT  25.35 59.83 26.585 92.92 ;
      RECT  18.35 17.71 24.65 20.3575 ;
      RECT  18.35 20.3575 24.65 20.39 ;
      RECT  24.65 17.71 25.35 20.3575 ;
      RECT  25.35 17.71 26.585 20.3575 ;
      RECT  25.35 20.3575 26.585 20.39 ;
      RECT  3.17 20.39 24.65 32.53 ;
      RECT  25.35 20.39 26.585 32.53 ;
      RECT  129.455 108.4 140.58 110.45 ;
      RECT  141.28 108.4 147.105 110.45 ;
      RECT  129.455 92.92 140.58 95.35 ;
      RECT  129.455 95.35 140.58 97.82 ;
      RECT  140.58 92.92 141.28 95.35 ;
      RECT  129.455 97.82 140.58 101.0225 ;
      RECT  129.455 101.0225 140.58 108.4 ;
      RECT  141.28 101.0225 146.1375 108.4 ;
      RECT  132.175 21.09 144.075 78.0275 ;
      RECT  132.175 78.0275 144.075 78.06 ;
      RECT  144.075 21.09 144.775 78.0275 ;
      RECT  144.775 21.09 146.1375 78.0275 ;
      RECT  144.775 78.0275 146.1375 78.06 ;
      RECT  144.775 78.06 146.1375 92.92 ;
      RECT  141.28 92.92 144.075 95.35 ;
      RECT  144.775 92.92 146.1375 95.35 ;
      RECT  141.28 95.35 144.075 97.82 ;
      RECT  144.775 95.35 146.1375 97.82 ;
      RECT  141.28 97.82 144.075 100.99 ;
      RECT  141.28 100.99 144.075 101.0225 ;
      RECT  144.075 100.99 144.775 101.0225 ;
      RECT  144.775 97.82 146.1375 100.99 ;
      RECT  144.775 100.99 146.1375 101.0225 ;
      RECT  15.63 32.53 17.79 44.245 ;
      RECT  15.63 44.245 17.79 44.31 ;
      RECT  17.79 32.53 18.49 44.245 ;
      RECT  18.49 32.53 24.65 44.245 ;
      RECT  18.49 44.245 24.65 44.31 ;
      RECT  15.63 44.31 17.79 59.83 ;
      RECT  18.49 44.31 24.65 59.83 ;
      RECT  15.63 59.83 17.79 59.895 ;
      RECT  15.63 59.895 17.79 92.92 ;
      RECT  17.79 59.895 18.49 92.92 ;
      RECT  18.49 59.83 24.65 59.895 ;
      RECT  18.49 59.895 24.65 92.92 ;
      RECT  1.1075 0.14 5.825 2.19 ;
      RECT  6.525 0.14 17.65 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 17.65 9.5675 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  6.525 9.5675 17.65 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  3.17 15.24 5.825 17.71 ;
      RECT  5.825 15.24 6.525 17.71 ;
      RECT  6.525 9.6 17.65 15.24 ;
      RECT  6.525 15.24 17.65 17.71 ;
      RECT  27.285 0.14 128.615 5.505 ;
      RECT  27.285 5.505 128.615 5.57 ;
      RECT  128.615 0.14 129.315 5.505 ;
      RECT  129.315 0.14 131.475 5.505 ;
      RECT  129.315 5.505 131.475 5.57 ;
      RECT  32.99 5.57 128.615 17.22 ;
      RECT  129.315 5.57 131.475 17.22 ;
      RECT  129.315 20.39 131.475 21.09 ;
      RECT  128.615 21.155 129.315 78.06 ;
      RECT  129.315 21.09 131.475 21.155 ;
      RECT  129.315 21.155 131.475 78.06 ;
      RECT  119.765 17.22 128.615 20.3575 ;
      RECT  129.315 17.22 131.475 20.3575 ;
      RECT  129.315 20.3575 131.475 20.39 ;
      RECT  33.45 92.92 113.46 95.77 ;
      RECT  33.45 17.22 113.46 20.39 ;
      RECT  33.45 78.06 113.46 92.92 ;
      RECT  33.45 20.39 113.46 21.09 ;
      RECT  33.45 21.09 113.46 78.06 ;
      RECT  120.325 78.06 121.56 92.92 ;
      RECT  122.26 78.06 144.075 92.92 ;
      RECT  120.325 20.39 121.56 21.09 ;
      RECT  122.26 20.39 128.615 21.09 ;
      RECT  120.325 21.09 121.56 21.155 ;
      RECT  122.26 21.09 128.615 21.155 ;
      RECT  120.325 21.155 121.56 78.06 ;
      RECT  122.26 21.155 128.615 78.06 ;
      RECT  119.765 20.3575 121.56 20.39 ;
      RECT  122.26 20.3575 128.615 20.39 ;
   END
END    freepdk45_sram_1w1r_96x32_32
END    LIBRARY
