/home/yl996/proj/mcp-eda-example/libraries/FreePDK45/OpenRAM/macros/freepdk45_sram_1w1r_256x48_12/freepdk45_sram_1w1r_256x48_12.lef