../macros/freepdk45_sram_1rw0r_128x44/freepdk45_sram_1rw0r_128x44.lef