../macros/freepdk45_sram_1w1r_32x32/freepdk45_sram_1w1r_32x32.lef