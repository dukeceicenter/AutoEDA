VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_256x4_1
   CLASS BLOCK ;
   SIZE 94.805 BY 107.625 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.91 1.105 35.045 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.77 1.105 37.905 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.63 1.105 40.765 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.49 1.105 43.625 1.24 ;
      END
   END din0[3]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14.89 1.105 15.025 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.75 1.105 17.885 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.61 1.105 20.745 1.24 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.17 52.41 9.305 52.545 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.17 55.14 9.305 55.275 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.17 57.35 9.305 57.485 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.17 60.08 9.305 60.215 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.17 62.29 9.305 62.425 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.78 106.385 76.915 106.52 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.92 106.385 74.055 106.52 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.06 106.385 71.195 106.52 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.36 29.27 85.495 29.405 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.36 26.54 85.495 26.675 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.36 24.33 85.495 24.465 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.36 21.6 85.495 21.735 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.36 19.39 85.495 19.525 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 10.81 0.42 10.945 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.385 95.13 94.52 95.265 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 10.895 6.3825 11.03 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.2825 95.045 88.4175 95.18 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.47 1.105 23.605 1.24 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.33 1.105 26.465 1.24 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.19 1.105 29.325 1.24 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.05 1.105 32.185 1.24 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.4025 92.1575 28.5375 92.2925 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.8025 92.1575 37.9375 92.2925 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.2025 92.1575 47.3375 92.2925 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.6025 92.1575 56.7375 92.2925 ;
      END
   END dout1[3]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  15.6125 31.87 15.7475 32.005 ;
         LAYER metal3 ;
         RECT  70.2625 79.71 70.3975 79.845 ;
         LAYER metal3 ;
         RECT  15.2675 43.83 15.4025 43.965 ;
         LAYER metal3 ;
         RECT  15.2675 46.82 15.4025 46.955 ;
         LAYER metal4 ;
         RECT  0.6875 19.55 0.8275 41.9525 ;
         LAYER metal4 ;
         RECT  82.92 83.8825 83.06 93.9025 ;
         LAYER metal3 ;
         RECT  65.9675 16.37 66.1025 16.505 ;
         LAYER metal3 ;
         RECT  79.0675 43.83 79.2025 43.965 ;
         LAYER metal3 ;
         RECT  92.245 93.765 92.38 93.9 ;
         LAYER metal3 ;
         RECT  25.0825 16.37 25.2175 16.505 ;
         LAYER metal3 ;
         RECT  79.0675 49.81 79.2025 49.945 ;
         LAYER metal4 ;
         RECT  85.64 17.9575 85.78 30.5125 ;
         LAYER metal3 ;
         RECT  78.7225 31.87 78.8575 32.005 ;
         LAYER metal3 ;
         RECT  23.1875 2.47 23.3225 2.605 ;
         LAYER metal4 ;
         RECT  70.26 30.3725 70.4 78.3525 ;
         LAYER metal3 ;
         RECT  79.0675 46.82 79.2025 46.955 ;
         LAYER metal3 ;
         RECT  79.0675 40.84 79.2025 40.975 ;
         LAYER metal3 ;
         RECT  72.895 78.9225 73.03 79.0575 ;
         LAYER metal3 ;
         RECT  25.2175 17.3375 57.4075 17.4075 ;
         LAYER metal3 ;
         RECT  14.6075 2.47 14.7425 2.605 ;
         LAYER metal3 ;
         RECT  15.6125 34.86 15.7475 34.995 ;
         LAYER metal3 ;
         RECT  25.2175 89.6 57.4075 89.67 ;
         LAYER metal3 ;
         RECT  15.2675 40.84 15.4025 40.975 ;
         LAYER metal4 ;
         RECT  69.18 27.2025 69.32 81.2725 ;
         LAYER metal4 ;
         RECT  20.82 30.3725 20.96 78.4225 ;
         LAYER metal3 ;
         RECT  77.0625 105.02 77.1975 105.155 ;
         LAYER metal4 ;
         RECT  18.2 4.285 18.34 24.185 ;
         LAYER metal3 ;
         RECT  21.44 29.6675 21.575 29.8025 ;
         LAYER metal3 ;
         RECT  25.2175 81.9675 67.2775 82.0375 ;
         LAYER metal4 ;
         RECT  93.9775 64.1225 94.1175 86.525 ;
         LAYER metal4 ;
         RECT  24.07 30.3725 24.21 78.3525 ;
         LAYER metal4 ;
         RECT  76.13 84.36 76.27 104.26 ;
         LAYER metal3 ;
         RECT  2.425 12.175 2.56 12.31 ;
         LAYER metal3 ;
         RECT  78.7225 34.86 78.8575 34.995 ;
         LAYER metal4 ;
         RECT  73.51 30.3725 73.65 78.4225 ;
         LAYER metal4 ;
         RECT  11.605 12.1725 11.745 27.1325 ;
         LAYER metal3 ;
         RECT  24.0725 28.88 24.2075 29.015 ;
         LAYER metal3 ;
         RECT  34.6275 2.47 34.7625 2.605 ;
         LAYER metal4 ;
         RECT  25.15 27.2025 25.29 81.2725 ;
         LAYER metal3 ;
         RECT  25.2175 26.5075 66.1025 26.5775 ;
         LAYER metal3 ;
         RECT  15.2675 49.81 15.4025 49.945 ;
         LAYER metal4 ;
         RECT  8.885 51.3025 9.025 63.8575 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  82.78 18.0225 82.92 30.5775 ;
         LAYER metal3 ;
         RECT  65.9675 14.55 66.1025 14.685 ;
         LAYER metal4 ;
         RECT  19.23 30.34 19.37 78.4225 ;
         LAYER metal4 ;
         RECT  6.105 9.7025 6.245 24.6625 ;
         LAYER metal3 ;
         RECT  80.875 42.335 81.01 42.47 ;
         LAYER metal3 ;
         RECT  13.46 45.325 13.595 45.46 ;
         LAYER metal3 ;
         RECT  25.0825 14.55 25.2175 14.685 ;
         LAYER metal3 ;
         RECT  14.085 36.355 14.22 36.49 ;
         LAYER metal3 ;
         RECT  25.2175 87.7075 57.4425 87.7775 ;
         LAYER metal3 ;
         RECT  25.2175 84.5875 66.135 84.6575 ;
         LAYER metal3 ;
         RECT  74.2025 107.49 74.3375 107.625 ;
         LAYER metal3 ;
         RECT  25.2175 19.3875 57.4075 19.4575 ;
         LAYER metal4 ;
         RECT  72.95 30.34 73.09 78.385 ;
         LAYER metal3 ;
         RECT  80.875 48.315 81.01 48.45 ;
         LAYER metal3 ;
         RECT  13.46 39.345 13.595 39.48 ;
         LAYER metal3 ;
         RECT  80.875 51.305 81.01 51.44 ;
         LAYER metal3 ;
         RECT  80.25 33.365 80.385 33.5 ;
         LAYER metal4 ;
         RECT  78.0725 84.2925 78.2125 104.3275 ;
         LAYER metal3 ;
         RECT  13.46 42.335 13.595 42.47 ;
         LAYER metal4 ;
         RECT  25.61 27.2025 25.75 81.2725 ;
         LAYER metal3 ;
         RECT  80.875 45.325 81.01 45.46 ;
         LAYER metal4 ;
         RECT  11.745 51.2375 11.885 63.7925 ;
         LAYER metal3 ;
         RECT  25.2175 23.8875 66.135 23.9575 ;
         LAYER metal3 ;
         RECT  17.4675 0.0 17.6025 0.135 ;
         LAYER metal3 ;
         RECT  14.085 30.375 14.22 30.51 ;
         LAYER metal3 ;
         RECT  26.0475 0.0 26.1825 0.135 ;
         LAYER metal3 ;
         RECT  14.085 33.365 14.22 33.5 ;
         LAYER metal3 ;
         RECT  13.46 48.315 13.595 48.45 ;
         LAYER metal4 ;
         RECT  75.1 30.34 75.24 78.4225 ;
         LAYER metal3 ;
         RECT  80.25 36.355 80.385 36.49 ;
         LAYER metal4 ;
         RECT  91.915 64.09 92.055 86.4925 ;
         LAYER metal3 ;
         RECT  13.46 51.305 13.595 51.44 ;
         LAYER metal3 ;
         RECT  92.245 96.235 92.38 96.37 ;
         LAYER metal3 ;
         RECT  80.25 30.375 80.385 30.51 ;
         LAYER metal4 ;
         RECT  68.72 27.2025 68.86 81.2725 ;
         LAYER metal4 ;
         RECT  2.75 19.5825 2.89 41.985 ;
         LAYER metal4 ;
         RECT  21.38 30.34 21.52 78.385 ;
         LAYER metal4 ;
         RECT  88.42 81.4125 88.56 96.3725 ;
         LAYER metal3 ;
         RECT  2.425 9.705 2.56 9.84 ;
         LAYER metal3 ;
         RECT  37.4875 0.0 37.6225 0.135 ;
         LAYER metal3 ;
         RECT  80.875 39.345 81.01 39.48 ;
         LAYER metal4 ;
         RECT  16.2575 4.2175 16.3975 24.2525 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 94.665 107.485 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 94.665 107.485 ;
   LAYER  metal3 ;
      RECT  34.77 0.14 35.185 0.965 ;
      RECT  35.185 0.965 37.63 1.38 ;
      RECT  38.045 0.965 40.49 1.38 ;
      RECT  40.905 0.965 43.35 1.38 ;
      RECT  43.765 0.965 94.665 1.38 ;
      RECT  0.14 0.965 14.75 1.38 ;
      RECT  15.165 0.965 17.61 1.38 ;
      RECT  18.025 0.965 20.47 1.38 ;
      RECT  0.14 52.27 9.03 52.685 ;
      RECT  0.14 52.685 9.03 107.485 ;
      RECT  9.03 1.38 9.445 52.27 ;
      RECT  9.445 52.27 34.77 52.685 ;
      RECT  9.03 52.685 9.445 55.0 ;
      RECT  9.03 55.415 9.445 57.21 ;
      RECT  9.03 57.625 9.445 59.94 ;
      RECT  9.03 60.355 9.445 62.15 ;
      RECT  9.03 62.565 9.445 107.485 ;
      RECT  76.64 106.66 77.055 107.485 ;
      RECT  77.055 106.245 94.665 106.66 ;
      RECT  77.055 106.66 94.665 107.485 ;
      RECT  74.195 106.245 76.64 106.66 ;
      RECT  35.185 106.245 70.92 106.66 ;
      RECT  71.335 106.245 73.78 106.66 ;
      RECT  77.055 1.38 85.22 29.13 ;
      RECT  77.055 29.13 85.22 29.545 ;
      RECT  85.22 29.545 85.635 106.245 ;
      RECT  85.635 1.38 94.665 29.13 ;
      RECT  85.635 29.13 94.665 29.545 ;
      RECT  85.22 26.815 85.635 29.13 ;
      RECT  85.22 24.605 85.635 26.4 ;
      RECT  85.22 21.875 85.635 24.19 ;
      RECT  85.22 1.38 85.635 19.25 ;
      RECT  85.22 19.665 85.635 21.46 ;
      RECT  0.14 1.38 0.145 10.67 ;
      RECT  0.14 10.67 0.145 11.085 ;
      RECT  0.14 11.085 0.145 52.27 ;
      RECT  0.145 1.38 0.56 10.67 ;
      RECT  0.145 11.085 0.56 52.27 ;
      RECT  94.245 29.545 94.66 94.99 ;
      RECT  94.245 95.405 94.66 106.245 ;
      RECT  94.66 29.545 94.665 94.99 ;
      RECT  94.66 94.99 94.665 95.405 ;
      RECT  94.66 95.405 94.665 106.245 ;
      RECT  0.56 10.67 6.1075 10.755 ;
      RECT  0.56 10.755 6.1075 11.085 ;
      RECT  6.1075 10.67 6.5225 10.755 ;
      RECT  6.5225 10.67 9.03 10.755 ;
      RECT  6.5225 10.755 9.03 11.085 ;
      RECT  0.56 11.085 6.1075 11.17 ;
      RECT  6.1075 11.17 6.5225 52.27 ;
      RECT  6.5225 11.085 9.03 11.17 ;
      RECT  6.5225 11.17 9.03 52.27 ;
      RECT  85.635 29.545 88.1425 94.905 ;
      RECT  85.635 94.905 88.1425 94.99 ;
      RECT  88.1425 29.545 88.5575 94.905 ;
      RECT  88.5575 94.905 94.245 94.99 ;
      RECT  85.635 94.99 88.1425 95.32 ;
      RECT  85.635 95.32 88.1425 95.405 ;
      RECT  88.1425 95.32 88.5575 95.405 ;
      RECT  88.5575 94.99 94.245 95.32 ;
      RECT  88.5575 95.32 94.245 95.405 ;
      RECT  20.885 0.965 23.33 1.38 ;
      RECT  23.745 0.965 26.19 1.38 ;
      RECT  26.605 0.965 29.05 1.38 ;
      RECT  29.465 0.965 31.91 1.38 ;
      RECT  32.325 0.965 34.77 1.38 ;
      RECT  9.445 92.0175 28.2625 92.4325 ;
      RECT  9.445 92.4325 28.2625 107.485 ;
      RECT  28.2625 92.4325 28.6775 107.485 ;
      RECT  28.6775 92.0175 34.77 92.4325 ;
      RECT  28.6775 92.4325 34.77 107.485 ;
      RECT  35.185 92.0175 37.6625 92.4325 ;
      RECT  35.185 92.4325 37.6625 106.245 ;
      RECT  37.6625 92.4325 38.0775 106.245 ;
      RECT  38.0775 92.4325 76.64 106.245 ;
      RECT  38.0775 92.0175 47.0625 92.4325 ;
      RECT  47.4775 92.0175 56.4625 92.4325 ;
      RECT  56.8775 92.0175 76.64 92.4325 ;
      RECT  9.445 31.73 15.4725 32.145 ;
      RECT  15.4725 1.38 15.8875 31.73 ;
      RECT  15.8875 31.73 34.77 32.145 ;
      RECT  15.8875 32.145 34.77 52.27 ;
      RECT  38.0775 79.57 70.1225 79.985 ;
      RECT  70.1225 1.38 70.5375 79.57 ;
      RECT  70.1225 79.985 70.5375 92.0175 ;
      RECT  70.5375 79.57 76.64 79.985 ;
      RECT  70.5375 79.985 76.64 92.0175 ;
      RECT  9.445 43.69 15.1275 44.105 ;
      RECT  15.5425 43.69 15.8875 44.105 ;
      RECT  15.5425 44.105 15.8875 52.27 ;
      RECT  15.1275 44.105 15.4725 46.68 ;
      RECT  15.4725 44.105 15.5425 46.68 ;
      RECT  38.0775 1.38 65.8275 16.23 ;
      RECT  38.0775 16.23 65.8275 16.645 ;
      RECT  66.2425 1.38 70.1225 16.23 ;
      RECT  66.2425 16.23 70.1225 16.645 ;
      RECT  77.055 43.69 78.9275 44.105 ;
      RECT  79.3425 43.69 85.22 44.105 ;
      RECT  88.5575 29.545 92.105 93.625 ;
      RECT  88.5575 93.625 92.105 94.04 ;
      RECT  88.5575 94.04 92.105 94.905 ;
      RECT  92.105 29.545 92.52 93.625 ;
      RECT  92.105 94.04 92.52 94.905 ;
      RECT  92.52 29.545 94.245 93.625 ;
      RECT  92.52 93.625 94.245 94.04 ;
      RECT  92.52 94.04 94.245 94.905 ;
      RECT  15.8875 16.23 24.9425 16.645 ;
      RECT  25.3575 16.23 34.77 16.645 ;
      RECT  78.9275 50.085 79.3425 106.245 ;
      RECT  77.055 29.545 78.5825 31.73 ;
      RECT  77.055 31.73 78.5825 32.145 ;
      RECT  77.055 32.145 78.5825 43.69 ;
      RECT  78.5825 29.545 78.9275 31.73 ;
      RECT  78.9275 29.545 78.9975 31.73 ;
      RECT  78.9975 29.545 79.3425 31.73 ;
      RECT  78.9975 31.73 79.3425 32.145 ;
      RECT  15.8875 1.38 23.0475 2.33 ;
      RECT  15.8875 2.33 23.0475 2.745 ;
      RECT  15.8875 2.745 23.0475 16.23 ;
      RECT  23.0475 1.38 23.4625 2.33 ;
      RECT  23.0475 2.745 23.4625 16.23 ;
      RECT  23.4625 1.38 24.9425 2.33 ;
      RECT  23.4625 2.33 24.9425 2.745 ;
      RECT  23.4625 2.745 24.9425 16.23 ;
      RECT  78.9275 44.105 79.3425 46.68 ;
      RECT  78.9275 47.095 79.3425 49.67 ;
      RECT  78.9275 41.115 78.9975 43.69 ;
      RECT  78.9975 32.145 79.3425 40.7 ;
      RECT  78.9975 41.115 79.3425 43.69 ;
      RECT  70.5375 1.38 72.755 78.7825 ;
      RECT  70.5375 78.7825 72.755 79.1975 ;
      RECT  70.5375 79.1975 72.755 79.57 ;
      RECT  72.755 1.38 73.17 78.7825 ;
      RECT  72.755 79.1975 73.17 79.57 ;
      RECT  73.17 1.38 76.64 78.7825 ;
      RECT  73.17 78.7825 76.64 79.1975 ;
      RECT  73.17 79.1975 76.64 79.57 ;
      RECT  35.185 1.38 37.6625 17.1975 ;
      RECT  37.6625 1.38 38.0775 17.1975 ;
      RECT  38.0775 16.645 57.5475 17.1975 ;
      RECT  57.5475 16.645 65.8275 17.1975 ;
      RECT  57.5475 17.1975 65.8275 17.5475 ;
      RECT  24.9425 16.645 25.0775 17.1975 ;
      RECT  24.9425 17.1975 25.0775 17.5475 ;
      RECT  24.9425 17.5475 25.0775 31.73 ;
      RECT  25.0775 16.645 25.3575 17.1975 ;
      RECT  25.3575 16.645 34.77 17.1975 ;
      RECT  9.445 1.38 14.4675 2.33 ;
      RECT  9.445 2.33 14.4675 2.745 ;
      RECT  14.4675 1.38 14.8825 2.33 ;
      RECT  14.4675 2.745 14.8825 31.73 ;
      RECT  14.8825 1.38 15.4725 2.33 ;
      RECT  14.8825 2.33 15.4725 2.745 ;
      RECT  14.8825 2.745 15.4725 31.73 ;
      RECT  15.4725 32.145 15.5425 34.72 ;
      RECT  15.5425 32.145 15.8875 34.72 ;
      RECT  15.5425 35.135 15.8875 43.69 ;
      RECT  9.445 52.685 25.0775 89.46 ;
      RECT  9.445 89.46 25.0775 89.81 ;
      RECT  9.445 89.81 25.0775 92.0175 ;
      RECT  25.0775 89.81 28.2625 92.0175 ;
      RECT  28.2625 89.81 28.6775 92.0175 ;
      RECT  28.6775 89.81 34.77 92.0175 ;
      RECT  38.0775 89.81 57.5475 92.0175 ;
      RECT  57.5475 89.46 70.1225 89.81 ;
      RECT  57.5475 89.81 70.1225 92.0175 ;
      RECT  34.77 89.81 35.185 107.485 ;
      RECT  35.185 89.81 37.6625 92.0175 ;
      RECT  37.6625 89.81 38.0775 92.0175 ;
      RECT  15.1275 32.145 15.4725 40.7 ;
      RECT  15.1275 41.115 15.4725 43.69 ;
      RECT  15.4725 35.135 15.5425 40.7 ;
      RECT  15.4725 41.115 15.5425 43.69 ;
      RECT  76.64 1.38 76.9225 104.88 ;
      RECT  76.64 104.88 76.9225 105.295 ;
      RECT  76.64 105.295 76.9225 106.245 ;
      RECT  76.9225 1.38 77.055 104.88 ;
      RECT  76.9225 105.295 77.055 106.245 ;
      RECT  77.055 44.105 77.3375 104.88 ;
      RECT  77.055 105.295 77.3375 106.245 ;
      RECT  77.3375 44.105 78.9275 104.88 ;
      RECT  77.3375 104.88 78.9275 105.295 ;
      RECT  77.3375 105.295 78.9275 106.245 ;
      RECT  15.8875 16.645 21.3 29.5275 ;
      RECT  15.8875 29.5275 21.3 29.9425 ;
      RECT  15.8875 29.9425 21.3 31.73 ;
      RECT  21.3 16.645 21.715 29.5275 ;
      RECT  21.3 29.9425 21.715 31.73 ;
      RECT  21.715 29.5275 24.9425 29.9425 ;
      RECT  21.715 29.9425 24.9425 31.73 ;
      RECT  25.0775 52.685 28.2625 81.8275 ;
      RECT  28.2625 52.685 28.6775 81.8275 ;
      RECT  28.6775 52.685 34.77 81.8275 ;
      RECT  38.0775 79.985 57.5475 81.8275 ;
      RECT  57.5475 79.985 67.4175 81.8275 ;
      RECT  67.4175 79.985 70.1225 81.8275 ;
      RECT  67.4175 81.8275 70.1225 82.1775 ;
      RECT  67.4175 82.1775 70.1225 89.46 ;
      RECT  0.56 11.17 2.285 12.035 ;
      RECT  0.56 12.035 2.285 12.45 ;
      RECT  0.56 12.45 2.285 52.27 ;
      RECT  2.285 11.17 2.7 12.035 ;
      RECT  2.285 12.45 2.7 52.27 ;
      RECT  2.7 11.17 6.1075 12.035 ;
      RECT  2.7 12.035 6.1075 12.45 ;
      RECT  2.7 12.45 6.1075 52.27 ;
      RECT  78.5825 32.145 78.9275 34.72 ;
      RECT  78.5825 35.135 78.9275 43.69 ;
      RECT  78.9275 32.145 78.9975 34.72 ;
      RECT  78.9275 35.135 78.9975 40.7 ;
      RECT  21.715 16.645 23.9325 28.74 ;
      RECT  21.715 28.74 23.9325 29.155 ;
      RECT  21.715 29.155 23.9325 29.5275 ;
      RECT  23.9325 16.645 24.3475 28.74 ;
      RECT  23.9325 29.155 24.3475 29.5275 ;
      RECT  24.3475 16.645 24.9425 28.74 ;
      RECT  24.3475 28.74 24.9425 29.155 ;
      RECT  24.3475 29.155 24.9425 29.5275 ;
      RECT  25.3575 1.38 34.4875 2.33 ;
      RECT  25.3575 2.33 34.4875 2.745 ;
      RECT  25.3575 2.745 34.4875 16.23 ;
      RECT  34.4875 1.38 34.77 2.33 ;
      RECT  34.4875 2.745 34.77 16.23 ;
      RECT  34.77 1.38 34.9025 2.33 ;
      RECT  34.77 2.745 34.9025 17.1975 ;
      RECT  34.9025 1.38 35.185 2.33 ;
      RECT  34.9025 2.33 35.185 2.745 ;
      RECT  34.9025 2.745 35.185 17.1975 ;
      RECT  65.8275 26.7175 66.2425 79.57 ;
      RECT  38.0775 26.7175 57.5475 79.57 ;
      RECT  57.5475 26.7175 65.8275 79.57 ;
      RECT  25.0775 26.7175 25.3575 31.73 ;
      RECT  25.3575 26.7175 34.77 31.73 ;
      RECT  34.77 26.7175 35.185 81.8275 ;
      RECT  35.185 26.7175 37.6625 81.8275 ;
      RECT  37.6625 26.7175 38.0775 81.8275 ;
      RECT  15.1275 47.095 15.4725 49.67 ;
      RECT  15.1275 50.085 15.4725 52.27 ;
      RECT  15.4725 47.095 15.5425 49.67 ;
      RECT  15.4725 50.085 15.5425 52.27 ;
      RECT  65.8275 1.38 66.2425 14.41 ;
      RECT  65.8275 14.825 66.2425 16.23 ;
      RECT  79.3425 42.195 80.735 42.61 ;
      RECT  79.3425 42.61 80.735 43.69 ;
      RECT  80.735 42.61 81.15 43.69 ;
      RECT  81.15 29.545 85.22 42.195 ;
      RECT  81.15 42.195 85.22 42.61 ;
      RECT  81.15 42.61 85.22 43.69 ;
      RECT  9.445 44.105 13.32 45.185 ;
      RECT  9.445 45.185 13.32 45.6 ;
      RECT  9.445 45.6 13.32 52.27 ;
      RECT  13.32 44.105 13.735 45.185 ;
      RECT  13.735 44.105 15.1275 45.185 ;
      RECT  13.735 45.185 15.1275 45.6 ;
      RECT  13.735 45.6 15.1275 52.27 ;
      RECT  24.9425 1.38 25.3575 14.41 ;
      RECT  24.9425 14.825 25.3575 16.23 ;
      RECT  9.445 32.145 13.945 36.215 ;
      RECT  9.445 36.215 13.945 36.63 ;
      RECT  13.945 36.63 14.36 43.69 ;
      RECT  14.36 32.145 15.1275 36.215 ;
      RECT  14.36 36.215 15.1275 36.63 ;
      RECT  14.36 36.63 15.1275 43.69 ;
      RECT  25.0775 87.9175 28.2625 89.46 ;
      RECT  28.2625 87.9175 28.6775 89.46 ;
      RECT  28.6775 87.9175 34.77 89.46 ;
      RECT  38.0775 87.9175 57.5475 89.46 ;
      RECT  57.5475 87.9175 57.5825 89.46 ;
      RECT  57.5825 87.5675 67.4175 87.9175 ;
      RECT  57.5825 87.9175 67.4175 89.46 ;
      RECT  34.77 87.9175 35.185 89.46 ;
      RECT  35.185 87.9175 37.6625 89.46 ;
      RECT  37.6625 87.9175 38.0775 89.46 ;
      RECT  25.0775 82.1775 28.2625 84.4475 ;
      RECT  25.0775 84.7975 28.2625 87.5675 ;
      RECT  28.2625 82.1775 28.6775 84.4475 ;
      RECT  28.2625 84.7975 28.6775 87.5675 ;
      RECT  28.6775 82.1775 34.77 84.4475 ;
      RECT  28.6775 84.7975 34.77 87.5675 ;
      RECT  38.0775 82.1775 57.5475 84.4475 ;
      RECT  38.0775 84.7975 57.5475 87.5675 ;
      RECT  57.5475 82.1775 57.5825 84.4475 ;
      RECT  57.5475 84.7975 57.5825 87.5675 ;
      RECT  57.5825 82.1775 66.275 84.4475 ;
      RECT  57.5825 84.7975 66.275 87.5675 ;
      RECT  66.275 82.1775 67.4175 84.4475 ;
      RECT  66.275 84.4475 67.4175 84.7975 ;
      RECT  66.275 84.7975 67.4175 87.5675 ;
      RECT  34.77 82.1775 35.185 84.4475 ;
      RECT  34.77 84.7975 35.185 87.5675 ;
      RECT  35.185 82.1775 37.6625 84.4475 ;
      RECT  35.185 84.7975 37.6625 87.5675 ;
      RECT  37.6625 82.1775 38.0775 84.4475 ;
      RECT  37.6625 84.7975 38.0775 87.5675 ;
      RECT  35.185 106.66 74.0625 107.35 ;
      RECT  35.185 107.35 74.0625 107.485 ;
      RECT  74.0625 106.66 74.4775 107.35 ;
      RECT  74.4775 106.66 76.64 107.35 ;
      RECT  74.4775 107.35 76.64 107.485 ;
      RECT  38.0775 17.5475 57.5475 19.2475 ;
      RECT  25.0775 17.5475 25.3575 19.2475 ;
      RECT  25.3575 17.5475 34.77 19.2475 ;
      RECT  34.77 17.5475 35.185 19.2475 ;
      RECT  35.185 17.5475 37.6625 19.2475 ;
      RECT  37.6625 17.5475 38.0775 19.2475 ;
      RECT  79.3425 44.105 80.735 48.175 ;
      RECT  79.3425 48.175 80.735 48.59 ;
      RECT  79.3425 48.59 80.735 106.245 ;
      RECT  81.15 44.105 85.22 48.175 ;
      RECT  81.15 48.175 85.22 48.59 ;
      RECT  81.15 48.59 85.22 106.245 ;
      RECT  9.445 36.63 13.32 39.205 ;
      RECT  9.445 39.205 13.32 39.62 ;
      RECT  9.445 39.62 13.32 43.69 ;
      RECT  13.32 36.63 13.735 39.205 ;
      RECT  13.735 36.63 13.945 39.205 ;
      RECT  13.735 39.205 13.945 39.62 ;
      RECT  13.735 39.62 13.945 43.69 ;
      RECT  80.735 48.59 81.15 51.165 ;
      RECT  80.735 51.58 81.15 106.245 ;
      RECT  79.3425 29.545 80.11 33.225 ;
      RECT  79.3425 33.225 80.11 33.64 ;
      RECT  79.3425 33.64 80.11 42.195 ;
      RECT  80.525 29.545 80.735 33.225 ;
      RECT  80.525 33.225 80.735 33.64 ;
      RECT  80.525 33.64 80.735 42.195 ;
      RECT  13.32 39.62 13.735 42.195 ;
      RECT  13.32 42.61 13.735 43.69 ;
      RECT  80.735 44.105 81.15 45.185 ;
      RECT  80.735 45.6 81.15 48.175 ;
      RECT  66.2425 16.645 66.275 23.7475 ;
      RECT  66.2425 24.0975 66.275 79.57 ;
      RECT  66.275 16.645 70.1225 23.7475 ;
      RECT  66.275 23.7475 70.1225 24.0975 ;
      RECT  66.275 24.0975 70.1225 79.57 ;
      RECT  65.8275 16.645 66.2425 23.7475 ;
      RECT  65.8275 24.0975 66.2425 26.3675 ;
      RECT  57.5475 17.5475 65.8275 23.7475 ;
      RECT  57.5475 24.0975 65.8275 26.3675 ;
      RECT  38.0775 19.5975 57.5475 23.7475 ;
      RECT  38.0775 24.0975 57.5475 26.3675 ;
      RECT  25.0775 19.5975 25.3575 23.7475 ;
      RECT  25.0775 24.0975 25.3575 26.3675 ;
      RECT  25.3575 19.5975 34.77 23.7475 ;
      RECT  25.3575 24.0975 34.77 26.3675 ;
      RECT  34.77 19.5975 35.185 23.7475 ;
      RECT  34.77 24.0975 35.185 26.3675 ;
      RECT  35.185 19.5975 37.6625 23.7475 ;
      RECT  35.185 24.0975 37.6625 26.3675 ;
      RECT  37.6625 19.5975 38.0775 23.7475 ;
      RECT  37.6625 24.0975 38.0775 26.3675 ;
      RECT  0.14 0.14 17.3275 0.275 ;
      RECT  0.14 0.275 17.3275 0.965 ;
      RECT  17.3275 0.275 17.7425 0.965 ;
      RECT  17.7425 0.275 34.77 0.965 ;
      RECT  9.445 2.745 13.945 30.235 ;
      RECT  9.445 30.235 13.945 30.65 ;
      RECT  9.445 30.65 13.945 31.73 ;
      RECT  13.945 2.745 14.36 30.235 ;
      RECT  13.945 30.65 14.36 31.73 ;
      RECT  14.36 2.745 14.4675 30.235 ;
      RECT  14.36 30.235 14.4675 30.65 ;
      RECT  14.36 30.65 14.4675 31.73 ;
      RECT  17.7425 0.14 25.9075 0.275 ;
      RECT  26.3225 0.14 34.77 0.275 ;
      RECT  13.945 32.145 14.36 33.225 ;
      RECT  13.945 33.64 14.36 36.215 ;
      RECT  13.32 45.6 13.735 48.175 ;
      RECT  80.11 33.64 80.525 36.215 ;
      RECT  80.11 36.63 80.525 42.195 ;
      RECT  13.32 48.59 13.735 51.165 ;
      RECT  13.32 51.58 13.735 52.27 ;
      RECT  85.635 95.405 92.105 96.095 ;
      RECT  85.635 96.095 92.105 96.51 ;
      RECT  85.635 96.51 92.105 106.245 ;
      RECT  92.105 95.405 92.52 96.095 ;
      RECT  92.105 96.51 92.52 106.245 ;
      RECT  92.52 95.405 94.245 96.095 ;
      RECT  92.52 96.095 94.245 96.51 ;
      RECT  92.52 96.51 94.245 106.245 ;
      RECT  80.11 29.545 80.525 30.235 ;
      RECT  80.11 30.65 80.525 33.225 ;
      RECT  0.56 1.38 2.285 9.565 ;
      RECT  0.56 9.565 2.285 9.98 ;
      RECT  0.56 9.98 2.285 10.67 ;
      RECT  2.285 1.38 2.7 9.565 ;
      RECT  2.285 9.98 2.7 10.67 ;
      RECT  2.7 1.38 9.03 9.565 ;
      RECT  2.7 9.565 9.03 9.98 ;
      RECT  2.7 9.98 9.03 10.67 ;
      RECT  35.185 0.14 37.3475 0.275 ;
      RECT  35.185 0.275 37.3475 0.965 ;
      RECT  37.3475 0.275 37.7625 0.965 ;
      RECT  37.7625 0.14 94.665 0.275 ;
      RECT  37.7625 0.275 94.665 0.965 ;
      RECT  80.735 29.545 81.15 39.205 ;
      RECT  80.735 39.62 81.15 42.195 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 0.4075 19.27 ;
      RECT  0.14 19.27 0.4075 42.2325 ;
      RECT  0.14 42.2325 0.4075 107.485 ;
      RECT  0.4075 0.14 1.1075 19.27 ;
      RECT  0.4075 42.2325 1.1075 107.485 ;
      RECT  82.64 42.2325 83.34 83.6025 ;
      RECT  82.64 94.1825 83.34 107.485 ;
      RECT  85.36 0.14 86.06 17.6775 ;
      RECT  86.06 0.14 94.665 17.6775 ;
      RECT  86.06 17.6775 94.665 19.27 ;
      RECT  85.36 30.7925 86.06 42.2325 ;
      RECT  86.06 19.27 94.665 30.7925 ;
      RECT  86.06 30.7925 94.665 42.2325 ;
      RECT  69.98 78.6325 70.68 83.6025 ;
      RECT  69.98 19.27 70.68 30.0925 ;
      RECT  69.6 42.2325 69.98 78.6325 ;
      RECT  1.1075 81.5525 68.9 83.6025 ;
      RECT  68.9 81.5525 69.6 83.6025 ;
      RECT  69.6 78.6325 69.98 81.5525 ;
      RECT  69.6 81.5525 69.98 83.6025 ;
      RECT  68.9 19.27 69.6 26.9225 ;
      RECT  69.6 19.27 69.98 26.9225 ;
      RECT  69.6 26.9225 69.98 30.0925 ;
      RECT  69.6 30.0925 69.98 30.7925 ;
      RECT  69.6 30.7925 69.98 42.2325 ;
      RECT  1.1075 78.7025 20.54 81.5525 ;
      RECT  20.54 78.7025 21.24 81.5525 ;
      RECT  17.92 0.14 18.62 4.005 ;
      RECT  18.62 0.14 85.36 4.005 ;
      RECT  18.62 4.005 85.36 17.6775 ;
      RECT  17.92 24.465 18.62 26.9225 ;
      RECT  18.62 19.27 68.9 24.465 ;
      RECT  18.62 24.465 68.9 26.9225 ;
      RECT  93.6975 42.2325 94.3975 63.8425 ;
      RECT  94.3975 42.2325 94.665 63.8425 ;
      RECT  94.3975 63.8425 94.665 83.6025 ;
      RECT  93.6975 86.805 94.3975 94.1825 ;
      RECT  94.3975 83.6025 94.665 86.805 ;
      RECT  94.3975 86.805 94.665 94.1825 ;
      RECT  1.1075 83.6025 75.85 84.08 ;
      RECT  1.1075 84.08 75.85 94.1825 ;
      RECT  75.85 83.6025 76.55 84.08 ;
      RECT  1.1075 94.1825 75.85 104.54 ;
      RECT  1.1075 104.54 75.85 107.485 ;
      RECT  75.85 104.54 76.55 107.485 ;
      RECT  70.68 78.7025 73.23 83.6025 ;
      RECT  73.23 78.7025 73.93 83.6025 ;
      RECT  73.93 78.7025 82.64 83.6025 ;
      RECT  11.325 27.4125 12.025 30.0925 ;
      RECT  11.325 4.005 12.025 11.8925 ;
      RECT  21.24 78.7025 24.87 81.5525 ;
      RECT  24.49 42.2325 24.87 78.6325 ;
      RECT  24.49 30.0925 24.87 30.7925 ;
      RECT  24.49 30.7925 24.87 42.2325 ;
      RECT  12.025 26.9225 24.87 27.4125 ;
      RECT  1.1075 51.0225 8.605 64.1375 ;
      RECT  1.1075 64.1375 8.605 78.6325 ;
      RECT  8.605 42.2325 9.305 51.0225 ;
      RECT  8.605 64.1375 9.305 78.6325 ;
      RECT  83.2 19.27 85.36 30.0925 ;
      RECT  18.62 17.6775 82.5 17.7425 ;
      RECT  18.62 17.7425 82.5 19.27 ;
      RECT  82.5 17.6775 83.2 17.7425 ;
      RECT  83.2 17.6775 85.36 17.7425 ;
      RECT  83.2 17.7425 85.36 19.27 ;
      RECT  83.2 30.0925 85.36 30.7925 ;
      RECT  82.5 30.8575 83.2 42.2325 ;
      RECT  83.2 30.7925 85.36 30.8575 ;
      RECT  83.2 30.8575 85.36 42.2325 ;
      RECT  1.1075 78.6325 18.95 78.7025 ;
      RECT  19.65 78.6325 20.54 78.7025 ;
      RECT  19.65 30.0925 20.54 30.7925 ;
      RECT  19.65 30.7925 20.54 42.2325 ;
      RECT  12.025 27.4125 18.95 30.06 ;
      RECT  12.025 30.06 18.95 30.0925 ;
      RECT  18.95 27.4125 19.65 30.06 ;
      RECT  19.65 27.4125 24.87 30.06 ;
      RECT  19.65 42.2325 20.54 51.0225 ;
      RECT  19.65 51.0225 20.54 64.1375 ;
      RECT  9.305 64.1375 18.95 78.6325 ;
      RECT  19.65 64.1375 20.54 78.6325 ;
      RECT  1.1075 4.005 5.825 9.4225 ;
      RECT  1.1075 9.4225 5.825 11.8925 ;
      RECT  5.825 4.005 6.525 9.4225 ;
      RECT  6.525 4.005 11.325 9.4225 ;
      RECT  6.525 9.4225 11.325 11.8925 ;
      RECT  1.1075 11.8925 5.825 17.6775 ;
      RECT  6.525 11.8925 11.325 17.6775 ;
      RECT  1.1075 17.6775 5.825 19.27 ;
      RECT  6.525 17.6775 11.325 19.27 ;
      RECT  6.525 19.27 11.325 24.465 ;
      RECT  5.825 24.9425 6.525 26.9225 ;
      RECT  6.525 24.465 11.325 24.9425 ;
      RECT  6.525 24.9425 11.325 26.9225 ;
      RECT  70.68 42.2325 72.67 78.6325 ;
      RECT  70.68 78.6325 72.67 78.665 ;
      RECT  70.68 78.665 72.67 78.7025 ;
      RECT  72.67 78.665 73.23 78.7025 ;
      RECT  70.68 30.0925 72.67 30.7925 ;
      RECT  70.68 30.7925 72.67 42.2325 ;
      RECT  70.68 19.27 72.67 30.06 ;
      RECT  70.68 30.06 72.67 30.0925 ;
      RECT  72.67 19.27 73.37 30.06 ;
      RECT  73.37 19.27 82.5 30.06 ;
      RECT  76.55 83.6025 77.7925 84.0125 ;
      RECT  76.55 84.0125 77.7925 84.08 ;
      RECT  77.7925 83.6025 78.4925 84.0125 ;
      RECT  78.4925 83.6025 82.64 84.0125 ;
      RECT  78.4925 84.0125 82.64 84.08 ;
      RECT  76.55 84.08 77.7925 94.1825 ;
      RECT  78.4925 84.08 82.64 94.1825 ;
      RECT  76.55 94.1825 77.7925 104.54 ;
      RECT  78.4925 94.1825 82.64 104.54 ;
      RECT  76.55 104.54 77.7925 104.6075 ;
      RECT  76.55 104.6075 77.7925 107.485 ;
      RECT  77.7925 104.6075 78.4925 107.485 ;
      RECT  78.4925 104.54 82.64 104.6075 ;
      RECT  78.4925 104.6075 82.64 107.485 ;
      RECT  9.305 42.2325 11.465 50.9575 ;
      RECT  9.305 50.9575 11.465 51.0225 ;
      RECT  11.465 42.2325 12.165 50.9575 ;
      RECT  12.165 42.2325 18.95 50.9575 ;
      RECT  12.165 50.9575 18.95 51.0225 ;
      RECT  9.305 51.0225 11.465 64.0725 ;
      RECT  9.305 64.0725 11.465 64.1375 ;
      RECT  11.465 64.0725 12.165 64.1375 ;
      RECT  12.165 51.0225 18.95 64.0725 ;
      RECT  12.165 64.0725 18.95 64.1375 ;
      RECT  73.93 42.2325 74.82 78.6325 ;
      RECT  75.52 42.2325 82.64 78.6325 ;
      RECT  73.93 78.6325 74.82 78.7025 ;
      RECT  75.52 78.6325 82.64 78.7025 ;
      RECT  73.93 30.0925 74.82 30.7925 ;
      RECT  75.52 30.0925 82.5 30.7925 ;
      RECT  73.93 30.7925 74.82 30.8575 ;
      RECT  75.52 30.7925 82.5 30.8575 ;
      RECT  73.93 30.8575 74.82 42.2325 ;
      RECT  75.52 30.8575 82.5 42.2325 ;
      RECT  73.37 30.06 74.82 30.0925 ;
      RECT  75.52 30.06 82.5 30.0925 ;
      RECT  83.34 42.2325 91.635 63.81 ;
      RECT  83.34 63.81 91.635 63.8425 ;
      RECT  91.635 42.2325 92.335 63.81 ;
      RECT  92.335 42.2325 93.6975 63.81 ;
      RECT  92.335 63.81 93.6975 63.8425 ;
      RECT  92.335 63.8425 93.6975 83.6025 ;
      RECT  91.635 86.7725 92.335 86.805 ;
      RECT  92.335 83.6025 93.6975 86.7725 ;
      RECT  92.335 86.7725 93.6975 86.805 ;
      RECT  26.03 78.6325 68.44 78.7025 ;
      RECT  26.03 78.7025 68.44 81.5525 ;
      RECT  26.03 42.2325 68.44 78.6325 ;
      RECT  26.03 30.0925 68.44 30.7925 ;
      RECT  26.03 30.7925 68.44 42.2325 ;
      RECT  26.03 26.9225 68.44 27.4125 ;
      RECT  26.03 27.4125 68.44 30.0925 ;
      RECT  1.1075 26.9225 2.47 27.4125 ;
      RECT  3.17 26.9225 11.325 27.4125 ;
      RECT  1.1075 27.4125 2.47 30.0925 ;
      RECT  3.17 27.4125 11.325 30.0925 ;
      RECT  1.1075 42.2325 2.47 42.265 ;
      RECT  1.1075 42.265 2.47 51.0225 ;
      RECT  2.47 42.265 3.17 51.0225 ;
      RECT  3.17 42.2325 8.605 42.265 ;
      RECT  3.17 42.265 8.605 51.0225 ;
      RECT  1.1075 30.0925 2.47 30.7925 ;
      RECT  3.17 30.0925 18.95 30.7925 ;
      RECT  1.1075 30.7925 2.47 42.2325 ;
      RECT  3.17 30.7925 18.95 42.2325 ;
      RECT  1.1075 19.27 2.47 19.3025 ;
      RECT  1.1075 19.3025 2.47 24.465 ;
      RECT  2.47 19.27 3.17 19.3025 ;
      RECT  3.17 19.27 5.825 19.3025 ;
      RECT  3.17 19.3025 5.825 24.465 ;
      RECT  1.1075 24.465 2.47 24.9425 ;
      RECT  3.17 24.465 5.825 24.9425 ;
      RECT  1.1075 24.9425 2.47 26.9225 ;
      RECT  3.17 24.9425 5.825 26.9225 ;
      RECT  21.8 42.2325 23.79 78.6325 ;
      RECT  21.8 30.0925 23.79 30.7925 ;
      RECT  21.8 30.7925 23.79 42.2325 ;
      RECT  21.24 78.665 21.8 78.7025 ;
      RECT  21.8 78.6325 24.87 78.665 ;
      RECT  21.8 78.665 24.87 78.7025 ;
      RECT  19.65 30.06 21.1 30.0925 ;
      RECT  21.8 30.06 24.87 30.0925 ;
      RECT  83.34 94.1825 88.14 96.6525 ;
      RECT  83.34 96.6525 88.14 107.485 ;
      RECT  88.14 96.6525 88.84 107.485 ;
      RECT  88.84 94.1825 94.665 96.6525 ;
      RECT  88.84 96.6525 94.665 107.485 ;
      RECT  83.34 86.805 88.14 94.1825 ;
      RECT  88.84 86.805 93.6975 94.1825 ;
      RECT  83.34 63.8425 88.14 81.1325 ;
      RECT  83.34 81.1325 88.14 83.6025 ;
      RECT  88.14 63.8425 88.84 81.1325 ;
      RECT  88.84 63.8425 91.635 81.1325 ;
      RECT  88.84 81.1325 91.635 83.6025 ;
      RECT  83.34 83.6025 88.14 86.7725 ;
      RECT  88.84 83.6025 91.635 86.7725 ;
      RECT  83.34 86.7725 88.14 86.805 ;
      RECT  88.84 86.7725 91.635 86.805 ;
      RECT  1.1075 0.14 15.9775 3.9375 ;
      RECT  1.1075 3.9375 15.9775 4.005 ;
      RECT  15.9775 0.14 16.6775 3.9375 ;
      RECT  16.6775 0.14 17.92 3.9375 ;
      RECT  16.6775 3.9375 17.92 4.005 ;
      RECT  12.025 4.005 15.9775 11.8925 ;
      RECT  16.6775 4.005 17.92 11.8925 ;
      RECT  12.025 11.8925 15.9775 17.6775 ;
      RECT  16.6775 11.8925 17.92 17.6775 ;
      RECT  12.025 17.6775 15.9775 19.27 ;
      RECT  16.6775 17.6775 17.92 19.27 ;
      RECT  12.025 19.27 15.9775 24.465 ;
      RECT  16.6775 19.27 17.92 24.465 ;
      RECT  12.025 24.465 15.9775 24.5325 ;
      RECT  12.025 24.5325 15.9775 26.9225 ;
      RECT  15.9775 24.5325 16.6775 26.9225 ;
      RECT  16.6775 24.465 17.92 24.5325 ;
      RECT  16.6775 24.5325 17.92 26.9225 ;
   END
END    freepdk45_sram_1w1r_256x4_1
END    LIBRARY
