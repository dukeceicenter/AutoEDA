../macros/freepdk45_sram_1rw0r_64x176_22/freepdk45_sram_1rw0r_64x176_22.lef