VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_32x240
   CLASS BLOCK ;
   SIZE 752.775 BY 116.3125 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.59 1.105 66.725 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.45 1.105 69.585 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.31 1.105 72.445 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.17 1.105 75.305 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.03 1.105 78.165 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.89 1.105 81.025 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.75 1.105 83.885 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.61 1.105 86.745 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.47 1.105 89.605 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.33 1.105 92.465 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.19 1.105 95.325 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.05 1.105 98.185 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.91 1.105 101.045 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.77 1.105 103.905 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.63 1.105 106.765 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.49 1.105 109.625 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.35 1.105 112.485 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.21 1.105 115.345 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.07 1.105 118.205 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.93 1.105 121.065 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.79 1.105 123.925 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.65 1.105 126.785 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.51 1.105 129.645 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.37 1.105 132.505 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.23 1.105 135.365 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.09 1.105 138.225 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.95 1.105 141.085 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.81 1.105 143.945 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.67 1.105 146.805 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.53 1.105 149.665 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.39 1.105 152.525 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.25 1.105 155.385 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.11 1.105 158.245 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.97 1.105 161.105 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.83 1.105 163.965 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.69 1.105 166.825 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.55 1.105 169.685 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.41 1.105 172.545 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.27 1.105 175.405 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.13 1.105 178.265 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.99 1.105 181.125 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.85 1.105 183.985 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.71 1.105 186.845 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.57 1.105 189.705 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.43 1.105 192.565 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.29 1.105 195.425 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.15 1.105 198.285 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.01 1.105 201.145 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.87 1.105 204.005 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.73 1.105 206.865 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.59 1.105 209.725 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.45 1.105 212.585 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.31 1.105 215.445 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.17 1.105 218.305 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.03 1.105 221.165 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.89 1.105 224.025 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.75 1.105 226.885 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.61 1.105 229.745 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.47 1.105 232.605 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.33 1.105 235.465 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.19 1.105 238.325 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.05 1.105 241.185 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.91 1.105 244.045 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.77 1.105 246.905 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.63 1.105 249.765 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.49 1.105 252.625 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.35 1.105 255.485 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.21 1.105 258.345 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.07 1.105 261.205 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.93 1.105 264.065 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.79 1.105 266.925 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.65 1.105 269.785 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.51 1.105 272.645 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.37 1.105 275.505 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.23 1.105 278.365 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.09 1.105 281.225 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.95 1.105 284.085 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.81 1.105 286.945 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.67 1.105 289.805 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.53 1.105 292.665 1.24 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.39 1.105 295.525 1.24 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.25 1.105 298.385 1.24 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.11 1.105 301.245 1.24 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.97 1.105 304.105 1.24 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.83 1.105 306.965 1.24 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.69 1.105 309.825 1.24 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.55 1.105 312.685 1.24 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.41 1.105 315.545 1.24 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.27 1.105 318.405 1.24 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.13 1.105 321.265 1.24 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.99 1.105 324.125 1.24 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.85 1.105 326.985 1.24 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.71 1.105 329.845 1.24 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.57 1.105 332.705 1.24 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.43 1.105 335.565 1.24 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.29 1.105 338.425 1.24 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.15 1.105 341.285 1.24 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.01 1.105 344.145 1.24 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.87 1.105 347.005 1.24 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.73 1.105 349.865 1.24 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.59 1.105 352.725 1.24 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.45 1.105 355.585 1.24 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.31 1.105 358.445 1.24 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.17 1.105 361.305 1.24 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.03 1.105 364.165 1.24 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.89 1.105 367.025 1.24 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.75 1.105 369.885 1.24 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.61 1.105 372.745 1.24 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.47 1.105 375.605 1.24 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.33 1.105 378.465 1.24 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.19 1.105 381.325 1.24 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.05 1.105 384.185 1.24 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.91 1.105 387.045 1.24 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.77 1.105 389.905 1.24 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.63 1.105 392.765 1.24 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.49 1.105 395.625 1.24 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.35 1.105 398.485 1.24 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.21 1.105 401.345 1.24 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.07 1.105 404.205 1.24 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.93 1.105 407.065 1.24 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.79 1.105 409.925 1.24 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.65 1.105 412.785 1.24 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.51 1.105 415.645 1.24 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.37 1.105 418.505 1.24 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.23 1.105 421.365 1.24 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.09 1.105 424.225 1.24 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.95 1.105 427.085 1.24 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.81 1.105 429.945 1.24 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.67 1.105 432.805 1.24 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.53 1.105 435.665 1.24 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.39 1.105 438.525 1.24 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.25 1.105 441.385 1.24 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.11 1.105 444.245 1.24 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.97 1.105 447.105 1.24 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.83 1.105 449.965 1.24 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.69 1.105 452.825 1.24 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.55 1.105 455.685 1.24 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.41 1.105 458.545 1.24 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.27 1.105 461.405 1.24 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.13 1.105 464.265 1.24 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.99 1.105 467.125 1.24 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.85 1.105 469.985 1.24 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.71 1.105 472.845 1.24 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.57 1.105 475.705 1.24 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.43 1.105 478.565 1.24 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.29 1.105 481.425 1.24 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.15 1.105 484.285 1.24 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.01 1.105 487.145 1.24 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.87 1.105 490.005 1.24 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.73 1.105 492.865 1.24 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.59 1.105 495.725 1.24 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.45 1.105 498.585 1.24 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.31 1.105 501.445 1.24 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.17 1.105 504.305 1.24 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.03 1.105 507.165 1.24 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.89 1.105 510.025 1.24 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.75 1.105 512.885 1.24 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.61 1.105 515.745 1.24 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.47 1.105 518.605 1.24 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.33 1.105 521.465 1.24 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  524.19 1.105 524.325 1.24 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.05 1.105 527.185 1.24 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  529.91 1.105 530.045 1.24 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  532.77 1.105 532.905 1.24 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  535.63 1.105 535.765 1.24 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  538.49 1.105 538.625 1.24 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  541.35 1.105 541.485 1.24 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  544.21 1.105 544.345 1.24 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  547.07 1.105 547.205 1.24 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  549.93 1.105 550.065 1.24 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  552.79 1.105 552.925 1.24 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  555.65 1.105 555.785 1.24 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  558.51 1.105 558.645 1.24 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  561.37 1.105 561.505 1.24 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  564.23 1.105 564.365 1.24 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  567.09 1.105 567.225 1.24 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  569.95 1.105 570.085 1.24 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  572.81 1.105 572.945 1.24 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  575.67 1.105 575.805 1.24 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  578.53 1.105 578.665 1.24 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  581.39 1.105 581.525 1.24 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  584.25 1.105 584.385 1.24 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  587.11 1.105 587.245 1.24 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  589.97 1.105 590.105 1.24 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  592.83 1.105 592.965 1.24 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  595.69 1.105 595.825 1.24 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  598.55 1.105 598.685 1.24 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  601.41 1.105 601.545 1.24 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  604.27 1.105 604.405 1.24 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  607.13 1.105 607.265 1.24 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  609.99 1.105 610.125 1.24 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  612.85 1.105 612.985 1.24 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  615.71 1.105 615.845 1.24 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  618.57 1.105 618.705 1.24 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  621.43 1.105 621.565 1.24 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  624.29 1.105 624.425 1.24 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  627.15 1.105 627.285 1.24 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  630.01 1.105 630.145 1.24 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  632.87 1.105 633.005 1.24 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  635.73 1.105 635.865 1.24 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  638.59 1.105 638.725 1.24 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  641.45 1.105 641.585 1.24 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  644.31 1.105 644.445 1.24 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  647.17 1.105 647.305 1.24 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  650.03 1.105 650.165 1.24 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  652.89 1.105 653.025 1.24 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  655.75 1.105 655.885 1.24 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  658.61 1.105 658.745 1.24 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  661.47 1.105 661.605 1.24 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  664.33 1.105 664.465 1.24 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  667.19 1.105 667.325 1.24 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  670.05 1.105 670.185 1.24 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  672.91 1.105 673.045 1.24 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  675.77 1.105 675.905 1.24 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  678.63 1.105 678.765 1.24 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  681.49 1.105 681.625 1.24 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  684.35 1.105 684.485 1.24 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  687.21 1.105 687.345 1.24 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  690.07 1.105 690.205 1.24 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  692.93 1.105 693.065 1.24 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  695.79 1.105 695.925 1.24 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  698.65 1.105 698.785 1.24 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  701.51 1.105 701.645 1.24 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  704.37 1.105 704.505 1.24 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  707.23 1.105 707.365 1.24 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  710.09 1.105 710.225 1.24 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  712.95 1.105 713.085 1.24 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  715.81 1.105 715.945 1.24 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  718.67 1.105 718.805 1.24 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  721.53 1.105 721.665 1.24 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  724.39 1.105 724.525 1.24 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  727.25 1.105 727.385 1.24 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  730.11 1.105 730.245 1.24 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  732.97 1.105 733.105 1.24 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  735.83 1.105 735.965 1.24 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  738.69 1.105 738.825 1.24 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  741.55 1.105 741.685 1.24 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  744.41 1.105 744.545 1.24 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  747.27 1.105 747.405 1.24 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  750.13 1.105 750.265 1.24 ;
      END
   END din0[239]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 72.35 61.005 72.485 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 75.08 61.005 75.215 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 77.29 61.005 77.425 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 80.02 61.005 80.155 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.87 82.23 61.005 82.365 ;
      END
   END addr0[4]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.61 49.21 399.745 49.345 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.61 46.48 399.745 46.615 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.61 44.27 399.745 44.405 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.61 41.54 399.745 41.675 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.61 39.33 399.745 39.465 ;
      END
   END addr1[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 30.75 0.42 30.885 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  460.335 115.07 460.47 115.205 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 30.835 6.3825 30.97 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  454.2325 114.985 454.3675 115.12 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.1775 108.3625 89.3125 108.4975 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.3525 108.3625 90.4875 108.4975 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.5275 108.3625 91.6625 108.4975 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.7025 108.3625 92.8375 108.4975 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.8775 108.3625 94.0125 108.4975 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.0525 108.3625 95.1875 108.4975 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.2275 108.3625 96.3625 108.4975 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.4025 108.3625 97.5375 108.4975 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.5775 108.3625 98.7125 108.4975 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.7525 108.3625 99.8875 108.4975 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.9275 108.3625 101.0625 108.4975 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.1025 108.3625 102.2375 108.4975 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.2775 108.3625 103.4125 108.4975 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.4525 108.3625 104.5875 108.4975 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.6275 108.3625 105.7625 108.4975 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.8025 108.3625 106.9375 108.4975 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.9775 108.3625 108.1125 108.4975 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.1525 108.3625 109.2875 108.4975 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.3275 108.3625 110.4625 108.4975 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.5025 108.3625 111.6375 108.4975 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.6775 108.3625 112.8125 108.4975 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.8525 108.3625 113.9875 108.4975 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.0275 108.3625 115.1625 108.4975 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.2025 108.3625 116.3375 108.4975 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.3775 108.3625 117.5125 108.4975 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.5525 108.3625 118.6875 108.4975 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.7275 108.3625 119.8625 108.4975 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.9025 108.3625 121.0375 108.4975 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.0775 108.3625 122.2125 108.4975 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.2525 108.3625 123.3875 108.4975 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.4275 108.3625 124.5625 108.4975 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.6025 108.3625 125.7375 108.4975 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.7775 108.3625 126.9125 108.4975 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.9525 108.3625 128.0875 108.4975 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.1275 108.3625 129.2625 108.4975 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.3025 108.3625 130.4375 108.4975 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.4775 108.3625 131.6125 108.4975 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.6525 108.3625 132.7875 108.4975 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.8275 108.3625 133.9625 108.4975 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.0025 108.3625 135.1375 108.4975 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.1775 108.3625 136.3125 108.4975 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.3525 108.3625 137.4875 108.4975 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.5275 108.3625 138.6625 108.4975 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.7025 108.3625 139.8375 108.4975 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.8775 108.3625 141.0125 108.4975 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.0525 108.3625 142.1875 108.4975 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.2275 108.3625 143.3625 108.4975 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.4025 108.3625 144.5375 108.4975 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.5775 108.3625 145.7125 108.4975 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.7525 108.3625 146.8875 108.4975 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.9275 108.3625 148.0625 108.4975 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.1025 108.3625 149.2375 108.4975 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.2775 108.3625 150.4125 108.4975 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.4525 108.3625 151.5875 108.4975 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.6275 108.3625 152.7625 108.4975 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.8025 108.3625 153.9375 108.4975 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.9775 108.3625 155.1125 108.4975 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.1525 108.3625 156.2875 108.4975 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.3275 108.3625 157.4625 108.4975 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.5025 108.3625 158.6375 108.4975 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.6775 108.3625 159.8125 108.4975 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.8525 108.3625 160.9875 108.4975 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.0275 108.3625 162.1625 108.4975 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.2025 108.3625 163.3375 108.4975 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.3775 108.3625 164.5125 108.4975 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.5525 108.3625 165.6875 108.4975 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.7275 108.3625 166.8625 108.4975 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.9025 108.3625 168.0375 108.4975 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.0775 108.3625 169.2125 108.4975 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.2525 108.3625 170.3875 108.4975 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.4275 108.3625 171.5625 108.4975 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.6025 108.3625 172.7375 108.4975 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.7775 108.3625 173.9125 108.4975 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.9525 108.3625 175.0875 108.4975 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.1275 108.3625 176.2625 108.4975 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.3025 108.3625 177.4375 108.4975 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.4775 108.3625 178.6125 108.4975 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.6525 108.3625 179.7875 108.4975 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.8275 108.3625 180.9625 108.4975 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.0025 108.3625 182.1375 108.4975 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.1775 108.3625 183.3125 108.4975 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.3525 108.3625 184.4875 108.4975 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.5275 108.3625 185.6625 108.4975 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.7025 108.3625 186.8375 108.4975 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.8775 108.3625 188.0125 108.4975 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.0525 108.3625 189.1875 108.4975 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.2275 108.3625 190.3625 108.4975 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.4025 108.3625 191.5375 108.4975 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.5775 108.3625 192.7125 108.4975 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.7525 108.3625 193.8875 108.4975 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.9275 108.3625 195.0625 108.4975 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.1025 108.3625 196.2375 108.4975 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.2775 108.3625 197.4125 108.4975 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.4525 108.3625 198.5875 108.4975 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.6275 108.3625 199.7625 108.4975 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.8025 108.3625 200.9375 108.4975 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.9775 108.3625 202.1125 108.4975 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.1525 108.3625 203.2875 108.4975 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.3275 108.3625 204.4625 108.4975 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.5025 108.3625 205.6375 108.4975 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.6775 108.3625 206.8125 108.4975 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.8525 108.3625 207.9875 108.4975 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.0275 108.3625 209.1625 108.4975 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.2025 108.3625 210.3375 108.4975 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.3775 108.3625 211.5125 108.4975 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.5525 108.3625 212.6875 108.4975 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.7275 108.3625 213.8625 108.4975 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.9025 108.3625 215.0375 108.4975 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.0775 108.3625 216.2125 108.4975 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.2525 108.3625 217.3875 108.4975 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.4275 108.3625 218.5625 108.4975 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.6025 108.3625 219.7375 108.4975 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.7775 108.3625 220.9125 108.4975 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.9525 108.3625 222.0875 108.4975 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.1275 108.3625 223.2625 108.4975 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.3025 108.3625 224.4375 108.4975 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.4775 108.3625 225.6125 108.4975 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.6525 108.3625 226.7875 108.4975 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.8275 108.3625 227.9625 108.4975 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.0025 108.3625 229.1375 108.4975 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.1775 108.3625 230.3125 108.4975 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.3525 108.3625 231.4875 108.4975 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.5275 108.3625 232.6625 108.4975 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.7025 108.3625 233.8375 108.4975 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.8775 108.3625 235.0125 108.4975 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.0525 108.3625 236.1875 108.4975 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.2275 108.3625 237.3625 108.4975 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.4025 108.3625 238.5375 108.4975 ;
      END
   END dout1[127]
   PIN dout1[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.5775 108.3625 239.7125 108.4975 ;
      END
   END dout1[128]
   PIN dout1[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.7525 108.3625 240.8875 108.4975 ;
      END
   END dout1[129]
   PIN dout1[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.9275 108.3625 242.0625 108.4975 ;
      END
   END dout1[130]
   PIN dout1[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.1025 108.3625 243.2375 108.4975 ;
      END
   END dout1[131]
   PIN dout1[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.2775 108.3625 244.4125 108.4975 ;
      END
   END dout1[132]
   PIN dout1[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.4525 108.3625 245.5875 108.4975 ;
      END
   END dout1[133]
   PIN dout1[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.6275 108.3625 246.7625 108.4975 ;
      END
   END dout1[134]
   PIN dout1[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.8025 108.3625 247.9375 108.4975 ;
      END
   END dout1[135]
   PIN dout1[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.9775 108.3625 249.1125 108.4975 ;
      END
   END dout1[136]
   PIN dout1[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.1525 108.3625 250.2875 108.4975 ;
      END
   END dout1[137]
   PIN dout1[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.3275 108.3625 251.4625 108.4975 ;
      END
   END dout1[138]
   PIN dout1[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.5025 108.3625 252.6375 108.4975 ;
      END
   END dout1[139]
   PIN dout1[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.6775 108.3625 253.8125 108.4975 ;
      END
   END dout1[140]
   PIN dout1[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.8525 108.3625 254.9875 108.4975 ;
      END
   END dout1[141]
   PIN dout1[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.0275 108.3625 256.1625 108.4975 ;
      END
   END dout1[142]
   PIN dout1[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.2025 108.3625 257.3375 108.4975 ;
      END
   END dout1[143]
   PIN dout1[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.3775 108.3625 258.5125 108.4975 ;
      END
   END dout1[144]
   PIN dout1[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.5525 108.3625 259.6875 108.4975 ;
      END
   END dout1[145]
   PIN dout1[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.7275 108.3625 260.8625 108.4975 ;
      END
   END dout1[146]
   PIN dout1[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.9025 108.3625 262.0375 108.4975 ;
      END
   END dout1[147]
   PIN dout1[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.0775 108.3625 263.2125 108.4975 ;
      END
   END dout1[148]
   PIN dout1[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.2525 108.3625 264.3875 108.4975 ;
      END
   END dout1[149]
   PIN dout1[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.4275 108.3625 265.5625 108.4975 ;
      END
   END dout1[150]
   PIN dout1[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.6025 108.3625 266.7375 108.4975 ;
      END
   END dout1[151]
   PIN dout1[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.7775 108.3625 267.9125 108.4975 ;
      END
   END dout1[152]
   PIN dout1[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.9525 108.3625 269.0875 108.4975 ;
      END
   END dout1[153]
   PIN dout1[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.1275 108.3625 270.2625 108.4975 ;
      END
   END dout1[154]
   PIN dout1[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.3025 108.3625 271.4375 108.4975 ;
      END
   END dout1[155]
   PIN dout1[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.4775 108.3625 272.6125 108.4975 ;
      END
   END dout1[156]
   PIN dout1[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.6525 108.3625 273.7875 108.4975 ;
      END
   END dout1[157]
   PIN dout1[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.8275 108.3625 274.9625 108.4975 ;
      END
   END dout1[158]
   PIN dout1[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.0025 108.3625 276.1375 108.4975 ;
      END
   END dout1[159]
   PIN dout1[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.1775 108.3625 277.3125 108.4975 ;
      END
   END dout1[160]
   PIN dout1[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.3525 108.3625 278.4875 108.4975 ;
      END
   END dout1[161]
   PIN dout1[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.5275 108.3625 279.6625 108.4975 ;
      END
   END dout1[162]
   PIN dout1[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.7025 108.3625 280.8375 108.4975 ;
      END
   END dout1[163]
   PIN dout1[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.8775 108.3625 282.0125 108.4975 ;
      END
   END dout1[164]
   PIN dout1[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.0525 108.3625 283.1875 108.4975 ;
      END
   END dout1[165]
   PIN dout1[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.2275 108.3625 284.3625 108.4975 ;
      END
   END dout1[166]
   PIN dout1[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.4025 108.3625 285.5375 108.4975 ;
      END
   END dout1[167]
   PIN dout1[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.5775 108.3625 286.7125 108.4975 ;
      END
   END dout1[168]
   PIN dout1[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.7525 108.3625 287.8875 108.4975 ;
      END
   END dout1[169]
   PIN dout1[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.9275 108.3625 289.0625 108.4975 ;
      END
   END dout1[170]
   PIN dout1[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.1025 108.3625 290.2375 108.4975 ;
      END
   END dout1[171]
   PIN dout1[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.2775 108.3625 291.4125 108.4975 ;
      END
   END dout1[172]
   PIN dout1[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.4525 108.3625 292.5875 108.4975 ;
      END
   END dout1[173]
   PIN dout1[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.6275 108.3625 293.7625 108.4975 ;
      END
   END dout1[174]
   PIN dout1[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.8025 108.3625 294.9375 108.4975 ;
      END
   END dout1[175]
   PIN dout1[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.9775 108.3625 296.1125 108.4975 ;
      END
   END dout1[176]
   PIN dout1[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.1525 108.3625 297.2875 108.4975 ;
      END
   END dout1[177]
   PIN dout1[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.3275 108.3625 298.4625 108.4975 ;
      END
   END dout1[178]
   PIN dout1[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.5025 108.3625 299.6375 108.4975 ;
      END
   END dout1[179]
   PIN dout1[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.6775 108.3625 300.8125 108.4975 ;
      END
   END dout1[180]
   PIN dout1[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.8525 108.3625 301.9875 108.4975 ;
      END
   END dout1[181]
   PIN dout1[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.0275 108.3625 303.1625 108.4975 ;
      END
   END dout1[182]
   PIN dout1[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.2025 108.3625 304.3375 108.4975 ;
      END
   END dout1[183]
   PIN dout1[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.3775 108.3625 305.5125 108.4975 ;
      END
   END dout1[184]
   PIN dout1[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.5525 108.3625 306.6875 108.4975 ;
      END
   END dout1[185]
   PIN dout1[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.7275 108.3625 307.8625 108.4975 ;
      END
   END dout1[186]
   PIN dout1[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.9025 108.3625 309.0375 108.4975 ;
      END
   END dout1[187]
   PIN dout1[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.0775 108.3625 310.2125 108.4975 ;
      END
   END dout1[188]
   PIN dout1[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.2525 108.3625 311.3875 108.4975 ;
      END
   END dout1[189]
   PIN dout1[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.4275 108.3625 312.5625 108.4975 ;
      END
   END dout1[190]
   PIN dout1[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.6025 108.3625 313.7375 108.4975 ;
      END
   END dout1[191]
   PIN dout1[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.7775 108.3625 314.9125 108.4975 ;
      END
   END dout1[192]
   PIN dout1[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.9525 108.3625 316.0875 108.4975 ;
      END
   END dout1[193]
   PIN dout1[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.1275 108.3625 317.2625 108.4975 ;
      END
   END dout1[194]
   PIN dout1[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.3025 108.3625 318.4375 108.4975 ;
      END
   END dout1[195]
   PIN dout1[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.4775 108.3625 319.6125 108.4975 ;
      END
   END dout1[196]
   PIN dout1[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.6525 108.3625 320.7875 108.4975 ;
      END
   END dout1[197]
   PIN dout1[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.8275 108.3625 321.9625 108.4975 ;
      END
   END dout1[198]
   PIN dout1[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.0025 108.3625 323.1375 108.4975 ;
      END
   END dout1[199]
   PIN dout1[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.1775 108.3625 324.3125 108.4975 ;
      END
   END dout1[200]
   PIN dout1[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.3525 108.3625 325.4875 108.4975 ;
      END
   END dout1[201]
   PIN dout1[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.5275 108.3625 326.6625 108.4975 ;
      END
   END dout1[202]
   PIN dout1[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.7025 108.3625 327.8375 108.4975 ;
      END
   END dout1[203]
   PIN dout1[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.8775 108.3625 329.0125 108.4975 ;
      END
   END dout1[204]
   PIN dout1[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.0525 108.3625 330.1875 108.4975 ;
      END
   END dout1[205]
   PIN dout1[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.2275 108.3625 331.3625 108.4975 ;
      END
   END dout1[206]
   PIN dout1[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.4025 108.3625 332.5375 108.4975 ;
      END
   END dout1[207]
   PIN dout1[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.5775 108.3625 333.7125 108.4975 ;
      END
   END dout1[208]
   PIN dout1[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.7525 108.3625 334.8875 108.4975 ;
      END
   END dout1[209]
   PIN dout1[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.9275 108.3625 336.0625 108.4975 ;
      END
   END dout1[210]
   PIN dout1[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.1025 108.3625 337.2375 108.4975 ;
      END
   END dout1[211]
   PIN dout1[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.2775 108.3625 338.4125 108.4975 ;
      END
   END dout1[212]
   PIN dout1[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.4525 108.3625 339.5875 108.4975 ;
      END
   END dout1[213]
   PIN dout1[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.6275 108.3625 340.7625 108.4975 ;
      END
   END dout1[214]
   PIN dout1[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.8025 108.3625 341.9375 108.4975 ;
      END
   END dout1[215]
   PIN dout1[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.9775 108.3625 343.1125 108.4975 ;
      END
   END dout1[216]
   PIN dout1[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.1525 108.3625 344.2875 108.4975 ;
      END
   END dout1[217]
   PIN dout1[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.3275 108.3625 345.4625 108.4975 ;
      END
   END dout1[218]
   PIN dout1[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.5025 108.3625 346.6375 108.4975 ;
      END
   END dout1[219]
   PIN dout1[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.6775 108.3625 347.8125 108.4975 ;
      END
   END dout1[220]
   PIN dout1[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.8525 108.3625 348.9875 108.4975 ;
      END
   END dout1[221]
   PIN dout1[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.0275 108.3625 350.1625 108.4975 ;
      END
   END dout1[222]
   PIN dout1[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  351.2025 108.3625 351.3375 108.4975 ;
      END
   END dout1[223]
   PIN dout1[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.3775 108.3625 352.5125 108.4975 ;
      END
   END dout1[224]
   PIN dout1[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.5525 108.3625 353.6875 108.4975 ;
      END
   END dout1[225]
   PIN dout1[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.7275 108.3625 354.8625 108.4975 ;
      END
   END dout1[226]
   PIN dout1[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.9025 108.3625 356.0375 108.4975 ;
      END
   END dout1[227]
   PIN dout1[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.0775 108.3625 357.2125 108.4975 ;
      END
   END dout1[228]
   PIN dout1[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.2525 108.3625 358.3875 108.4975 ;
      END
   END dout1[229]
   PIN dout1[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.4275 108.3625 359.5625 108.4975 ;
      END
   END dout1[230]
   PIN dout1[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.6025 108.3625 360.7375 108.4975 ;
      END
   END dout1[231]
   PIN dout1[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.7775 108.3625 361.9125 108.4975 ;
      END
   END dout1[232]
   PIN dout1[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.9525 108.3625 363.0875 108.4975 ;
      END
   END dout1[233]
   PIN dout1[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.1275 108.3625 364.2625 108.4975 ;
      END
   END dout1[234]
   PIN dout1[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.3025 108.3625 365.4375 108.4975 ;
      END
   END dout1[235]
   PIN dout1[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.4775 108.3625 366.6125 108.4975 ;
      END
   END dout1[236]
   PIN dout1[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.6525 108.3625 367.7875 108.4975 ;
      END
   END dout1[237]
   PIN dout1[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.8275 108.3625 368.9625 108.4975 ;
      END
   END dout1[238]
   PIN dout1[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.0025 108.3625 370.1375 108.4975 ;
      END
   END dout1[239]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  638.3075 2.47 638.4425 2.605 ;
         LAYER metal3 ;
         RECT  523.9075 2.47 524.0425 2.605 ;
         LAYER metal3 ;
         RECT  375.1875 2.47 375.3225 2.605 ;
         LAYER metal4 ;
         RECT  397.17 103.8225 397.31 113.8425 ;
         LAYER metal3 ;
         RECT  558.2275 2.47 558.3625 2.605 ;
         LAYER metal4 ;
         RECT  85.925 47.1425 86.065 101.2125 ;
         LAYER metal3 ;
         RECT  661.1875 2.47 661.3225 2.605 ;
         LAYER metal3 ;
         RECT  478.1475 2.47 478.2825 2.605 ;
         LAYER metal3 ;
         RECT  249.3475 2.47 249.4825 2.605 ;
         LAYER metal3 ;
         RECT  203.5875 2.47 203.7225 2.605 ;
         LAYER metal4 ;
         RECT  84.845 50.3125 84.985 98.2925 ;
         LAYER metal3 ;
         RECT  85.9925 41.0125 370.8075 41.0825 ;
         LAYER metal3 ;
         RECT  66.9675 69.75 67.1025 69.885 ;
         LAYER metal3 ;
         RECT  112.0675 2.47 112.2025 2.605 ;
         LAYER metal3 ;
         RECT  489.5875 2.47 489.7225 2.605 ;
         LAYER metal3 ;
         RECT  695.5075 2.47 695.6425 2.605 ;
         LAYER metal3 ;
         RECT  66.9675 60.78 67.1025 60.915 ;
         LAYER metal3 ;
         RECT  393.3175 63.77 393.4525 63.905 ;
         LAYER metal4 ;
         RECT  72.52 50.3125 72.66 98.3625 ;
         LAYER metal3 ;
         RECT  432.3875 2.47 432.5225 2.605 ;
         LAYER metal3 ;
         RECT  393.3175 66.76 393.4525 66.895 ;
         LAYER metal3 ;
         RECT  317.9875 2.47 318.1225 2.605 ;
         LAYER metal3 ;
         RECT  123.5075 2.47 123.6425 2.605 ;
         LAYER metal3 ;
         RECT  649.7475 2.47 649.8825 2.605 ;
         LAYER metal3 ;
         RECT  684.0675 2.47 684.2025 2.605 ;
         LAYER metal3 ;
         RECT  100.6275 2.47 100.7625 2.605 ;
         LAYER metal3 ;
         RECT  215.0275 2.47 215.1625 2.605 ;
         LAYER metal3 ;
         RECT  420.9475 2.47 421.0825 2.605 ;
         LAYER metal3 ;
         RECT  535.3475 2.47 535.4825 2.605 ;
         LAYER metal3 ;
         RECT  84.8475 48.82 84.9825 48.955 ;
         LAYER metal3 ;
         RECT  386.6275 2.47 386.7625 2.605 ;
         LAYER metal3 ;
         RECT  466.7075 2.47 466.8425 2.605 ;
         LAYER metal3 ;
         RECT  134.9475 2.47 135.0825 2.605 ;
         LAYER metal3 ;
         RECT  77.7475 2.47 77.8825 2.605 ;
         LAYER metal4 ;
         RECT  375.435 50.3125 375.575 98.2925 ;
         LAYER metal3 ;
         RECT  512.4675 2.47 512.6025 2.605 ;
         LAYER metal3 ;
         RECT  392.9725 51.81 393.1075 51.945 ;
         LAYER metal3 ;
         RECT  85.9925 46.4475 371.2775 46.5175 ;
         LAYER metal3 ;
         RECT  672.6275 2.47 672.7625 2.605 ;
         LAYER metal3 ;
         RECT  73.14 49.6075 73.275 49.7425 ;
         LAYER metal3 ;
         RECT  306.5475 2.47 306.6825 2.605 ;
         LAYER metal3 ;
         RECT  443.8275 2.47 443.9625 2.605 ;
         LAYER metal3 ;
         RECT  85.9925 101.9075 372.4525 101.9775 ;
         LAYER metal3 ;
         RECT  226.4675 2.47 226.6025 2.605 ;
         LAYER metal3 ;
         RECT  375.4375 99.65 375.5725 99.785 ;
         LAYER metal3 ;
         RECT  741.2675 2.47 741.4025 2.605 ;
         LAYER metal3 ;
         RECT  352.3075 2.47 352.4425 2.605 ;
         LAYER metal3 ;
         RECT  409.5075 2.47 409.6425 2.605 ;
         LAYER metal3 ;
         RECT  85.9925 105.805 370.8075 105.875 ;
         LAYER metal3 ;
         RECT  272.2275 2.47 272.3625 2.605 ;
         LAYER metal3 ;
         RECT  66.9675 66.76 67.1025 66.895 ;
         LAYER metal4 ;
         RECT  387.76 50.3125 387.9 98.3625 ;
         LAYER metal3 ;
         RECT  392.9725 54.8 393.1075 54.935 ;
         LAYER metal3 ;
         RECT  2.425 32.115 2.56 32.25 ;
         LAYER metal3 ;
         RECT  581.1075 2.47 581.2425 2.605 ;
         LAYER metal4 ;
         RECT  459.9275 84.0625 460.0675 106.465 ;
         LAYER metal3 ;
         RECT  67.3125 54.8 67.4475 54.935 ;
         LAYER metal3 ;
         RECT  66.9675 63.77 67.1025 63.905 ;
         LAYER metal3 ;
         RECT  387.145 98.8625 387.28 98.9975 ;
         LAYER metal3 ;
         RECT  615.4275 2.47 615.5625 2.605 ;
         LAYER metal3 ;
         RECT  329.4275 2.47 329.5625 2.605 ;
         LAYER metal3 ;
         RECT  569.6675 2.47 569.8025 2.605 ;
         LAYER metal3 ;
         RECT  169.2675 2.47 169.4025 2.605 ;
         LAYER metal3 ;
         RECT  157.8275 2.47 157.9625 2.605 ;
         LAYER metal3 ;
         RECT  501.0275 2.47 501.1625 2.605 ;
         LAYER metal3 ;
         RECT  626.8675 2.47 627.0025 2.605 ;
         LAYER metal3 ;
         RECT  67.3125 51.81 67.4475 51.945 ;
         LAYER metal4 ;
         RECT  399.89 37.8975 400.03 50.4525 ;
         LAYER metal3 ;
         RECT  363.7475 2.47 363.8825 2.605 ;
         LAYER metal3 ;
         RECT  393.3175 60.78 393.4525 60.915 ;
         LAYER metal3 ;
         RECT  180.7075 2.47 180.8425 2.605 ;
         LAYER metal4 ;
         RECT  374.355 47.1425 374.495 101.2125 ;
         LAYER metal3 ;
         RECT  146.3875 2.47 146.5225 2.605 ;
         LAYER metal3 ;
         RECT  546.7875 2.47 546.9225 2.605 ;
         LAYER metal3 ;
         RECT  706.9475 2.47 707.0825 2.605 ;
         LAYER metal3 ;
         RECT  192.1475 2.47 192.2825 2.605 ;
         LAYER metal3 ;
         RECT  89.1875 2.47 89.3225 2.605 ;
         LAYER metal3 ;
         RECT  393.3175 69.75 393.4525 69.885 ;
         LAYER metal4 ;
         RECT  60.585 71.2425 60.725 83.7975 ;
         LAYER metal3 ;
         RECT  729.8275 2.47 729.9625 2.605 ;
         LAYER metal3 ;
         RECT  398.0675 2.47 398.2025 2.605 ;
         LAYER metal3 ;
         RECT  295.1075 2.47 295.2425 2.605 ;
         LAYER metal3 ;
         RECT  260.7875 2.47 260.9225 2.605 ;
         LAYER metal3 ;
         RECT  592.5475 2.47 592.6825 2.605 ;
         LAYER metal3 ;
         RECT  458.195 113.705 458.33 113.84 ;
         LAYER metal3 ;
         RECT  66.3075 2.47 66.4425 2.605 ;
         LAYER metal3 ;
         RECT  340.8675 2.47 341.0025 2.605 ;
         LAYER metal3 ;
         RECT  718.3875 2.47 718.5225 2.605 ;
         LAYER metal3 ;
         RECT  237.9075 2.47 238.0425 2.605 ;
         LAYER metal3 ;
         RECT  603.9875 2.47 604.1225 2.605 ;
         LAYER metal3 ;
         RECT  283.6675 2.47 283.8025 2.605 ;
         LAYER metal3 ;
         RECT  455.2675 2.47 455.4025 2.605 ;
         LAYER metal4 ;
         RECT  63.305 32.1125 63.445 47.0725 ;
         LAYER metal4 ;
         RECT  0.6875 39.49 0.8275 61.8925 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  149.2475 0.0 149.3825 0.135 ;
         LAYER metal3 ;
         RECT  469.5675 0.0 469.7025 0.135 ;
         LAYER metal3 ;
         RECT  309.4075 0.0 309.5425 0.135 ;
         LAYER metal3 ;
         RECT  549.6475 0.0 549.7825 0.135 ;
         LAYER metal3 ;
         RECT  378.0475 0.0 378.1825 0.135 ;
         LAYER metal4 ;
         RECT  63.445 71.1775 63.585 83.7325 ;
         LAYER metal4 ;
         RECT  397.03 37.9625 397.17 50.5175 ;
         LAYER metal3 ;
         RECT  641.1675 0.0 641.3025 0.135 ;
         LAYER metal3 ;
         RECT  515.3275 0.0 515.4625 0.135 ;
         LAYER metal3 ;
         RECT  561.0875 0.0 561.2225 0.135 ;
         LAYER metal3 ;
         RECT  458.195 116.175 458.33 116.31 ;
         LAYER metal3 ;
         RECT  160.6875 0.0 160.8225 0.135 ;
         LAYER metal3 ;
         RECT  395.125 59.285 395.26 59.42 ;
         LAYER metal3 ;
         RECT  395.125 62.275 395.26 62.41 ;
         LAYER metal3 ;
         RECT  92.0475 0.0 92.1825 0.135 ;
         LAYER metal3 ;
         RECT  389.4875 0.0 389.6225 0.135 ;
         LAYER metal4 ;
         RECT  86.385 47.1425 86.525 101.2125 ;
         LAYER metal3 ;
         RECT  366.6075 0.0 366.7425 0.135 ;
         LAYER metal3 ;
         RECT  183.5675 0.0 183.7025 0.135 ;
         LAYER metal3 ;
         RECT  252.2075 0.0 252.3425 0.135 ;
         LAYER metal3 ;
         RECT  229.3275 0.0 229.4625 0.135 ;
         LAYER metal3 ;
         RECT  395.125 68.255 395.26 68.39 ;
         LAYER metal4 ;
         RECT  457.865 84.03 458.005 106.4325 ;
         LAYER metal3 ;
         RECT  503.8875 0.0 504.0225 0.135 ;
         LAYER metal3 ;
         RECT  343.7275 0.0 343.8625 0.135 ;
         LAYER metal3 ;
         RECT  65.785 56.295 65.92 56.43 ;
         LAYER metal3 ;
         RECT  395.125 65.265 395.26 65.4 ;
         LAYER metal3 ;
         RECT  583.9675 0.0 584.1025 0.135 ;
         LAYER metal3 ;
         RECT  103.4875 0.0 103.6225 0.135 ;
         LAYER metal3 ;
         RECT  652.6075 0.0 652.7425 0.135 ;
         LAYER metal3 ;
         RECT  394.5 50.315 394.635 50.45 ;
         LAYER metal3 ;
         RECT  618.2875 0.0 618.4225 0.135 ;
         LAYER metal3 ;
         RECT  332.2875 0.0 332.4225 0.135 ;
         LAYER metal3 ;
         RECT  698.3675 0.0 698.5025 0.135 ;
         LAYER metal4 ;
         RECT  2.75 39.5225 2.89 61.925 ;
         LAYER metal3 ;
         RECT  65.16 62.275 65.295 62.41 ;
         LAYER metal3 ;
         RECT  297.9675 0.0 298.1025 0.135 ;
         LAYER metal3 ;
         RECT  744.1275 0.0 744.2625 0.135 ;
         LAYER metal4 ;
         RECT  73.08 50.28 73.22 98.325 ;
         LAYER metal3 ;
         RECT  286.5275 0.0 286.6625 0.135 ;
         LAYER metal3 ;
         RECT  69.1675 0.0 69.3025 0.135 ;
         LAYER metal3 ;
         RECT  85.9925 43.0625 370.8075 43.1325 ;
         LAYER metal3 ;
         RECT  526.7675 0.0 526.9025 0.135 ;
         LAYER metal3 ;
         RECT  423.8075 0.0 423.9425 0.135 ;
         LAYER metal3 ;
         RECT  65.16 71.245 65.295 71.38 ;
         LAYER metal3 ;
         RECT  686.9275 0.0 687.0625 0.135 ;
         LAYER metal3 ;
         RECT  435.2475 0.0 435.3825 0.135 ;
         LAYER metal3 ;
         RECT  263.6475 0.0 263.7825 0.135 ;
         LAYER metal3 ;
         RECT  65.785 50.315 65.92 50.45 ;
         LAYER metal4 ;
         RECT  70.93 50.28 71.07 98.3625 ;
         LAYER metal3 ;
         RECT  412.3675 0.0 412.5025 0.135 ;
         LAYER metal4 ;
         RECT  387.2 50.28 387.34 98.325 ;
         LAYER metal3 ;
         RECT  629.7275 0.0 629.8625 0.135 ;
         LAYER metal3 ;
         RECT  709.8075 0.0 709.9425 0.135 ;
         LAYER metal3 ;
         RECT  400.9275 0.0 401.0625 0.135 ;
         LAYER metal3 ;
         RECT  394.5 56.295 394.635 56.43 ;
         LAYER metal4 ;
         RECT  389.35 50.28 389.49 98.3625 ;
         LAYER metal4 ;
         RECT  6.105 29.6425 6.245 44.6025 ;
         LAYER metal3 ;
         RECT  206.4475 0.0 206.5825 0.135 ;
         LAYER metal3 ;
         RECT  446.6875 0.0 446.8225 0.135 ;
         LAYER metal3 ;
         RECT  492.4475 0.0 492.5825 0.135 ;
         LAYER metal3 ;
         RECT  458.1275 0.0 458.2625 0.135 ;
         LAYER metal3 ;
         RECT  355.1675 0.0 355.3025 0.135 ;
         LAYER metal3 ;
         RECT  275.0875 0.0 275.2225 0.135 ;
         LAYER metal3 ;
         RECT  172.1275 0.0 172.2625 0.135 ;
         LAYER metal3 ;
         RECT  595.4075 0.0 595.5425 0.135 ;
         LAYER metal3 ;
         RECT  675.4875 0.0 675.6225 0.135 ;
         LAYER metal3 ;
         RECT  85.9925 103.9125 370.8425 103.9825 ;
         LAYER metal3 ;
         RECT  195.0075 0.0 195.1425 0.135 ;
         LAYER metal3 ;
         RECT  65.16 65.265 65.295 65.4 ;
         LAYER metal3 ;
         RECT  65.16 59.285 65.295 59.42 ;
         LAYER metal3 ;
         RECT  217.8875 0.0 218.0225 0.135 ;
         LAYER metal3 ;
         RECT  65.16 68.255 65.295 68.39 ;
         LAYER metal3 ;
         RECT  606.8475 0.0 606.9825 0.135 ;
         LAYER metal4 ;
         RECT  454.37 101.3525 454.51 116.3125 ;
         LAYER metal3 ;
         RECT  572.5275 0.0 572.6625 0.135 ;
         LAYER metal3 ;
         RECT  126.3675 0.0 126.5025 0.135 ;
         LAYER metal3 ;
         RECT  664.0475 0.0 664.1825 0.135 ;
         LAYER metal3 ;
         RECT  320.8475 0.0 320.9825 0.135 ;
         LAYER metal3 ;
         RECT  732.6875 0.0 732.8225 0.135 ;
         LAYER metal3 ;
         RECT  80.6075 0.0 80.7425 0.135 ;
         LAYER metal3 ;
         RECT  394.5 53.305 394.635 53.44 ;
         LAYER metal3 ;
         RECT  65.785 53.305 65.92 53.44 ;
         LAYER metal3 ;
         RECT  240.7675 0.0 240.9025 0.135 ;
         LAYER metal3 ;
         RECT  721.2475 0.0 721.3825 0.135 ;
         LAYER metal3 ;
         RECT  395.125 71.245 395.26 71.38 ;
         LAYER metal3 ;
         RECT  137.8075 0.0 137.9425 0.135 ;
         LAYER metal3 ;
         RECT  114.9275 0.0 115.0625 0.135 ;
         LAYER metal3 ;
         RECT  2.425 29.645 2.56 29.78 ;
         LAYER metal3 ;
         RECT  538.2075 0.0 538.3425 0.135 ;
         LAYER metal4 ;
         RECT  373.895 47.1425 374.035 101.2125 ;
         LAYER metal3 ;
         RECT  481.0075 0.0 481.1425 0.135 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 752.635 116.1725 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 752.635 116.1725 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 66.45 0.965 ;
      RECT  0.14 0.965 66.45 1.38 ;
      RECT  66.45 0.14 66.865 0.965 ;
      RECT  66.865 0.965 69.31 1.38 ;
      RECT  69.725 0.965 72.17 1.38 ;
      RECT  72.585 0.965 75.03 1.38 ;
      RECT  75.445 0.965 77.89 1.38 ;
      RECT  78.305 0.965 80.75 1.38 ;
      RECT  81.165 0.965 83.61 1.38 ;
      RECT  84.025 0.965 86.47 1.38 ;
      RECT  86.885 0.965 89.33 1.38 ;
      RECT  89.745 0.965 92.19 1.38 ;
      RECT  92.605 0.965 95.05 1.38 ;
      RECT  95.465 0.965 97.91 1.38 ;
      RECT  98.325 0.965 100.77 1.38 ;
      RECT  101.185 0.965 103.63 1.38 ;
      RECT  104.045 0.965 106.49 1.38 ;
      RECT  106.905 0.965 109.35 1.38 ;
      RECT  109.765 0.965 112.21 1.38 ;
      RECT  112.625 0.965 115.07 1.38 ;
      RECT  115.485 0.965 117.93 1.38 ;
      RECT  118.345 0.965 120.79 1.38 ;
      RECT  121.205 0.965 123.65 1.38 ;
      RECT  124.065 0.965 126.51 1.38 ;
      RECT  126.925 0.965 129.37 1.38 ;
      RECT  129.785 0.965 132.23 1.38 ;
      RECT  132.645 0.965 135.09 1.38 ;
      RECT  135.505 0.965 137.95 1.38 ;
      RECT  138.365 0.965 140.81 1.38 ;
      RECT  141.225 0.965 143.67 1.38 ;
      RECT  144.085 0.965 146.53 1.38 ;
      RECT  146.945 0.965 149.39 1.38 ;
      RECT  149.805 0.965 152.25 1.38 ;
      RECT  152.665 0.965 155.11 1.38 ;
      RECT  155.525 0.965 157.97 1.38 ;
      RECT  158.385 0.965 160.83 1.38 ;
      RECT  161.245 0.965 163.69 1.38 ;
      RECT  164.105 0.965 166.55 1.38 ;
      RECT  166.965 0.965 169.41 1.38 ;
      RECT  169.825 0.965 172.27 1.38 ;
      RECT  172.685 0.965 175.13 1.38 ;
      RECT  175.545 0.965 177.99 1.38 ;
      RECT  178.405 0.965 180.85 1.38 ;
      RECT  181.265 0.965 183.71 1.38 ;
      RECT  184.125 0.965 186.57 1.38 ;
      RECT  186.985 0.965 189.43 1.38 ;
      RECT  189.845 0.965 192.29 1.38 ;
      RECT  192.705 0.965 195.15 1.38 ;
      RECT  195.565 0.965 198.01 1.38 ;
      RECT  198.425 0.965 200.87 1.38 ;
      RECT  201.285 0.965 203.73 1.38 ;
      RECT  204.145 0.965 206.59 1.38 ;
      RECT  207.005 0.965 209.45 1.38 ;
      RECT  209.865 0.965 212.31 1.38 ;
      RECT  212.725 0.965 215.17 1.38 ;
      RECT  215.585 0.965 218.03 1.38 ;
      RECT  218.445 0.965 220.89 1.38 ;
      RECT  221.305 0.965 223.75 1.38 ;
      RECT  224.165 0.965 226.61 1.38 ;
      RECT  227.025 0.965 229.47 1.38 ;
      RECT  229.885 0.965 232.33 1.38 ;
      RECT  232.745 0.965 235.19 1.38 ;
      RECT  235.605 0.965 238.05 1.38 ;
      RECT  238.465 0.965 240.91 1.38 ;
      RECT  241.325 0.965 243.77 1.38 ;
      RECT  244.185 0.965 246.63 1.38 ;
      RECT  247.045 0.965 249.49 1.38 ;
      RECT  249.905 0.965 252.35 1.38 ;
      RECT  252.765 0.965 255.21 1.38 ;
      RECT  255.625 0.965 258.07 1.38 ;
      RECT  258.485 0.965 260.93 1.38 ;
      RECT  261.345 0.965 263.79 1.38 ;
      RECT  264.205 0.965 266.65 1.38 ;
      RECT  267.065 0.965 269.51 1.38 ;
      RECT  269.925 0.965 272.37 1.38 ;
      RECT  272.785 0.965 275.23 1.38 ;
      RECT  275.645 0.965 278.09 1.38 ;
      RECT  278.505 0.965 280.95 1.38 ;
      RECT  281.365 0.965 283.81 1.38 ;
      RECT  284.225 0.965 286.67 1.38 ;
      RECT  287.085 0.965 289.53 1.38 ;
      RECT  289.945 0.965 292.39 1.38 ;
      RECT  292.805 0.965 295.25 1.38 ;
      RECT  295.665 0.965 298.11 1.38 ;
      RECT  298.525 0.965 300.97 1.38 ;
      RECT  301.385 0.965 303.83 1.38 ;
      RECT  304.245 0.965 306.69 1.38 ;
      RECT  307.105 0.965 309.55 1.38 ;
      RECT  309.965 0.965 312.41 1.38 ;
      RECT  312.825 0.965 315.27 1.38 ;
      RECT  315.685 0.965 318.13 1.38 ;
      RECT  318.545 0.965 320.99 1.38 ;
      RECT  321.405 0.965 323.85 1.38 ;
      RECT  324.265 0.965 326.71 1.38 ;
      RECT  327.125 0.965 329.57 1.38 ;
      RECT  329.985 0.965 332.43 1.38 ;
      RECT  332.845 0.965 335.29 1.38 ;
      RECT  335.705 0.965 338.15 1.38 ;
      RECT  338.565 0.965 341.01 1.38 ;
      RECT  341.425 0.965 343.87 1.38 ;
      RECT  344.285 0.965 346.73 1.38 ;
      RECT  347.145 0.965 349.59 1.38 ;
      RECT  350.005 0.965 352.45 1.38 ;
      RECT  352.865 0.965 355.31 1.38 ;
      RECT  355.725 0.965 358.17 1.38 ;
      RECT  358.585 0.965 361.03 1.38 ;
      RECT  361.445 0.965 363.89 1.38 ;
      RECT  364.305 0.965 366.75 1.38 ;
      RECT  367.165 0.965 369.61 1.38 ;
      RECT  370.025 0.965 372.47 1.38 ;
      RECT  372.885 0.965 375.33 1.38 ;
      RECT  375.745 0.965 378.19 1.38 ;
      RECT  378.605 0.965 381.05 1.38 ;
      RECT  381.465 0.965 383.91 1.38 ;
      RECT  384.325 0.965 386.77 1.38 ;
      RECT  387.185 0.965 389.63 1.38 ;
      RECT  390.045 0.965 392.49 1.38 ;
      RECT  392.905 0.965 395.35 1.38 ;
      RECT  395.765 0.965 398.21 1.38 ;
      RECT  398.625 0.965 401.07 1.38 ;
      RECT  401.485 0.965 403.93 1.38 ;
      RECT  404.345 0.965 406.79 1.38 ;
      RECT  407.205 0.965 409.65 1.38 ;
      RECT  410.065 0.965 412.51 1.38 ;
      RECT  412.925 0.965 415.37 1.38 ;
      RECT  415.785 0.965 418.23 1.38 ;
      RECT  418.645 0.965 421.09 1.38 ;
      RECT  421.505 0.965 423.95 1.38 ;
      RECT  424.365 0.965 426.81 1.38 ;
      RECT  427.225 0.965 429.67 1.38 ;
      RECT  430.085 0.965 432.53 1.38 ;
      RECT  432.945 0.965 435.39 1.38 ;
      RECT  435.805 0.965 438.25 1.38 ;
      RECT  438.665 0.965 441.11 1.38 ;
      RECT  441.525 0.965 443.97 1.38 ;
      RECT  444.385 0.965 446.83 1.38 ;
      RECT  447.245 0.965 449.69 1.38 ;
      RECT  450.105 0.965 452.55 1.38 ;
      RECT  452.965 0.965 455.41 1.38 ;
      RECT  455.825 0.965 458.27 1.38 ;
      RECT  458.685 0.965 461.13 1.38 ;
      RECT  461.545 0.965 463.99 1.38 ;
      RECT  464.405 0.965 466.85 1.38 ;
      RECT  467.265 0.965 469.71 1.38 ;
      RECT  470.125 0.965 472.57 1.38 ;
      RECT  472.985 0.965 475.43 1.38 ;
      RECT  475.845 0.965 478.29 1.38 ;
      RECT  478.705 0.965 481.15 1.38 ;
      RECT  481.565 0.965 484.01 1.38 ;
      RECT  484.425 0.965 486.87 1.38 ;
      RECT  487.285 0.965 489.73 1.38 ;
      RECT  490.145 0.965 492.59 1.38 ;
      RECT  493.005 0.965 495.45 1.38 ;
      RECT  495.865 0.965 498.31 1.38 ;
      RECT  498.725 0.965 501.17 1.38 ;
      RECT  501.585 0.965 504.03 1.38 ;
      RECT  504.445 0.965 506.89 1.38 ;
      RECT  507.305 0.965 509.75 1.38 ;
      RECT  510.165 0.965 512.61 1.38 ;
      RECT  513.025 0.965 515.47 1.38 ;
      RECT  515.885 0.965 518.33 1.38 ;
      RECT  518.745 0.965 521.19 1.38 ;
      RECT  521.605 0.965 524.05 1.38 ;
      RECT  524.465 0.965 526.91 1.38 ;
      RECT  527.325 0.965 529.77 1.38 ;
      RECT  530.185 0.965 532.63 1.38 ;
      RECT  533.045 0.965 535.49 1.38 ;
      RECT  535.905 0.965 538.35 1.38 ;
      RECT  538.765 0.965 541.21 1.38 ;
      RECT  541.625 0.965 544.07 1.38 ;
      RECT  544.485 0.965 546.93 1.38 ;
      RECT  547.345 0.965 549.79 1.38 ;
      RECT  550.205 0.965 552.65 1.38 ;
      RECT  553.065 0.965 555.51 1.38 ;
      RECT  555.925 0.965 558.37 1.38 ;
      RECT  558.785 0.965 561.23 1.38 ;
      RECT  561.645 0.965 564.09 1.38 ;
      RECT  564.505 0.965 566.95 1.38 ;
      RECT  567.365 0.965 569.81 1.38 ;
      RECT  570.225 0.965 572.67 1.38 ;
      RECT  573.085 0.965 575.53 1.38 ;
      RECT  575.945 0.965 578.39 1.38 ;
      RECT  578.805 0.965 581.25 1.38 ;
      RECT  581.665 0.965 584.11 1.38 ;
      RECT  584.525 0.965 586.97 1.38 ;
      RECT  587.385 0.965 589.83 1.38 ;
      RECT  590.245 0.965 592.69 1.38 ;
      RECT  593.105 0.965 595.55 1.38 ;
      RECT  595.965 0.965 598.41 1.38 ;
      RECT  598.825 0.965 601.27 1.38 ;
      RECT  601.685 0.965 604.13 1.38 ;
      RECT  604.545 0.965 606.99 1.38 ;
      RECT  607.405 0.965 609.85 1.38 ;
      RECT  610.265 0.965 612.71 1.38 ;
      RECT  613.125 0.965 615.57 1.38 ;
      RECT  615.985 0.965 618.43 1.38 ;
      RECT  618.845 0.965 621.29 1.38 ;
      RECT  621.705 0.965 624.15 1.38 ;
      RECT  624.565 0.965 627.01 1.38 ;
      RECT  627.425 0.965 629.87 1.38 ;
      RECT  630.285 0.965 632.73 1.38 ;
      RECT  633.145 0.965 635.59 1.38 ;
      RECT  636.005 0.965 638.45 1.38 ;
      RECT  638.865 0.965 641.31 1.38 ;
      RECT  641.725 0.965 644.17 1.38 ;
      RECT  644.585 0.965 647.03 1.38 ;
      RECT  647.445 0.965 649.89 1.38 ;
      RECT  650.305 0.965 652.75 1.38 ;
      RECT  653.165 0.965 655.61 1.38 ;
      RECT  656.025 0.965 658.47 1.38 ;
      RECT  658.885 0.965 661.33 1.38 ;
      RECT  661.745 0.965 664.19 1.38 ;
      RECT  664.605 0.965 667.05 1.38 ;
      RECT  667.465 0.965 669.91 1.38 ;
      RECT  670.325 0.965 672.77 1.38 ;
      RECT  673.185 0.965 675.63 1.38 ;
      RECT  676.045 0.965 678.49 1.38 ;
      RECT  678.905 0.965 681.35 1.38 ;
      RECT  681.765 0.965 684.21 1.38 ;
      RECT  684.625 0.965 687.07 1.38 ;
      RECT  687.485 0.965 689.93 1.38 ;
      RECT  690.345 0.965 692.79 1.38 ;
      RECT  693.205 0.965 695.65 1.38 ;
      RECT  696.065 0.965 698.51 1.38 ;
      RECT  698.925 0.965 701.37 1.38 ;
      RECT  701.785 0.965 704.23 1.38 ;
      RECT  704.645 0.965 707.09 1.38 ;
      RECT  707.505 0.965 709.95 1.38 ;
      RECT  710.365 0.965 712.81 1.38 ;
      RECT  713.225 0.965 715.67 1.38 ;
      RECT  716.085 0.965 718.53 1.38 ;
      RECT  718.945 0.965 721.39 1.38 ;
      RECT  721.805 0.965 724.25 1.38 ;
      RECT  724.665 0.965 727.11 1.38 ;
      RECT  727.525 0.965 729.97 1.38 ;
      RECT  730.385 0.965 732.83 1.38 ;
      RECT  733.245 0.965 735.69 1.38 ;
      RECT  736.105 0.965 738.55 1.38 ;
      RECT  738.965 0.965 741.41 1.38 ;
      RECT  741.825 0.965 744.27 1.38 ;
      RECT  744.685 0.965 747.13 1.38 ;
      RECT  747.545 0.965 749.99 1.38 ;
      RECT  750.405 0.965 752.635 1.38 ;
      RECT  0.14 72.21 60.73 72.625 ;
      RECT  0.14 72.625 60.73 116.1725 ;
      RECT  60.73 1.38 61.145 72.21 ;
      RECT  61.145 72.21 66.45 72.625 ;
      RECT  61.145 72.625 66.45 116.1725 ;
      RECT  60.73 72.625 61.145 74.94 ;
      RECT  60.73 75.355 61.145 77.15 ;
      RECT  60.73 77.565 61.145 79.88 ;
      RECT  60.73 80.295 61.145 82.09 ;
      RECT  60.73 82.505 61.145 116.1725 ;
      RECT  399.47 49.485 399.885 116.1725 ;
      RECT  399.885 49.07 752.635 49.485 ;
      RECT  399.47 46.755 399.885 49.07 ;
      RECT  399.47 44.545 399.885 46.34 ;
      RECT  399.47 41.815 399.885 44.13 ;
      RECT  399.47 1.38 399.885 39.19 ;
      RECT  399.47 39.605 399.885 41.4 ;
      RECT  0.14 1.38 0.145 30.61 ;
      RECT  0.14 30.61 0.145 31.025 ;
      RECT  0.14 31.025 0.145 72.21 ;
      RECT  0.145 1.38 0.56 30.61 ;
      RECT  0.145 31.025 0.56 72.21 ;
      RECT  460.195 49.485 460.61 114.93 ;
      RECT  460.195 115.345 460.61 116.1725 ;
      RECT  460.61 49.485 752.635 114.93 ;
      RECT  460.61 114.93 752.635 115.345 ;
      RECT  460.61 115.345 752.635 116.1725 ;
      RECT  0.56 30.61 6.1075 30.695 ;
      RECT  0.56 30.695 6.1075 31.025 ;
      RECT  6.1075 30.61 6.5225 30.695 ;
      RECT  6.5225 30.61 60.73 30.695 ;
      RECT  6.5225 30.695 60.73 31.025 ;
      RECT  0.56 31.025 6.1075 31.11 ;
      RECT  6.1075 31.11 6.5225 72.21 ;
      RECT  6.5225 31.025 60.73 31.11 ;
      RECT  6.5225 31.11 60.73 72.21 ;
      RECT  399.885 49.485 454.0925 114.845 ;
      RECT  399.885 114.845 454.0925 114.93 ;
      RECT  454.0925 49.485 454.5075 114.845 ;
      RECT  454.5075 114.845 460.195 114.93 ;
      RECT  399.885 114.93 454.0925 115.26 ;
      RECT  399.885 115.26 454.0925 115.345 ;
      RECT  454.0925 115.26 454.5075 115.345 ;
      RECT  454.5075 114.93 460.195 115.26 ;
      RECT  454.5075 115.26 460.195 115.345 ;
      RECT  66.865 108.2225 89.0375 108.6375 ;
      RECT  66.865 108.6375 89.0375 116.1725 ;
      RECT  89.0375 108.6375 89.4525 116.1725 ;
      RECT  89.4525 108.6375 399.47 116.1725 ;
      RECT  89.4525 108.2225 90.2125 108.6375 ;
      RECT  90.6275 108.2225 91.3875 108.6375 ;
      RECT  91.8025 108.2225 92.5625 108.6375 ;
      RECT  92.9775 108.2225 93.7375 108.6375 ;
      RECT  94.1525 108.2225 94.9125 108.6375 ;
      RECT  95.3275 108.2225 96.0875 108.6375 ;
      RECT  96.5025 108.2225 97.2625 108.6375 ;
      RECT  97.6775 108.2225 98.4375 108.6375 ;
      RECT  98.8525 108.2225 99.6125 108.6375 ;
      RECT  100.0275 108.2225 100.7875 108.6375 ;
      RECT  101.2025 108.2225 101.9625 108.6375 ;
      RECT  102.3775 108.2225 103.1375 108.6375 ;
      RECT  103.5525 108.2225 104.3125 108.6375 ;
      RECT  104.7275 108.2225 105.4875 108.6375 ;
      RECT  105.9025 108.2225 106.6625 108.6375 ;
      RECT  107.0775 108.2225 107.8375 108.6375 ;
      RECT  108.2525 108.2225 109.0125 108.6375 ;
      RECT  109.4275 108.2225 110.1875 108.6375 ;
      RECT  110.6025 108.2225 111.3625 108.6375 ;
      RECT  111.7775 108.2225 112.5375 108.6375 ;
      RECT  112.9525 108.2225 113.7125 108.6375 ;
      RECT  114.1275 108.2225 114.8875 108.6375 ;
      RECT  115.3025 108.2225 116.0625 108.6375 ;
      RECT  116.4775 108.2225 117.2375 108.6375 ;
      RECT  117.6525 108.2225 118.4125 108.6375 ;
      RECT  118.8275 108.2225 119.5875 108.6375 ;
      RECT  120.0025 108.2225 120.7625 108.6375 ;
      RECT  121.1775 108.2225 121.9375 108.6375 ;
      RECT  122.3525 108.2225 123.1125 108.6375 ;
      RECT  123.5275 108.2225 124.2875 108.6375 ;
      RECT  124.7025 108.2225 125.4625 108.6375 ;
      RECT  125.8775 108.2225 126.6375 108.6375 ;
      RECT  127.0525 108.2225 127.8125 108.6375 ;
      RECT  128.2275 108.2225 128.9875 108.6375 ;
      RECT  129.4025 108.2225 130.1625 108.6375 ;
      RECT  130.5775 108.2225 131.3375 108.6375 ;
      RECT  131.7525 108.2225 132.5125 108.6375 ;
      RECT  132.9275 108.2225 133.6875 108.6375 ;
      RECT  134.1025 108.2225 134.8625 108.6375 ;
      RECT  135.2775 108.2225 136.0375 108.6375 ;
      RECT  136.4525 108.2225 137.2125 108.6375 ;
      RECT  137.6275 108.2225 138.3875 108.6375 ;
      RECT  138.8025 108.2225 139.5625 108.6375 ;
      RECT  139.9775 108.2225 140.7375 108.6375 ;
      RECT  141.1525 108.2225 141.9125 108.6375 ;
      RECT  142.3275 108.2225 143.0875 108.6375 ;
      RECT  143.5025 108.2225 144.2625 108.6375 ;
      RECT  144.6775 108.2225 145.4375 108.6375 ;
      RECT  145.8525 108.2225 146.6125 108.6375 ;
      RECT  147.0275 108.2225 147.7875 108.6375 ;
      RECT  148.2025 108.2225 148.9625 108.6375 ;
      RECT  149.3775 108.2225 150.1375 108.6375 ;
      RECT  150.5525 108.2225 151.3125 108.6375 ;
      RECT  151.7275 108.2225 152.4875 108.6375 ;
      RECT  152.9025 108.2225 153.6625 108.6375 ;
      RECT  154.0775 108.2225 154.8375 108.6375 ;
      RECT  155.2525 108.2225 156.0125 108.6375 ;
      RECT  156.4275 108.2225 157.1875 108.6375 ;
      RECT  157.6025 108.2225 158.3625 108.6375 ;
      RECT  158.7775 108.2225 159.5375 108.6375 ;
      RECT  159.9525 108.2225 160.7125 108.6375 ;
      RECT  161.1275 108.2225 161.8875 108.6375 ;
      RECT  162.3025 108.2225 163.0625 108.6375 ;
      RECT  163.4775 108.2225 164.2375 108.6375 ;
      RECT  164.6525 108.2225 165.4125 108.6375 ;
      RECT  165.8275 108.2225 166.5875 108.6375 ;
      RECT  167.0025 108.2225 167.7625 108.6375 ;
      RECT  168.1775 108.2225 168.9375 108.6375 ;
      RECT  169.3525 108.2225 170.1125 108.6375 ;
      RECT  170.5275 108.2225 171.2875 108.6375 ;
      RECT  171.7025 108.2225 172.4625 108.6375 ;
      RECT  172.8775 108.2225 173.6375 108.6375 ;
      RECT  174.0525 108.2225 174.8125 108.6375 ;
      RECT  175.2275 108.2225 175.9875 108.6375 ;
      RECT  176.4025 108.2225 177.1625 108.6375 ;
      RECT  177.5775 108.2225 178.3375 108.6375 ;
      RECT  178.7525 108.2225 179.5125 108.6375 ;
      RECT  179.9275 108.2225 180.6875 108.6375 ;
      RECT  181.1025 108.2225 181.8625 108.6375 ;
      RECT  182.2775 108.2225 183.0375 108.6375 ;
      RECT  183.4525 108.2225 184.2125 108.6375 ;
      RECT  184.6275 108.2225 185.3875 108.6375 ;
      RECT  185.8025 108.2225 186.5625 108.6375 ;
      RECT  186.9775 108.2225 187.7375 108.6375 ;
      RECT  188.1525 108.2225 188.9125 108.6375 ;
      RECT  189.3275 108.2225 190.0875 108.6375 ;
      RECT  190.5025 108.2225 191.2625 108.6375 ;
      RECT  191.6775 108.2225 192.4375 108.6375 ;
      RECT  192.8525 108.2225 193.6125 108.6375 ;
      RECT  194.0275 108.2225 194.7875 108.6375 ;
      RECT  195.2025 108.2225 195.9625 108.6375 ;
      RECT  196.3775 108.2225 197.1375 108.6375 ;
      RECT  197.5525 108.2225 198.3125 108.6375 ;
      RECT  198.7275 108.2225 199.4875 108.6375 ;
      RECT  199.9025 108.2225 200.6625 108.6375 ;
      RECT  201.0775 108.2225 201.8375 108.6375 ;
      RECT  202.2525 108.2225 203.0125 108.6375 ;
      RECT  203.4275 108.2225 204.1875 108.6375 ;
      RECT  204.6025 108.2225 205.3625 108.6375 ;
      RECT  205.7775 108.2225 206.5375 108.6375 ;
      RECT  206.9525 108.2225 207.7125 108.6375 ;
      RECT  208.1275 108.2225 208.8875 108.6375 ;
      RECT  209.3025 108.2225 210.0625 108.6375 ;
      RECT  210.4775 108.2225 211.2375 108.6375 ;
      RECT  211.6525 108.2225 212.4125 108.6375 ;
      RECT  212.8275 108.2225 213.5875 108.6375 ;
      RECT  214.0025 108.2225 214.7625 108.6375 ;
      RECT  215.1775 108.2225 215.9375 108.6375 ;
      RECT  216.3525 108.2225 217.1125 108.6375 ;
      RECT  217.5275 108.2225 218.2875 108.6375 ;
      RECT  218.7025 108.2225 219.4625 108.6375 ;
      RECT  219.8775 108.2225 220.6375 108.6375 ;
      RECT  221.0525 108.2225 221.8125 108.6375 ;
      RECT  222.2275 108.2225 222.9875 108.6375 ;
      RECT  223.4025 108.2225 224.1625 108.6375 ;
      RECT  224.5775 108.2225 225.3375 108.6375 ;
      RECT  225.7525 108.2225 226.5125 108.6375 ;
      RECT  226.9275 108.2225 227.6875 108.6375 ;
      RECT  228.1025 108.2225 228.8625 108.6375 ;
      RECT  229.2775 108.2225 230.0375 108.6375 ;
      RECT  230.4525 108.2225 231.2125 108.6375 ;
      RECT  231.6275 108.2225 232.3875 108.6375 ;
      RECT  232.8025 108.2225 233.5625 108.6375 ;
      RECT  233.9775 108.2225 234.7375 108.6375 ;
      RECT  235.1525 108.2225 235.9125 108.6375 ;
      RECT  236.3275 108.2225 237.0875 108.6375 ;
      RECT  237.5025 108.2225 238.2625 108.6375 ;
      RECT  238.6775 108.2225 239.4375 108.6375 ;
      RECT  239.8525 108.2225 240.6125 108.6375 ;
      RECT  241.0275 108.2225 241.7875 108.6375 ;
      RECT  242.2025 108.2225 242.9625 108.6375 ;
      RECT  243.3775 108.2225 244.1375 108.6375 ;
      RECT  244.5525 108.2225 245.3125 108.6375 ;
      RECT  245.7275 108.2225 246.4875 108.6375 ;
      RECT  246.9025 108.2225 247.6625 108.6375 ;
      RECT  248.0775 108.2225 248.8375 108.6375 ;
      RECT  249.2525 108.2225 250.0125 108.6375 ;
      RECT  250.4275 108.2225 251.1875 108.6375 ;
      RECT  251.6025 108.2225 252.3625 108.6375 ;
      RECT  252.7775 108.2225 253.5375 108.6375 ;
      RECT  253.9525 108.2225 254.7125 108.6375 ;
      RECT  255.1275 108.2225 255.8875 108.6375 ;
      RECT  256.3025 108.2225 257.0625 108.6375 ;
      RECT  257.4775 108.2225 258.2375 108.6375 ;
      RECT  258.6525 108.2225 259.4125 108.6375 ;
      RECT  259.8275 108.2225 260.5875 108.6375 ;
      RECT  261.0025 108.2225 261.7625 108.6375 ;
      RECT  262.1775 108.2225 262.9375 108.6375 ;
      RECT  263.3525 108.2225 264.1125 108.6375 ;
      RECT  264.5275 108.2225 265.2875 108.6375 ;
      RECT  265.7025 108.2225 266.4625 108.6375 ;
      RECT  266.8775 108.2225 267.6375 108.6375 ;
      RECT  268.0525 108.2225 268.8125 108.6375 ;
      RECT  269.2275 108.2225 269.9875 108.6375 ;
      RECT  270.4025 108.2225 271.1625 108.6375 ;
      RECT  271.5775 108.2225 272.3375 108.6375 ;
      RECT  272.7525 108.2225 273.5125 108.6375 ;
      RECT  273.9275 108.2225 274.6875 108.6375 ;
      RECT  275.1025 108.2225 275.8625 108.6375 ;
      RECT  276.2775 108.2225 277.0375 108.6375 ;
      RECT  277.4525 108.2225 278.2125 108.6375 ;
      RECT  278.6275 108.2225 279.3875 108.6375 ;
      RECT  279.8025 108.2225 280.5625 108.6375 ;
      RECT  280.9775 108.2225 281.7375 108.6375 ;
      RECT  282.1525 108.2225 282.9125 108.6375 ;
      RECT  283.3275 108.2225 284.0875 108.6375 ;
      RECT  284.5025 108.2225 285.2625 108.6375 ;
      RECT  285.6775 108.2225 286.4375 108.6375 ;
      RECT  286.8525 108.2225 287.6125 108.6375 ;
      RECT  288.0275 108.2225 288.7875 108.6375 ;
      RECT  289.2025 108.2225 289.9625 108.6375 ;
      RECT  290.3775 108.2225 291.1375 108.6375 ;
      RECT  291.5525 108.2225 292.3125 108.6375 ;
      RECT  292.7275 108.2225 293.4875 108.6375 ;
      RECT  293.9025 108.2225 294.6625 108.6375 ;
      RECT  295.0775 108.2225 295.8375 108.6375 ;
      RECT  296.2525 108.2225 297.0125 108.6375 ;
      RECT  297.4275 108.2225 298.1875 108.6375 ;
      RECT  298.6025 108.2225 299.3625 108.6375 ;
      RECT  299.7775 108.2225 300.5375 108.6375 ;
      RECT  300.9525 108.2225 301.7125 108.6375 ;
      RECT  302.1275 108.2225 302.8875 108.6375 ;
      RECT  303.3025 108.2225 304.0625 108.6375 ;
      RECT  304.4775 108.2225 305.2375 108.6375 ;
      RECT  305.6525 108.2225 306.4125 108.6375 ;
      RECT  306.8275 108.2225 307.5875 108.6375 ;
      RECT  308.0025 108.2225 308.7625 108.6375 ;
      RECT  309.1775 108.2225 309.9375 108.6375 ;
      RECT  310.3525 108.2225 311.1125 108.6375 ;
      RECT  311.5275 108.2225 312.2875 108.6375 ;
      RECT  312.7025 108.2225 313.4625 108.6375 ;
      RECT  313.8775 108.2225 314.6375 108.6375 ;
      RECT  315.0525 108.2225 315.8125 108.6375 ;
      RECT  316.2275 108.2225 316.9875 108.6375 ;
      RECT  317.4025 108.2225 318.1625 108.6375 ;
      RECT  318.5775 108.2225 319.3375 108.6375 ;
      RECT  319.7525 108.2225 320.5125 108.6375 ;
      RECT  320.9275 108.2225 321.6875 108.6375 ;
      RECT  322.1025 108.2225 322.8625 108.6375 ;
      RECT  323.2775 108.2225 324.0375 108.6375 ;
      RECT  324.4525 108.2225 325.2125 108.6375 ;
      RECT  325.6275 108.2225 326.3875 108.6375 ;
      RECT  326.8025 108.2225 327.5625 108.6375 ;
      RECT  327.9775 108.2225 328.7375 108.6375 ;
      RECT  329.1525 108.2225 329.9125 108.6375 ;
      RECT  330.3275 108.2225 331.0875 108.6375 ;
      RECT  331.5025 108.2225 332.2625 108.6375 ;
      RECT  332.6775 108.2225 333.4375 108.6375 ;
      RECT  333.8525 108.2225 334.6125 108.6375 ;
      RECT  335.0275 108.2225 335.7875 108.6375 ;
      RECT  336.2025 108.2225 336.9625 108.6375 ;
      RECT  337.3775 108.2225 338.1375 108.6375 ;
      RECT  338.5525 108.2225 339.3125 108.6375 ;
      RECT  339.7275 108.2225 340.4875 108.6375 ;
      RECT  340.9025 108.2225 341.6625 108.6375 ;
      RECT  342.0775 108.2225 342.8375 108.6375 ;
      RECT  343.2525 108.2225 344.0125 108.6375 ;
      RECT  344.4275 108.2225 345.1875 108.6375 ;
      RECT  345.6025 108.2225 346.3625 108.6375 ;
      RECT  346.7775 108.2225 347.5375 108.6375 ;
      RECT  347.9525 108.2225 348.7125 108.6375 ;
      RECT  349.1275 108.2225 349.8875 108.6375 ;
      RECT  350.3025 108.2225 351.0625 108.6375 ;
      RECT  351.4775 108.2225 352.2375 108.6375 ;
      RECT  352.6525 108.2225 353.4125 108.6375 ;
      RECT  353.8275 108.2225 354.5875 108.6375 ;
      RECT  355.0025 108.2225 355.7625 108.6375 ;
      RECT  356.1775 108.2225 356.9375 108.6375 ;
      RECT  357.3525 108.2225 358.1125 108.6375 ;
      RECT  358.5275 108.2225 359.2875 108.6375 ;
      RECT  359.7025 108.2225 360.4625 108.6375 ;
      RECT  360.8775 108.2225 361.6375 108.6375 ;
      RECT  362.0525 108.2225 362.8125 108.6375 ;
      RECT  363.2275 108.2225 363.9875 108.6375 ;
      RECT  364.4025 108.2225 365.1625 108.6375 ;
      RECT  365.5775 108.2225 366.3375 108.6375 ;
      RECT  366.7525 108.2225 367.5125 108.6375 ;
      RECT  367.9275 108.2225 368.6875 108.6375 ;
      RECT  369.1025 108.2225 369.8625 108.6375 ;
      RECT  370.2775 108.2225 399.47 108.6375 ;
      RECT  399.885 1.38 638.1675 2.33 ;
      RECT  399.885 2.745 638.1675 49.07 ;
      RECT  638.1675 1.38 638.5825 2.33 ;
      RECT  638.1675 2.745 638.5825 49.07 ;
      RECT  638.5825 1.38 752.635 2.33 ;
      RECT  638.5825 2.745 752.635 49.07 ;
      RECT  66.865 1.38 375.0475 2.33 ;
      RECT  375.0475 1.38 375.4625 2.33 ;
      RECT  375.0475 2.745 375.4625 49.07 ;
      RECT  375.4625 1.38 399.47 2.33 ;
      RECT  375.4625 2.745 399.47 49.07 ;
      RECT  66.865 2.745 85.8525 40.8725 ;
      RECT  66.865 40.8725 85.8525 41.2225 ;
      RECT  85.8525 2.745 370.9475 40.8725 ;
      RECT  370.9475 2.745 375.0475 40.8725 ;
      RECT  370.9475 40.8725 375.0475 41.2225 ;
      RECT  66.45 69.61 66.8275 70.025 ;
      RECT  66.45 70.025 66.8275 116.1725 ;
      RECT  66.8275 70.025 66.865 116.1725 ;
      RECT  66.865 70.025 67.2425 108.2225 ;
      RECT  67.2425 69.61 89.0375 70.025 ;
      RECT  478.4225 2.33 489.4475 2.745 ;
      RECT  66.8275 1.38 66.865 60.64 ;
      RECT  89.4525 63.63 393.1775 64.045 ;
      RECT  393.5925 63.63 399.47 64.045 ;
      RECT  393.1775 64.045 393.5925 66.62 ;
      RECT  112.3425 2.33 123.3675 2.745 ;
      RECT  638.5825 2.33 649.6075 2.745 ;
      RECT  650.0225 2.33 661.0475 2.745 ;
      RECT  684.3425 2.33 695.3675 2.745 ;
      RECT  100.9025 2.33 111.9275 2.745 ;
      RECT  203.8625 2.33 214.8875 2.745 ;
      RECT  421.2225 2.33 432.2475 2.745 ;
      RECT  524.1825 2.33 535.2075 2.745 ;
      RECT  66.865 49.07 84.7075 49.095 ;
      RECT  84.7075 49.095 85.1225 49.485 ;
      RECT  85.1225 49.07 399.47 49.095 ;
      RECT  85.1225 49.095 399.47 49.485 ;
      RECT  66.865 41.2225 84.7075 48.68 ;
      RECT  66.865 48.68 84.7075 49.07 ;
      RECT  84.7075 41.2225 85.1225 48.68 ;
      RECT  85.1225 41.2225 85.8525 48.68 ;
      RECT  85.1225 48.68 85.8525 49.07 ;
      RECT  375.4625 2.33 386.4875 2.745 ;
      RECT  466.9825 2.33 478.0075 2.745 ;
      RECT  123.7825 2.33 134.8075 2.745 ;
      RECT  66.865 2.33 77.6075 2.745 ;
      RECT  512.7425 2.33 523.7675 2.745 ;
      RECT  89.4525 49.485 392.8325 51.67 ;
      RECT  89.4525 51.67 392.8325 52.085 ;
      RECT  89.4525 52.085 392.8325 63.63 ;
      RECT  392.8325 49.485 393.1775 51.67 ;
      RECT  393.1775 49.485 393.2475 51.67 ;
      RECT  393.2475 49.485 393.5925 51.67 ;
      RECT  393.2475 51.67 393.5925 52.085 ;
      RECT  85.8525 46.6575 370.9475 49.07 ;
      RECT  370.9475 41.2225 371.4175 46.3075 ;
      RECT  370.9475 46.6575 371.4175 49.07 ;
      RECT  371.4175 41.2225 375.0475 46.3075 ;
      RECT  371.4175 46.3075 375.0475 46.6575 ;
      RECT  371.4175 46.6575 375.0475 49.07 ;
      RECT  661.4625 2.33 672.4875 2.745 ;
      RECT  672.9025 2.33 683.9275 2.745 ;
      RECT  67.2425 49.485 73.0 49.8825 ;
      RECT  73.0 49.8825 73.415 69.61 ;
      RECT  73.415 49.485 89.0375 49.8825 ;
      RECT  73.415 49.8825 89.0375 69.61 ;
      RECT  66.865 49.095 73.0 49.4675 ;
      RECT  66.865 49.4675 73.0 49.485 ;
      RECT  73.0 49.095 73.415 49.4675 ;
      RECT  73.415 49.095 84.7075 49.4675 ;
      RECT  73.415 49.4675 84.7075 49.485 ;
      RECT  306.8225 2.33 317.8475 2.745 ;
      RECT  432.6625 2.33 443.6875 2.745 ;
      RECT  89.0375 49.485 89.4525 101.7675 ;
      RECT  67.2425 70.025 85.8525 101.7675 ;
      RECT  67.2425 101.7675 85.8525 102.1175 ;
      RECT  67.2425 102.1175 85.8525 108.2225 ;
      RECT  85.8525 70.025 89.0375 101.7675 ;
      RECT  89.4525 64.045 372.5925 101.7675 ;
      RECT  372.5925 101.7675 393.1775 102.1175 ;
      RECT  372.5925 102.1175 393.1775 108.2225 ;
      RECT  215.3025 2.33 226.3275 2.745 ;
      RECT  372.5925 64.045 375.2975 99.51 ;
      RECT  372.5925 99.51 375.2975 99.925 ;
      RECT  372.5925 99.925 375.2975 101.7675 ;
      RECT  375.2975 64.045 375.7125 99.51 ;
      RECT  375.2975 99.925 375.7125 101.7675 ;
      RECT  375.7125 99.51 393.1775 99.925 ;
      RECT  375.7125 99.925 393.1775 101.7675 ;
      RECT  741.5425 2.33 752.635 2.745 ;
      RECT  399.885 2.33 409.3675 2.745 ;
      RECT  409.7825 2.33 420.8075 2.745 ;
      RECT  89.0375 106.015 89.4525 108.2225 ;
      RECT  85.8525 106.015 89.0375 108.2225 ;
      RECT  89.4525 106.015 370.9475 108.2225 ;
      RECT  370.9475 105.665 372.5925 106.015 ;
      RECT  370.9475 106.015 372.5925 108.2225 ;
      RECT  66.8275 67.035 66.865 69.61 ;
      RECT  66.865 67.035 67.2425 69.61 ;
      RECT  392.8325 52.085 393.1775 54.66 ;
      RECT  392.8325 55.075 393.1775 63.63 ;
      RECT  393.1775 52.085 393.2475 54.66 ;
      RECT  0.56 31.11 2.285 31.975 ;
      RECT  0.56 31.975 2.285 32.39 ;
      RECT  0.56 32.39 2.285 72.21 ;
      RECT  2.285 31.11 2.7 31.975 ;
      RECT  2.285 32.39 2.7 72.21 ;
      RECT  2.7 31.11 6.1075 31.975 ;
      RECT  2.7 31.975 6.1075 32.39 ;
      RECT  2.7 32.39 6.1075 72.21 ;
      RECT  66.865 49.485 67.1725 54.66 ;
      RECT  66.865 54.66 67.1725 55.075 ;
      RECT  66.865 55.075 67.1725 60.64 ;
      RECT  67.1725 55.075 67.2425 60.64 ;
      RECT  67.2425 55.075 67.5875 69.61 ;
      RECT  67.5875 49.8825 73.0 54.66 ;
      RECT  67.5875 54.66 73.0 55.075 ;
      RECT  67.5875 55.075 73.0 69.61 ;
      RECT  66.8275 61.055 66.865 63.63 ;
      RECT  66.8275 64.045 66.865 66.62 ;
      RECT  66.865 61.055 67.2425 63.63 ;
      RECT  66.865 64.045 67.2425 66.62 ;
      RECT  375.7125 64.045 387.005 98.7225 ;
      RECT  375.7125 98.7225 387.005 99.1375 ;
      RECT  375.7125 99.1375 387.005 99.51 ;
      RECT  387.005 64.045 387.42 98.7225 ;
      RECT  387.005 99.1375 387.42 99.51 ;
      RECT  387.42 64.045 393.1775 98.7225 ;
      RECT  387.42 98.7225 393.1775 99.1375 ;
      RECT  387.42 99.1375 393.1775 99.51 ;
      RECT  318.2625 2.33 329.2875 2.745 ;
      RECT  558.5025 2.33 569.5275 2.745 ;
      RECT  569.9425 2.33 580.9675 2.745 ;
      RECT  158.1025 2.33 169.1275 2.745 ;
      RECT  489.8625 2.33 500.8875 2.745 ;
      RECT  501.3025 2.33 512.3275 2.745 ;
      RECT  615.7025 2.33 626.7275 2.745 ;
      RECT  627.1425 2.33 638.1675 2.745 ;
      RECT  67.1725 49.485 67.2425 51.67 ;
      RECT  67.1725 52.085 67.2425 54.66 ;
      RECT  67.2425 49.8825 67.5875 51.67 ;
      RECT  67.2425 52.085 67.5875 54.66 ;
      RECT  352.5825 2.33 363.6075 2.745 ;
      RECT  364.0225 2.33 375.0475 2.745 ;
      RECT  393.2475 52.085 393.5925 60.64 ;
      RECT  393.2475 61.055 393.5925 63.63 ;
      RECT  393.1775 55.075 393.2475 60.64 ;
      RECT  393.1775 61.055 393.2475 63.63 ;
      RECT  169.5425 2.33 180.5675 2.745 ;
      RECT  135.2225 2.33 146.2475 2.745 ;
      RECT  146.6625 2.33 157.6875 2.745 ;
      RECT  535.6225 2.33 546.6475 2.745 ;
      RECT  547.0625 2.33 558.0875 2.745 ;
      RECT  695.7825 2.33 706.8075 2.745 ;
      RECT  180.9825 2.33 192.0075 2.745 ;
      RECT  192.4225 2.33 203.4475 2.745 ;
      RECT  78.0225 2.33 89.0475 2.745 ;
      RECT  89.4625 2.33 100.4875 2.745 ;
      RECT  393.1775 67.035 393.5925 69.61 ;
      RECT  393.1775 70.025 393.5925 108.2225 ;
      RECT  730.1025 2.33 741.1275 2.745 ;
      RECT  386.9025 2.33 397.9275 2.745 ;
      RECT  398.3425 2.33 399.47 2.745 ;
      RECT  295.3825 2.33 306.4075 2.745 ;
      RECT  249.6225 2.33 260.6475 2.745 ;
      RECT  261.0625 2.33 272.0875 2.745 ;
      RECT  581.3825 2.33 592.4075 2.745 ;
      RECT  454.5075 49.485 458.055 113.565 ;
      RECT  454.5075 113.565 458.055 113.98 ;
      RECT  454.5075 113.98 458.055 114.845 ;
      RECT  458.055 49.485 458.47 113.565 ;
      RECT  458.055 113.98 458.47 114.845 ;
      RECT  458.47 49.485 460.195 113.565 ;
      RECT  458.47 113.565 460.195 113.98 ;
      RECT  458.47 113.98 460.195 114.845 ;
      RECT  61.145 1.38 66.1675 2.33 ;
      RECT  61.145 2.33 66.1675 2.745 ;
      RECT  66.1675 1.38 66.45 2.33 ;
      RECT  66.1675 2.745 66.45 72.21 ;
      RECT  66.45 1.38 66.5825 2.33 ;
      RECT  66.45 2.745 66.5825 69.61 ;
      RECT  66.5825 1.38 66.8275 2.33 ;
      RECT  66.5825 2.33 66.8275 2.745 ;
      RECT  66.5825 2.745 66.8275 69.61 ;
      RECT  329.7025 2.33 340.7275 2.745 ;
      RECT  341.1425 2.33 352.1675 2.745 ;
      RECT  707.2225 2.33 718.2475 2.745 ;
      RECT  718.6625 2.33 729.6875 2.745 ;
      RECT  226.7425 2.33 237.7675 2.745 ;
      RECT  238.1825 2.33 249.2075 2.745 ;
      RECT  592.8225 2.33 603.8475 2.745 ;
      RECT  604.2625 2.33 615.2875 2.745 ;
      RECT  272.5025 2.33 283.5275 2.745 ;
      RECT  283.9425 2.33 294.9675 2.745 ;
      RECT  444.1025 2.33 455.1275 2.745 ;
      RECT  455.5425 2.33 466.5675 2.745 ;
      RECT  66.865 0.275 149.1075 0.965 ;
      RECT  149.1075 0.275 149.5225 0.965 ;
      RECT  149.5225 0.275 752.635 0.965 ;
      RECT  549.9225 0.14 560.9475 0.275 ;
      RECT  399.885 115.345 458.055 116.035 ;
      RECT  399.885 116.035 458.055 116.1725 ;
      RECT  458.055 115.345 458.47 116.035 ;
      RECT  458.47 115.345 460.195 116.035 ;
      RECT  458.47 116.035 460.195 116.1725 ;
      RECT  149.5225 0.14 160.5475 0.275 ;
      RECT  393.5925 59.145 394.985 59.56 ;
      RECT  393.5925 59.56 394.985 63.63 ;
      RECT  394.985 49.485 395.4 59.145 ;
      RECT  395.4 49.485 399.47 59.145 ;
      RECT  395.4 59.145 399.47 59.56 ;
      RECT  395.4 59.56 399.47 63.63 ;
      RECT  394.985 59.56 395.4 62.135 ;
      RECT  394.985 62.55 395.4 63.63 ;
      RECT  378.3225 0.14 389.3475 0.275 ;
      RECT  366.8825 0.14 377.9075 0.275 ;
      RECT  393.5925 64.045 394.985 68.115 ;
      RECT  393.5925 68.115 394.985 68.53 ;
      RECT  393.5925 68.53 394.985 108.2225 ;
      RECT  395.4 64.045 399.47 68.115 ;
      RECT  395.4 68.115 399.47 68.53 ;
      RECT  395.4 68.53 399.47 108.2225 ;
      RECT  504.1625 0.14 515.1875 0.275 ;
      RECT  61.145 2.745 65.645 56.155 ;
      RECT  61.145 56.155 65.645 56.57 ;
      RECT  65.645 56.57 66.06 72.21 ;
      RECT  66.06 2.745 66.1675 56.155 ;
      RECT  66.06 56.155 66.1675 56.57 ;
      RECT  66.06 56.57 66.1675 72.21 ;
      RECT  394.985 64.045 395.4 65.125 ;
      RECT  394.985 65.54 395.4 68.115 ;
      RECT  92.3225 0.14 103.3475 0.275 ;
      RECT  641.4425 0.14 652.4675 0.275 ;
      RECT  393.5925 49.485 394.36 50.175 ;
      RECT  393.5925 50.175 394.36 50.59 ;
      RECT  393.5925 50.59 394.36 59.145 ;
      RECT  394.36 49.485 394.775 50.175 ;
      RECT  394.775 49.485 394.985 50.175 ;
      RECT  394.775 50.175 394.985 50.59 ;
      RECT  394.775 50.59 394.985 59.145 ;
      RECT  332.5625 0.14 343.5875 0.275 ;
      RECT  61.145 56.57 65.02 62.135 ;
      RECT  61.145 62.135 65.02 62.55 ;
      RECT  61.145 62.55 65.02 72.21 ;
      RECT  65.435 56.57 65.645 62.135 ;
      RECT  65.435 62.135 65.645 62.55 ;
      RECT  65.435 62.55 65.645 72.21 ;
      RECT  298.2425 0.14 309.2675 0.275 ;
      RECT  744.4025 0.14 752.635 0.275 ;
      RECT  286.8025 0.14 297.8275 0.275 ;
      RECT  66.865 0.14 69.0275 0.275 ;
      RECT  85.8525 41.2225 370.9475 42.9225 ;
      RECT  85.8525 43.2725 370.9475 46.3075 ;
      RECT  515.6025 0.14 526.6275 0.275 ;
      RECT  65.02 71.52 65.435 72.21 ;
      RECT  687.2025 0.14 698.2275 0.275 ;
      RECT  424.0825 0.14 435.1075 0.275 ;
      RECT  252.4825 0.14 263.5075 0.275 ;
      RECT  65.645 2.745 66.06 50.175 ;
      RECT  412.6425 0.14 423.6675 0.275 ;
      RECT  618.5625 0.14 629.5875 0.275 ;
      RECT  630.0025 0.14 641.0275 0.275 ;
      RECT  698.6425 0.14 709.6675 0.275 ;
      RECT  389.7625 0.14 400.7875 0.275 ;
      RECT  401.2025 0.14 412.2275 0.275 ;
      RECT  394.36 56.57 394.775 59.145 ;
      RECT  435.5225 0.14 446.5475 0.275 ;
      RECT  492.7225 0.14 503.7475 0.275 ;
      RECT  446.9625 0.14 457.9875 0.275 ;
      RECT  458.4025 0.14 469.4275 0.275 ;
      RECT  344.0025 0.14 355.0275 0.275 ;
      RECT  355.4425 0.14 366.4675 0.275 ;
      RECT  263.9225 0.14 274.9475 0.275 ;
      RECT  275.3625 0.14 286.3875 0.275 ;
      RECT  160.9625 0.14 171.9875 0.275 ;
      RECT  172.4025 0.14 183.4275 0.275 ;
      RECT  584.2425 0.14 595.2675 0.275 ;
      RECT  675.7625 0.14 686.7875 0.275 ;
      RECT  89.0375 102.1175 89.4525 103.7725 ;
      RECT  89.0375 104.1225 89.4525 105.665 ;
      RECT  85.8525 102.1175 89.0375 103.7725 ;
      RECT  85.8525 104.1225 89.0375 105.665 ;
      RECT  89.4525 102.1175 370.9475 103.7725 ;
      RECT  89.4525 104.1225 370.9475 105.665 ;
      RECT  370.9475 102.1175 370.9825 103.7725 ;
      RECT  370.9475 104.1225 370.9825 105.665 ;
      RECT  370.9825 102.1175 372.5925 103.7725 ;
      RECT  370.9825 103.7725 372.5925 104.1225 ;
      RECT  370.9825 104.1225 372.5925 105.665 ;
      RECT  183.8425 0.14 194.8675 0.275 ;
      RECT  195.2825 0.14 206.3075 0.275 ;
      RECT  65.02 62.55 65.435 65.125 ;
      RECT  65.02 56.57 65.435 59.145 ;
      RECT  65.02 59.56 65.435 62.135 ;
      RECT  206.7225 0.14 217.7475 0.275 ;
      RECT  218.1625 0.14 229.1875 0.275 ;
      RECT  65.02 65.54 65.435 68.115 ;
      RECT  65.02 68.53 65.435 71.105 ;
      RECT  595.6825 0.14 606.7075 0.275 ;
      RECT  607.1225 0.14 618.1475 0.275 ;
      RECT  561.3625 0.14 572.3875 0.275 ;
      RECT  572.8025 0.14 583.8275 0.275 ;
      RECT  652.8825 0.14 663.9075 0.275 ;
      RECT  664.3225 0.14 675.3475 0.275 ;
      RECT  309.6825 0.14 320.7075 0.275 ;
      RECT  321.1225 0.14 332.1475 0.275 ;
      RECT  732.9625 0.14 743.9875 0.275 ;
      RECT  69.4425 0.14 80.4675 0.275 ;
      RECT  80.8825 0.14 91.9075 0.275 ;
      RECT  394.36 50.59 394.775 53.165 ;
      RECT  394.36 53.58 394.775 56.155 ;
      RECT  65.645 50.59 66.06 53.165 ;
      RECT  65.645 53.58 66.06 56.155 ;
      RECT  229.6025 0.14 240.6275 0.275 ;
      RECT  241.0425 0.14 252.0675 0.275 ;
      RECT  710.0825 0.14 721.1075 0.275 ;
      RECT  721.5225 0.14 732.5475 0.275 ;
      RECT  394.985 68.53 395.4 71.105 ;
      RECT  394.985 71.52 395.4 108.2225 ;
      RECT  126.6425 0.14 137.6675 0.275 ;
      RECT  138.0825 0.14 149.1075 0.275 ;
      RECT  103.7625 0.14 114.7875 0.275 ;
      RECT  115.2025 0.14 126.2275 0.275 ;
      RECT  0.56 1.38 2.285 29.505 ;
      RECT  0.56 29.505 2.285 29.92 ;
      RECT  0.56 29.92 2.285 30.61 ;
      RECT  2.285 1.38 2.7 29.505 ;
      RECT  2.285 29.92 2.7 30.61 ;
      RECT  2.7 1.38 60.73 29.505 ;
      RECT  2.7 29.505 60.73 29.92 ;
      RECT  2.7 29.92 60.73 30.61 ;
      RECT  527.0425 0.14 538.0675 0.275 ;
      RECT  538.4825 0.14 549.5075 0.275 ;
      RECT  469.8425 0.14 480.8675 0.275 ;
      RECT  481.2825 0.14 492.3075 0.275 ;
   LAYER  metal4 ;
      RECT  0.14 103.5425 396.89 114.1225 ;
      RECT  0.14 114.1225 396.89 116.1725 ;
      RECT  396.89 114.1225 397.59 116.1725 ;
      RECT  0.14 101.4925 85.645 103.5425 ;
      RECT  85.645 0.14 86.345 46.8625 ;
      RECT  85.645 101.4925 86.345 103.5425 ;
      RECT  86.345 101.4925 396.89 103.5425 ;
      RECT  84.565 46.8625 85.265 50.0325 ;
      RECT  84.565 98.5725 85.265 101.4925 ;
      RECT  85.265 46.8625 85.645 50.0325 ;
      RECT  85.265 50.0325 85.645 98.5725 ;
      RECT  85.265 98.5725 85.645 101.4925 ;
      RECT  0.14 98.6425 72.24 101.4925 ;
      RECT  72.24 98.6425 72.94 101.4925 ;
      RECT  72.94 98.6425 84.565 101.4925 ;
      RECT  375.155 46.8625 375.855 50.0325 ;
      RECT  375.155 98.5725 375.855 101.4925 ;
      RECT  375.855 98.6425 387.48 101.4925 ;
      RECT  387.48 98.6425 388.18 101.4925 ;
      RECT  388.18 98.6425 396.89 101.4925 ;
      RECT  459.6475 0.14 460.3475 83.7825 ;
      RECT  460.3475 0.14 752.635 83.7825 ;
      RECT  460.3475 83.7825 752.635 103.5425 ;
      RECT  459.6475 106.745 460.3475 114.1225 ;
      RECT  460.3475 103.5425 752.635 106.745 ;
      RECT  460.3475 106.745 752.635 114.1225 ;
      RECT  397.59 0.14 399.61 37.6175 ;
      RECT  397.59 37.6175 399.61 50.7325 ;
      RECT  397.59 50.7325 399.61 83.7825 ;
      RECT  399.61 0.14 400.31 37.6175 ;
      RECT  399.61 50.7325 400.31 83.7825 ;
      RECT  400.31 0.14 459.6475 37.6175 ;
      RECT  400.31 37.6175 459.6475 50.7325 ;
      RECT  374.775 46.8625 375.155 50.0325 ;
      RECT  374.775 50.0325 375.155 98.5725 ;
      RECT  374.775 98.5725 375.155 101.4925 ;
      RECT  0.14 70.9625 60.305 84.0775 ;
      RECT  0.14 84.0775 60.305 98.5725 ;
      RECT  60.305 50.0325 61.005 70.9625 ;
      RECT  60.305 84.0775 61.005 98.5725 ;
      RECT  63.025 0.14 63.725 31.8325 ;
      RECT  63.725 0.14 85.645 31.8325 ;
      RECT  63.725 31.8325 85.645 46.8625 ;
      RECT  63.025 47.3525 63.725 50.0325 ;
      RECT  63.725 46.8625 84.565 47.3525 ;
      RECT  0.14 50.0325 0.4075 62.1725 ;
      RECT  0.14 62.1725 0.4075 70.9625 ;
      RECT  0.4075 62.1725 1.1075 70.9625 ;
      RECT  0.14 31.8325 0.4075 39.21 ;
      RECT  0.14 39.21 0.4075 46.8625 ;
      RECT  0.4075 31.8325 1.1075 39.21 ;
      RECT  0.14 46.8625 0.4075 47.3525 ;
      RECT  0.14 47.3525 0.4075 50.0325 ;
      RECT  61.005 50.0325 63.165 70.8975 ;
      RECT  61.005 70.8975 63.165 70.9625 ;
      RECT  63.165 50.0325 63.865 70.8975 ;
      RECT  61.005 70.9625 63.165 84.0125 ;
      RECT  61.005 84.0125 63.165 84.0775 ;
      RECT  63.165 84.0125 63.865 84.0775 ;
      RECT  396.89 0.14 397.45 37.6825 ;
      RECT  396.89 50.7975 397.45 103.5425 ;
      RECT  397.45 0.14 397.59 37.6825 ;
      RECT  397.45 37.6825 397.59 50.7975 ;
      RECT  397.45 50.7975 397.59 103.5425 ;
      RECT  86.345 0.14 396.75 37.6825 ;
      RECT  86.345 37.6825 396.75 46.8625 ;
      RECT  396.75 0.14 396.89 37.6825 ;
      RECT  396.75 50.7975 396.89 98.5725 ;
      RECT  458.285 83.7825 459.6475 103.5425 ;
      RECT  457.585 106.7125 458.285 106.745 ;
      RECT  458.285 103.5425 459.6475 106.7125 ;
      RECT  458.285 106.7125 459.6475 106.745 ;
      RECT  400.31 50.7325 457.585 83.75 ;
      RECT  400.31 83.75 457.585 83.7825 ;
      RECT  457.585 50.7325 458.285 83.75 ;
      RECT  458.285 50.7325 459.6475 83.75 ;
      RECT  458.285 83.75 459.6475 83.7825 ;
      RECT  1.1075 50.0325 2.47 62.1725 ;
      RECT  3.17 50.0325 60.305 62.1725 ;
      RECT  1.1075 62.1725 2.47 62.205 ;
      RECT  1.1075 62.205 2.47 70.9625 ;
      RECT  2.47 62.205 3.17 70.9625 ;
      RECT  3.17 62.1725 60.305 62.205 ;
      RECT  3.17 62.205 60.305 70.9625 ;
      RECT  1.1075 39.21 2.47 39.2425 ;
      RECT  1.1075 39.2425 2.47 46.8625 ;
      RECT  2.47 39.21 3.17 39.2425 ;
      RECT  1.1075 46.8625 2.47 47.3525 ;
      RECT  3.17 46.8625 63.025 47.3525 ;
      RECT  1.1075 47.3525 2.47 50.0325 ;
      RECT  3.17 47.3525 63.025 50.0325 ;
      RECT  73.5 50.0325 84.565 98.5725 ;
      RECT  72.94 98.605 73.5 98.6425 ;
      RECT  73.5 98.5725 84.565 98.605 ;
      RECT  73.5 98.605 84.565 98.6425 ;
      RECT  63.725 47.3525 72.8 50.0 ;
      RECT  72.8 47.3525 73.5 50.0 ;
      RECT  73.5 47.3525 84.565 50.0 ;
      RECT  73.5 50.0 84.565 50.0325 ;
      RECT  0.14 98.5725 70.65 98.6425 ;
      RECT  71.35 98.5725 72.24 98.6425 ;
      RECT  61.005 84.0775 70.65 98.5725 ;
      RECT  71.35 84.0775 72.24 98.5725 ;
      RECT  63.865 50.0325 70.65 70.8975 ;
      RECT  71.35 50.0325 72.24 70.8975 ;
      RECT  63.865 70.8975 70.65 70.9625 ;
      RECT  71.35 70.8975 72.24 70.9625 ;
      RECT  63.865 70.9625 70.65 84.0125 ;
      RECT  71.35 70.9625 72.24 84.0125 ;
      RECT  63.865 84.0125 70.65 84.0775 ;
      RECT  71.35 84.0125 72.24 84.0775 ;
      RECT  63.725 50.0 70.65 50.0325 ;
      RECT  71.35 50.0 72.8 50.0325 ;
      RECT  375.855 50.0325 386.92 98.5725 ;
      RECT  375.855 98.5725 386.92 98.605 ;
      RECT  375.855 98.605 386.92 98.6425 ;
      RECT  386.92 98.605 387.48 98.6425 ;
      RECT  375.855 46.8625 386.92 50.0 ;
      RECT  375.855 50.0 386.92 50.0325 ;
      RECT  386.92 46.8625 387.62 50.0 ;
      RECT  387.62 46.8625 396.75 50.0 ;
      RECT  388.18 98.5725 389.07 98.6425 ;
      RECT  389.77 98.5725 396.89 98.6425 ;
      RECT  388.18 50.0325 389.07 50.7975 ;
      RECT  389.77 50.0325 396.75 50.7975 ;
      RECT  388.18 50.7975 389.07 98.5725 ;
      RECT  389.77 50.7975 396.75 98.5725 ;
      RECT  387.62 50.0 389.07 50.0325 ;
      RECT  389.77 50.0 396.75 50.0325 ;
      RECT  0.14 0.14 5.825 29.3625 ;
      RECT  0.14 29.3625 5.825 31.8325 ;
      RECT  5.825 0.14 6.525 29.3625 ;
      RECT  6.525 0.14 63.025 29.3625 ;
      RECT  6.525 29.3625 63.025 31.8325 ;
      RECT  1.1075 31.8325 5.825 39.21 ;
      RECT  6.525 31.8325 63.025 39.21 ;
      RECT  3.17 39.21 5.825 39.2425 ;
      RECT  6.525 39.21 63.025 39.2425 ;
      RECT  3.17 39.2425 5.825 44.8825 ;
      RECT  3.17 44.8825 5.825 46.8625 ;
      RECT  5.825 44.8825 6.525 46.8625 ;
      RECT  6.525 39.2425 63.025 44.8825 ;
      RECT  6.525 44.8825 63.025 46.8625 ;
      RECT  397.59 114.1225 454.09 116.1725 ;
      RECT  454.79 114.1225 752.635 116.1725 ;
      RECT  397.59 106.745 454.09 114.1225 ;
      RECT  454.79 106.745 459.6475 114.1225 ;
      RECT  397.59 83.7825 454.09 101.0725 ;
      RECT  397.59 101.0725 454.09 103.5425 ;
      RECT  454.09 83.7825 454.79 101.0725 ;
      RECT  454.79 83.7825 457.585 101.0725 ;
      RECT  454.79 101.0725 457.585 103.5425 ;
      RECT  397.59 103.5425 454.09 106.7125 ;
      RECT  454.79 103.5425 457.585 106.7125 ;
      RECT  397.59 106.7125 454.09 106.745 ;
      RECT  454.79 106.7125 457.585 106.745 ;
      RECT  86.805 46.8625 373.615 50.0325 ;
      RECT  86.805 50.0325 373.615 98.5725 ;
      RECT  86.805 98.5725 373.615 101.4925 ;
   END
END    freepdk45_sram_1w1r_32x240
END    LIBRARY
