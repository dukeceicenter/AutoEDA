../macros/freepdk45_sram_1w1r_31x128/freepdk45_sram_1w1r_31x128.lef