VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1rw0r_64x512
   CLASS BLOCK ;
   SIZE 1593.9 BY 218.82 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.625 4.2375 126.76 4.3725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.485 4.2375 129.62 4.3725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.345 4.2375 132.48 4.3725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.205 4.2375 135.34 4.3725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.065 4.2375 138.2 4.3725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.925 4.2375 141.06 4.3725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.785 4.2375 143.92 4.3725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.645 4.2375 146.78 4.3725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.505 4.2375 149.64 4.3725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.365 4.2375 152.5 4.3725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.225 4.2375 155.36 4.3725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.085 4.2375 158.22 4.3725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.945 4.2375 161.08 4.3725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.805 4.2375 163.94 4.3725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.665 4.2375 166.8 4.3725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.525 4.2375 169.66 4.3725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.385 4.2375 172.52 4.3725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.245 4.2375 175.38 4.3725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.105 4.2375 178.24 4.3725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.965 4.2375 181.1 4.3725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.825 4.2375 183.96 4.3725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.685 4.2375 186.82 4.3725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.545 4.2375 189.68 4.3725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.405 4.2375 192.54 4.3725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.265 4.2375 195.4 4.3725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.125 4.2375 198.26 4.3725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.985 4.2375 201.12 4.3725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.845 4.2375 203.98 4.3725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.705 4.2375 206.84 4.3725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.565 4.2375 209.7 4.3725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.425 4.2375 212.56 4.3725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.285 4.2375 215.42 4.3725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.145 4.2375 218.28 4.3725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.005 4.2375 221.14 4.3725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.865 4.2375 224.0 4.3725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.725 4.2375 226.86 4.3725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.585 4.2375 229.72 4.3725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.445 4.2375 232.58 4.3725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.305 4.2375 235.44 4.3725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.165 4.2375 238.3 4.3725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.025 4.2375 241.16 4.3725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.885 4.2375 244.02 4.3725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.745 4.2375 246.88 4.3725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.605 4.2375 249.74 4.3725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.465 4.2375 252.6 4.3725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.325 4.2375 255.46 4.3725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.185 4.2375 258.32 4.3725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.045 4.2375 261.18 4.3725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.905 4.2375 264.04 4.3725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.765 4.2375 266.9 4.3725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.625 4.2375 269.76 4.3725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.485 4.2375 272.62 4.3725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.345 4.2375 275.48 4.3725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.205 4.2375 278.34 4.3725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.065 4.2375 281.2 4.3725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.925 4.2375 284.06 4.3725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.785 4.2375 286.92 4.3725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.645 4.2375 289.78 4.3725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.505 4.2375 292.64 4.3725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.365 4.2375 295.5 4.3725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.225 4.2375 298.36 4.3725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.085 4.2375 301.22 4.3725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.945 4.2375 304.08 4.3725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.805 4.2375 306.94 4.3725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.665 4.2375 309.8 4.3725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.525 4.2375 312.66 4.3725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.385 4.2375 315.52 4.3725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.245 4.2375 318.38 4.3725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.105 4.2375 321.24 4.3725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.965 4.2375 324.1 4.3725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.825 4.2375 326.96 4.3725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.685 4.2375 329.82 4.3725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.545 4.2375 332.68 4.3725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.405 4.2375 335.54 4.3725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.265 4.2375 338.4 4.3725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.125 4.2375 341.26 4.3725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.985 4.2375 344.12 4.3725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.845 4.2375 346.98 4.3725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.705 4.2375 349.84 4.3725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.565 4.2375 352.7 4.3725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.425 4.2375 355.56 4.3725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.285 4.2375 358.42 4.3725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.145 4.2375 361.28 4.3725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.005 4.2375 364.14 4.3725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.865 4.2375 367.0 4.3725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.725 4.2375 369.86 4.3725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.585 4.2375 372.72 4.3725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.445 4.2375 375.58 4.3725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.305 4.2375 378.44 4.3725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.165 4.2375 381.3 4.3725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.025 4.2375 384.16 4.3725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.885 4.2375 387.02 4.3725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.745 4.2375 389.88 4.3725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.605 4.2375 392.74 4.3725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.465 4.2375 395.6 4.3725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.325 4.2375 398.46 4.3725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.185 4.2375 401.32 4.3725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.045 4.2375 404.18 4.3725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.905 4.2375 407.04 4.3725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.765 4.2375 409.9 4.3725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.625 4.2375 412.76 4.3725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.485 4.2375 415.62 4.3725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.345 4.2375 418.48 4.3725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.205 4.2375 421.34 4.3725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.065 4.2375 424.2 4.3725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.925 4.2375 427.06 4.3725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.785 4.2375 429.92 4.3725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.645 4.2375 432.78 4.3725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.505 4.2375 435.64 4.3725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.365 4.2375 438.5 4.3725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.225 4.2375 441.36 4.3725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.085 4.2375 444.22 4.3725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.945 4.2375 447.08 4.3725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.805 4.2375 449.94 4.3725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.665 4.2375 452.8 4.3725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.525 4.2375 455.66 4.3725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.385 4.2375 458.52 4.3725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.245 4.2375 461.38 4.3725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.105 4.2375 464.24 4.3725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.965 4.2375 467.1 4.3725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.825 4.2375 469.96 4.3725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.685 4.2375 472.82 4.3725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.545 4.2375 475.68 4.3725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.405 4.2375 478.54 4.3725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.265 4.2375 481.4 4.3725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.125 4.2375 484.26 4.3725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.985 4.2375 487.12 4.3725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.845 4.2375 489.98 4.3725 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.705 4.2375 492.84 4.3725 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.565 4.2375 495.7 4.3725 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.425 4.2375 498.56 4.3725 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.285 4.2375 501.42 4.3725 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.145 4.2375 504.28 4.3725 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.005 4.2375 507.14 4.3725 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.865 4.2375 510.0 4.3725 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.725 4.2375 512.86 4.3725 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.585 4.2375 515.72 4.3725 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.445 4.2375 518.58 4.3725 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.305 4.2375 521.44 4.3725 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  524.165 4.2375 524.3 4.3725 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.025 4.2375 527.16 4.3725 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  529.885 4.2375 530.02 4.3725 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  532.745 4.2375 532.88 4.3725 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  535.605 4.2375 535.74 4.3725 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  538.465 4.2375 538.6 4.3725 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  541.325 4.2375 541.46 4.3725 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  544.185 4.2375 544.32 4.3725 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  547.045 4.2375 547.18 4.3725 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  549.905 4.2375 550.04 4.3725 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  552.765 4.2375 552.9 4.3725 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  555.625 4.2375 555.76 4.3725 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  558.485 4.2375 558.62 4.3725 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  561.345 4.2375 561.48 4.3725 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  564.205 4.2375 564.34 4.3725 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  567.065 4.2375 567.2 4.3725 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  569.925 4.2375 570.06 4.3725 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  572.785 4.2375 572.92 4.3725 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  575.645 4.2375 575.78 4.3725 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  578.505 4.2375 578.64 4.3725 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  581.365 4.2375 581.5 4.3725 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  584.225 4.2375 584.36 4.3725 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  587.085 4.2375 587.22 4.3725 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  589.945 4.2375 590.08 4.3725 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  592.805 4.2375 592.94 4.3725 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  595.665 4.2375 595.8 4.3725 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  598.525 4.2375 598.66 4.3725 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  601.385 4.2375 601.52 4.3725 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  604.245 4.2375 604.38 4.3725 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  607.105 4.2375 607.24 4.3725 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  609.965 4.2375 610.1 4.3725 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  612.825 4.2375 612.96 4.3725 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  615.685 4.2375 615.82 4.3725 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  618.545 4.2375 618.68 4.3725 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  621.405 4.2375 621.54 4.3725 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  624.265 4.2375 624.4 4.3725 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  627.125 4.2375 627.26 4.3725 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  629.985 4.2375 630.12 4.3725 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  632.845 4.2375 632.98 4.3725 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  635.705 4.2375 635.84 4.3725 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  638.565 4.2375 638.7 4.3725 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  641.425 4.2375 641.56 4.3725 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  644.285 4.2375 644.42 4.3725 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  647.145 4.2375 647.28 4.3725 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  650.005 4.2375 650.14 4.3725 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  652.865 4.2375 653.0 4.3725 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  655.725 4.2375 655.86 4.3725 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  658.585 4.2375 658.72 4.3725 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  661.445 4.2375 661.58 4.3725 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  664.305 4.2375 664.44 4.3725 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  667.165 4.2375 667.3 4.3725 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  670.025 4.2375 670.16 4.3725 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  672.885 4.2375 673.02 4.3725 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  675.745 4.2375 675.88 4.3725 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  678.605 4.2375 678.74 4.3725 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  681.465 4.2375 681.6 4.3725 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  684.325 4.2375 684.46 4.3725 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  687.185 4.2375 687.32 4.3725 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  690.045 4.2375 690.18 4.3725 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  692.905 4.2375 693.04 4.3725 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  695.765 4.2375 695.9 4.3725 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  698.625 4.2375 698.76 4.3725 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  701.485 4.2375 701.62 4.3725 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  704.345 4.2375 704.48 4.3725 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  707.205 4.2375 707.34 4.3725 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  710.065 4.2375 710.2 4.3725 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  712.925 4.2375 713.06 4.3725 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  715.785 4.2375 715.92 4.3725 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  718.645 4.2375 718.78 4.3725 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  721.505 4.2375 721.64 4.3725 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  724.365 4.2375 724.5 4.3725 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  727.225 4.2375 727.36 4.3725 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  730.085 4.2375 730.22 4.3725 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  732.945 4.2375 733.08 4.3725 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  735.805 4.2375 735.94 4.3725 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  738.665 4.2375 738.8 4.3725 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  741.525 4.2375 741.66 4.3725 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  744.385 4.2375 744.52 4.3725 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  747.245 4.2375 747.38 4.3725 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  750.105 4.2375 750.24 4.3725 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  752.965 4.2375 753.1 4.3725 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  755.825 4.2375 755.96 4.3725 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  758.685 4.2375 758.82 4.3725 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  761.545 4.2375 761.68 4.3725 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  764.405 4.2375 764.54 4.3725 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  767.265 4.2375 767.4 4.3725 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  770.125 4.2375 770.26 4.3725 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  772.985 4.2375 773.12 4.3725 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  775.845 4.2375 775.98 4.3725 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  778.705 4.2375 778.84 4.3725 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  781.565 4.2375 781.7 4.3725 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  784.425 4.2375 784.56 4.3725 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  787.285 4.2375 787.42 4.3725 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  790.145 4.2375 790.28 4.3725 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  793.005 4.2375 793.14 4.3725 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  795.865 4.2375 796.0 4.3725 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  798.725 4.2375 798.86 4.3725 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  801.585 4.2375 801.72 4.3725 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  804.445 4.2375 804.58 4.3725 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  807.305 4.2375 807.44 4.3725 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  810.165 4.2375 810.3 4.3725 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  813.025 4.2375 813.16 4.3725 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  815.885 4.2375 816.02 4.3725 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  818.745 4.2375 818.88 4.3725 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  821.605 4.2375 821.74 4.3725 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  824.465 4.2375 824.6 4.3725 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  827.325 4.2375 827.46 4.3725 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  830.185 4.2375 830.32 4.3725 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  833.045 4.2375 833.18 4.3725 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  835.905 4.2375 836.04 4.3725 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  838.765 4.2375 838.9 4.3725 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  841.625 4.2375 841.76 4.3725 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  844.485 4.2375 844.62 4.3725 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  847.345 4.2375 847.48 4.3725 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  850.205 4.2375 850.34 4.3725 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  853.065 4.2375 853.2 4.3725 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  855.925 4.2375 856.06 4.3725 ;
      END
   END din0[255]
   PIN din0[256]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  858.785 4.2375 858.92 4.3725 ;
      END
   END din0[256]
   PIN din0[257]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  861.645 4.2375 861.78 4.3725 ;
      END
   END din0[257]
   PIN din0[258]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  864.505 4.2375 864.64 4.3725 ;
      END
   END din0[258]
   PIN din0[259]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  867.365 4.2375 867.5 4.3725 ;
      END
   END din0[259]
   PIN din0[260]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  870.225 4.2375 870.36 4.3725 ;
      END
   END din0[260]
   PIN din0[261]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  873.085 4.2375 873.22 4.3725 ;
      END
   END din0[261]
   PIN din0[262]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  875.945 4.2375 876.08 4.3725 ;
      END
   END din0[262]
   PIN din0[263]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  878.805 4.2375 878.94 4.3725 ;
      END
   END din0[263]
   PIN din0[264]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  881.665 4.2375 881.8 4.3725 ;
      END
   END din0[264]
   PIN din0[265]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  884.525 4.2375 884.66 4.3725 ;
      END
   END din0[265]
   PIN din0[266]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  887.385 4.2375 887.52 4.3725 ;
      END
   END din0[266]
   PIN din0[267]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  890.245 4.2375 890.38 4.3725 ;
      END
   END din0[267]
   PIN din0[268]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  893.105 4.2375 893.24 4.3725 ;
      END
   END din0[268]
   PIN din0[269]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  895.965 4.2375 896.1 4.3725 ;
      END
   END din0[269]
   PIN din0[270]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  898.825 4.2375 898.96 4.3725 ;
      END
   END din0[270]
   PIN din0[271]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  901.685 4.2375 901.82 4.3725 ;
      END
   END din0[271]
   PIN din0[272]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  904.545 4.2375 904.68 4.3725 ;
      END
   END din0[272]
   PIN din0[273]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  907.405 4.2375 907.54 4.3725 ;
      END
   END din0[273]
   PIN din0[274]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  910.265 4.2375 910.4 4.3725 ;
      END
   END din0[274]
   PIN din0[275]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  913.125 4.2375 913.26 4.3725 ;
      END
   END din0[275]
   PIN din0[276]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  915.985 4.2375 916.12 4.3725 ;
      END
   END din0[276]
   PIN din0[277]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  918.845 4.2375 918.98 4.3725 ;
      END
   END din0[277]
   PIN din0[278]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  921.705 4.2375 921.84 4.3725 ;
      END
   END din0[278]
   PIN din0[279]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  924.565 4.2375 924.7 4.3725 ;
      END
   END din0[279]
   PIN din0[280]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  927.425 4.2375 927.56 4.3725 ;
      END
   END din0[280]
   PIN din0[281]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  930.285 4.2375 930.42 4.3725 ;
      END
   END din0[281]
   PIN din0[282]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  933.145 4.2375 933.28 4.3725 ;
      END
   END din0[282]
   PIN din0[283]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  936.005 4.2375 936.14 4.3725 ;
      END
   END din0[283]
   PIN din0[284]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  938.865 4.2375 939.0 4.3725 ;
      END
   END din0[284]
   PIN din0[285]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  941.725 4.2375 941.86 4.3725 ;
      END
   END din0[285]
   PIN din0[286]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  944.585 4.2375 944.72 4.3725 ;
      END
   END din0[286]
   PIN din0[287]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  947.445 4.2375 947.58 4.3725 ;
      END
   END din0[287]
   PIN din0[288]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  950.305 4.2375 950.44 4.3725 ;
      END
   END din0[288]
   PIN din0[289]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  953.165 4.2375 953.3 4.3725 ;
      END
   END din0[289]
   PIN din0[290]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  956.025 4.2375 956.16 4.3725 ;
      END
   END din0[290]
   PIN din0[291]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  958.885 4.2375 959.02 4.3725 ;
      END
   END din0[291]
   PIN din0[292]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  961.745 4.2375 961.88 4.3725 ;
      END
   END din0[292]
   PIN din0[293]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  964.605 4.2375 964.74 4.3725 ;
      END
   END din0[293]
   PIN din0[294]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  967.465 4.2375 967.6 4.3725 ;
      END
   END din0[294]
   PIN din0[295]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  970.325 4.2375 970.46 4.3725 ;
      END
   END din0[295]
   PIN din0[296]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  973.185 4.2375 973.32 4.3725 ;
      END
   END din0[296]
   PIN din0[297]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  976.045 4.2375 976.18 4.3725 ;
      END
   END din0[297]
   PIN din0[298]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  978.905 4.2375 979.04 4.3725 ;
      END
   END din0[298]
   PIN din0[299]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  981.765 4.2375 981.9 4.3725 ;
      END
   END din0[299]
   PIN din0[300]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  984.625 4.2375 984.76 4.3725 ;
      END
   END din0[300]
   PIN din0[301]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  987.485 4.2375 987.62 4.3725 ;
      END
   END din0[301]
   PIN din0[302]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  990.345 4.2375 990.48 4.3725 ;
      END
   END din0[302]
   PIN din0[303]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  993.205 4.2375 993.34 4.3725 ;
      END
   END din0[303]
   PIN din0[304]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  996.065 4.2375 996.2 4.3725 ;
      END
   END din0[304]
   PIN din0[305]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  998.925 4.2375 999.06 4.3725 ;
      END
   END din0[305]
   PIN din0[306]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1001.785 4.2375 1001.92 4.3725 ;
      END
   END din0[306]
   PIN din0[307]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1004.645 4.2375 1004.78 4.3725 ;
      END
   END din0[307]
   PIN din0[308]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1007.505 4.2375 1007.64 4.3725 ;
      END
   END din0[308]
   PIN din0[309]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1010.365 4.2375 1010.5 4.3725 ;
      END
   END din0[309]
   PIN din0[310]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1013.225 4.2375 1013.36 4.3725 ;
      END
   END din0[310]
   PIN din0[311]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1016.085 4.2375 1016.22 4.3725 ;
      END
   END din0[311]
   PIN din0[312]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1018.945 4.2375 1019.08 4.3725 ;
      END
   END din0[312]
   PIN din0[313]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1021.805 4.2375 1021.94 4.3725 ;
      END
   END din0[313]
   PIN din0[314]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1024.665 4.2375 1024.8 4.3725 ;
      END
   END din0[314]
   PIN din0[315]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1027.525 4.2375 1027.66 4.3725 ;
      END
   END din0[315]
   PIN din0[316]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1030.385 4.2375 1030.52 4.3725 ;
      END
   END din0[316]
   PIN din0[317]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1033.245 4.2375 1033.38 4.3725 ;
      END
   END din0[317]
   PIN din0[318]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1036.105 4.2375 1036.24 4.3725 ;
      END
   END din0[318]
   PIN din0[319]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1038.965 4.2375 1039.1 4.3725 ;
      END
   END din0[319]
   PIN din0[320]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1041.825 4.2375 1041.96 4.3725 ;
      END
   END din0[320]
   PIN din0[321]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1044.685 4.2375 1044.82 4.3725 ;
      END
   END din0[321]
   PIN din0[322]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1047.545 4.2375 1047.68 4.3725 ;
      END
   END din0[322]
   PIN din0[323]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1050.405 4.2375 1050.54 4.3725 ;
      END
   END din0[323]
   PIN din0[324]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1053.265 4.2375 1053.4 4.3725 ;
      END
   END din0[324]
   PIN din0[325]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1056.125 4.2375 1056.26 4.3725 ;
      END
   END din0[325]
   PIN din0[326]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1058.985 4.2375 1059.12 4.3725 ;
      END
   END din0[326]
   PIN din0[327]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1061.845 4.2375 1061.98 4.3725 ;
      END
   END din0[327]
   PIN din0[328]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1064.705 4.2375 1064.84 4.3725 ;
      END
   END din0[328]
   PIN din0[329]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1067.565 4.2375 1067.7 4.3725 ;
      END
   END din0[329]
   PIN din0[330]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1070.425 4.2375 1070.56 4.3725 ;
      END
   END din0[330]
   PIN din0[331]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1073.285 4.2375 1073.42 4.3725 ;
      END
   END din0[331]
   PIN din0[332]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1076.145 4.2375 1076.28 4.3725 ;
      END
   END din0[332]
   PIN din0[333]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1079.005 4.2375 1079.14 4.3725 ;
      END
   END din0[333]
   PIN din0[334]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1081.865 4.2375 1082.0 4.3725 ;
      END
   END din0[334]
   PIN din0[335]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1084.725 4.2375 1084.86 4.3725 ;
      END
   END din0[335]
   PIN din0[336]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1087.585 4.2375 1087.72 4.3725 ;
      END
   END din0[336]
   PIN din0[337]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1090.445 4.2375 1090.58 4.3725 ;
      END
   END din0[337]
   PIN din0[338]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1093.305 4.2375 1093.44 4.3725 ;
      END
   END din0[338]
   PIN din0[339]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1096.165 4.2375 1096.3 4.3725 ;
      END
   END din0[339]
   PIN din0[340]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1099.025 4.2375 1099.16 4.3725 ;
      END
   END din0[340]
   PIN din0[341]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1101.885 4.2375 1102.02 4.3725 ;
      END
   END din0[341]
   PIN din0[342]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1104.745 4.2375 1104.88 4.3725 ;
      END
   END din0[342]
   PIN din0[343]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1107.605 4.2375 1107.74 4.3725 ;
      END
   END din0[343]
   PIN din0[344]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1110.465 4.2375 1110.6 4.3725 ;
      END
   END din0[344]
   PIN din0[345]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1113.325 4.2375 1113.46 4.3725 ;
      END
   END din0[345]
   PIN din0[346]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1116.185 4.2375 1116.32 4.3725 ;
      END
   END din0[346]
   PIN din0[347]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1119.045 4.2375 1119.18 4.3725 ;
      END
   END din0[347]
   PIN din0[348]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1121.905 4.2375 1122.04 4.3725 ;
      END
   END din0[348]
   PIN din0[349]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1124.765 4.2375 1124.9 4.3725 ;
      END
   END din0[349]
   PIN din0[350]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1127.625 4.2375 1127.76 4.3725 ;
      END
   END din0[350]
   PIN din0[351]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1130.485 4.2375 1130.62 4.3725 ;
      END
   END din0[351]
   PIN din0[352]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1133.345 4.2375 1133.48 4.3725 ;
      END
   END din0[352]
   PIN din0[353]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1136.205 4.2375 1136.34 4.3725 ;
      END
   END din0[353]
   PIN din0[354]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1139.065 4.2375 1139.2 4.3725 ;
      END
   END din0[354]
   PIN din0[355]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1141.925 4.2375 1142.06 4.3725 ;
      END
   END din0[355]
   PIN din0[356]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1144.785 4.2375 1144.92 4.3725 ;
      END
   END din0[356]
   PIN din0[357]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1147.645 4.2375 1147.78 4.3725 ;
      END
   END din0[357]
   PIN din0[358]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1150.505 4.2375 1150.64 4.3725 ;
      END
   END din0[358]
   PIN din0[359]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1153.365 4.2375 1153.5 4.3725 ;
      END
   END din0[359]
   PIN din0[360]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1156.225 4.2375 1156.36 4.3725 ;
      END
   END din0[360]
   PIN din0[361]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1159.085 4.2375 1159.22 4.3725 ;
      END
   END din0[361]
   PIN din0[362]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1161.945 4.2375 1162.08 4.3725 ;
      END
   END din0[362]
   PIN din0[363]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1164.805 4.2375 1164.94 4.3725 ;
      END
   END din0[363]
   PIN din0[364]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1167.665 4.2375 1167.8 4.3725 ;
      END
   END din0[364]
   PIN din0[365]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1170.525 4.2375 1170.66 4.3725 ;
      END
   END din0[365]
   PIN din0[366]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1173.385 4.2375 1173.52 4.3725 ;
      END
   END din0[366]
   PIN din0[367]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1176.245 4.2375 1176.38 4.3725 ;
      END
   END din0[367]
   PIN din0[368]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1179.105 4.2375 1179.24 4.3725 ;
      END
   END din0[368]
   PIN din0[369]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1181.965 4.2375 1182.1 4.3725 ;
      END
   END din0[369]
   PIN din0[370]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1184.825 4.2375 1184.96 4.3725 ;
      END
   END din0[370]
   PIN din0[371]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1187.685 4.2375 1187.82 4.3725 ;
      END
   END din0[371]
   PIN din0[372]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1190.545 4.2375 1190.68 4.3725 ;
      END
   END din0[372]
   PIN din0[373]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1193.405 4.2375 1193.54 4.3725 ;
      END
   END din0[373]
   PIN din0[374]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1196.265 4.2375 1196.4 4.3725 ;
      END
   END din0[374]
   PIN din0[375]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1199.125 4.2375 1199.26 4.3725 ;
      END
   END din0[375]
   PIN din0[376]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1201.985 4.2375 1202.12 4.3725 ;
      END
   END din0[376]
   PIN din0[377]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1204.845 4.2375 1204.98 4.3725 ;
      END
   END din0[377]
   PIN din0[378]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1207.705 4.2375 1207.84 4.3725 ;
      END
   END din0[378]
   PIN din0[379]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1210.565 4.2375 1210.7 4.3725 ;
      END
   END din0[379]
   PIN din0[380]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1213.425 4.2375 1213.56 4.3725 ;
      END
   END din0[380]
   PIN din0[381]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1216.285 4.2375 1216.42 4.3725 ;
      END
   END din0[381]
   PIN din0[382]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1219.145 4.2375 1219.28 4.3725 ;
      END
   END din0[382]
   PIN din0[383]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1222.005 4.2375 1222.14 4.3725 ;
      END
   END din0[383]
   PIN din0[384]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1224.865 4.2375 1225.0 4.3725 ;
      END
   END din0[384]
   PIN din0[385]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1227.725 4.2375 1227.86 4.3725 ;
      END
   END din0[385]
   PIN din0[386]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1230.585 4.2375 1230.72 4.3725 ;
      END
   END din0[386]
   PIN din0[387]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1233.445 4.2375 1233.58 4.3725 ;
      END
   END din0[387]
   PIN din0[388]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1236.305 4.2375 1236.44 4.3725 ;
      END
   END din0[388]
   PIN din0[389]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1239.165 4.2375 1239.3 4.3725 ;
      END
   END din0[389]
   PIN din0[390]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1242.025 4.2375 1242.16 4.3725 ;
      END
   END din0[390]
   PIN din0[391]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1244.885 4.2375 1245.02 4.3725 ;
      END
   END din0[391]
   PIN din0[392]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1247.745 4.2375 1247.88 4.3725 ;
      END
   END din0[392]
   PIN din0[393]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1250.605 4.2375 1250.74 4.3725 ;
      END
   END din0[393]
   PIN din0[394]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1253.465 4.2375 1253.6 4.3725 ;
      END
   END din0[394]
   PIN din0[395]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1256.325 4.2375 1256.46 4.3725 ;
      END
   END din0[395]
   PIN din0[396]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1259.185 4.2375 1259.32 4.3725 ;
      END
   END din0[396]
   PIN din0[397]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1262.045 4.2375 1262.18 4.3725 ;
      END
   END din0[397]
   PIN din0[398]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1264.905 4.2375 1265.04 4.3725 ;
      END
   END din0[398]
   PIN din0[399]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1267.765 4.2375 1267.9 4.3725 ;
      END
   END din0[399]
   PIN din0[400]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1270.625 4.2375 1270.76 4.3725 ;
      END
   END din0[400]
   PIN din0[401]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1273.485 4.2375 1273.62 4.3725 ;
      END
   END din0[401]
   PIN din0[402]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1276.345 4.2375 1276.48 4.3725 ;
      END
   END din0[402]
   PIN din0[403]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1279.205 4.2375 1279.34 4.3725 ;
      END
   END din0[403]
   PIN din0[404]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1282.065 4.2375 1282.2 4.3725 ;
      END
   END din0[404]
   PIN din0[405]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1284.925 4.2375 1285.06 4.3725 ;
      END
   END din0[405]
   PIN din0[406]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1287.785 4.2375 1287.92 4.3725 ;
      END
   END din0[406]
   PIN din0[407]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1290.645 4.2375 1290.78 4.3725 ;
      END
   END din0[407]
   PIN din0[408]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1293.505 4.2375 1293.64 4.3725 ;
      END
   END din0[408]
   PIN din0[409]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1296.365 4.2375 1296.5 4.3725 ;
      END
   END din0[409]
   PIN din0[410]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1299.225 4.2375 1299.36 4.3725 ;
      END
   END din0[410]
   PIN din0[411]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1302.085 4.2375 1302.22 4.3725 ;
      END
   END din0[411]
   PIN din0[412]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1304.945 4.2375 1305.08 4.3725 ;
      END
   END din0[412]
   PIN din0[413]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1307.805 4.2375 1307.94 4.3725 ;
      END
   END din0[413]
   PIN din0[414]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1310.665 4.2375 1310.8 4.3725 ;
      END
   END din0[414]
   PIN din0[415]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1313.525 4.2375 1313.66 4.3725 ;
      END
   END din0[415]
   PIN din0[416]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1316.385 4.2375 1316.52 4.3725 ;
      END
   END din0[416]
   PIN din0[417]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1319.245 4.2375 1319.38 4.3725 ;
      END
   END din0[417]
   PIN din0[418]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1322.105 4.2375 1322.24 4.3725 ;
      END
   END din0[418]
   PIN din0[419]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1324.965 4.2375 1325.1 4.3725 ;
      END
   END din0[419]
   PIN din0[420]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1327.825 4.2375 1327.96 4.3725 ;
      END
   END din0[420]
   PIN din0[421]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1330.685 4.2375 1330.82 4.3725 ;
      END
   END din0[421]
   PIN din0[422]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1333.545 4.2375 1333.68 4.3725 ;
      END
   END din0[422]
   PIN din0[423]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1336.405 4.2375 1336.54 4.3725 ;
      END
   END din0[423]
   PIN din0[424]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1339.265 4.2375 1339.4 4.3725 ;
      END
   END din0[424]
   PIN din0[425]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1342.125 4.2375 1342.26 4.3725 ;
      END
   END din0[425]
   PIN din0[426]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1344.985 4.2375 1345.12 4.3725 ;
      END
   END din0[426]
   PIN din0[427]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1347.845 4.2375 1347.98 4.3725 ;
      END
   END din0[427]
   PIN din0[428]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1350.705 4.2375 1350.84 4.3725 ;
      END
   END din0[428]
   PIN din0[429]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1353.565 4.2375 1353.7 4.3725 ;
      END
   END din0[429]
   PIN din0[430]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1356.425 4.2375 1356.56 4.3725 ;
      END
   END din0[430]
   PIN din0[431]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1359.285 4.2375 1359.42 4.3725 ;
      END
   END din0[431]
   PIN din0[432]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1362.145 4.2375 1362.28 4.3725 ;
      END
   END din0[432]
   PIN din0[433]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1365.005 4.2375 1365.14 4.3725 ;
      END
   END din0[433]
   PIN din0[434]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1367.865 4.2375 1368.0 4.3725 ;
      END
   END din0[434]
   PIN din0[435]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1370.725 4.2375 1370.86 4.3725 ;
      END
   END din0[435]
   PIN din0[436]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1373.585 4.2375 1373.72 4.3725 ;
      END
   END din0[436]
   PIN din0[437]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1376.445 4.2375 1376.58 4.3725 ;
      END
   END din0[437]
   PIN din0[438]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1379.305 4.2375 1379.44 4.3725 ;
      END
   END din0[438]
   PIN din0[439]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1382.165 4.2375 1382.3 4.3725 ;
      END
   END din0[439]
   PIN din0[440]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1385.025 4.2375 1385.16 4.3725 ;
      END
   END din0[440]
   PIN din0[441]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1387.885 4.2375 1388.02 4.3725 ;
      END
   END din0[441]
   PIN din0[442]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1390.745 4.2375 1390.88 4.3725 ;
      END
   END din0[442]
   PIN din0[443]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1393.605 4.2375 1393.74 4.3725 ;
      END
   END din0[443]
   PIN din0[444]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1396.465 4.2375 1396.6 4.3725 ;
      END
   END din0[444]
   PIN din0[445]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1399.325 4.2375 1399.46 4.3725 ;
      END
   END din0[445]
   PIN din0[446]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1402.185 4.2375 1402.32 4.3725 ;
      END
   END din0[446]
   PIN din0[447]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1405.045 4.2375 1405.18 4.3725 ;
      END
   END din0[447]
   PIN din0[448]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1407.905 4.2375 1408.04 4.3725 ;
      END
   END din0[448]
   PIN din0[449]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1410.765 4.2375 1410.9 4.3725 ;
      END
   END din0[449]
   PIN din0[450]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1413.625 4.2375 1413.76 4.3725 ;
      END
   END din0[450]
   PIN din0[451]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1416.485 4.2375 1416.62 4.3725 ;
      END
   END din0[451]
   PIN din0[452]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1419.345 4.2375 1419.48 4.3725 ;
      END
   END din0[452]
   PIN din0[453]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1422.205 4.2375 1422.34 4.3725 ;
      END
   END din0[453]
   PIN din0[454]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1425.065 4.2375 1425.2 4.3725 ;
      END
   END din0[454]
   PIN din0[455]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1427.925 4.2375 1428.06 4.3725 ;
      END
   END din0[455]
   PIN din0[456]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1430.785 4.2375 1430.92 4.3725 ;
      END
   END din0[456]
   PIN din0[457]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1433.645 4.2375 1433.78 4.3725 ;
      END
   END din0[457]
   PIN din0[458]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1436.505 4.2375 1436.64 4.3725 ;
      END
   END din0[458]
   PIN din0[459]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1439.365 4.2375 1439.5 4.3725 ;
      END
   END din0[459]
   PIN din0[460]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1442.225 4.2375 1442.36 4.3725 ;
      END
   END din0[460]
   PIN din0[461]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1445.085 4.2375 1445.22 4.3725 ;
      END
   END din0[461]
   PIN din0[462]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1447.945 4.2375 1448.08 4.3725 ;
      END
   END din0[462]
   PIN din0[463]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1450.805 4.2375 1450.94 4.3725 ;
      END
   END din0[463]
   PIN din0[464]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1453.665 4.2375 1453.8 4.3725 ;
      END
   END din0[464]
   PIN din0[465]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1456.525 4.2375 1456.66 4.3725 ;
      END
   END din0[465]
   PIN din0[466]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1459.385 4.2375 1459.52 4.3725 ;
      END
   END din0[466]
   PIN din0[467]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1462.245 4.2375 1462.38 4.3725 ;
      END
   END din0[467]
   PIN din0[468]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1465.105 4.2375 1465.24 4.3725 ;
      END
   END din0[468]
   PIN din0[469]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1467.965 4.2375 1468.1 4.3725 ;
      END
   END din0[469]
   PIN din0[470]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1470.825 4.2375 1470.96 4.3725 ;
      END
   END din0[470]
   PIN din0[471]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1473.685 4.2375 1473.82 4.3725 ;
      END
   END din0[471]
   PIN din0[472]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1476.545 4.2375 1476.68 4.3725 ;
      END
   END din0[472]
   PIN din0[473]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1479.405 4.2375 1479.54 4.3725 ;
      END
   END din0[473]
   PIN din0[474]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1482.265 4.2375 1482.4 4.3725 ;
      END
   END din0[474]
   PIN din0[475]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1485.125 4.2375 1485.26 4.3725 ;
      END
   END din0[475]
   PIN din0[476]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1487.985 4.2375 1488.12 4.3725 ;
      END
   END din0[476]
   PIN din0[477]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1490.845 4.2375 1490.98 4.3725 ;
      END
   END din0[477]
   PIN din0[478]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1493.705 4.2375 1493.84 4.3725 ;
      END
   END din0[478]
   PIN din0[479]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1496.565 4.2375 1496.7 4.3725 ;
      END
   END din0[479]
   PIN din0[480]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1499.425 4.2375 1499.56 4.3725 ;
      END
   END din0[480]
   PIN din0[481]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1502.285 4.2375 1502.42 4.3725 ;
      END
   END din0[481]
   PIN din0[482]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1505.145 4.2375 1505.28 4.3725 ;
      END
   END din0[482]
   PIN din0[483]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1508.005 4.2375 1508.14 4.3725 ;
      END
   END din0[483]
   PIN din0[484]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1510.865 4.2375 1511.0 4.3725 ;
      END
   END din0[484]
   PIN din0[485]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1513.725 4.2375 1513.86 4.3725 ;
      END
   END din0[485]
   PIN din0[486]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1516.585 4.2375 1516.72 4.3725 ;
      END
   END din0[486]
   PIN din0[487]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1519.445 4.2375 1519.58 4.3725 ;
      END
   END din0[487]
   PIN din0[488]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1522.305 4.2375 1522.44 4.3725 ;
      END
   END din0[488]
   PIN din0[489]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1525.165 4.2375 1525.3 4.3725 ;
      END
   END din0[489]
   PIN din0[490]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1528.025 4.2375 1528.16 4.3725 ;
      END
   END din0[490]
   PIN din0[491]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1530.885 4.2375 1531.02 4.3725 ;
      END
   END din0[491]
   PIN din0[492]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1533.745 4.2375 1533.88 4.3725 ;
      END
   END din0[492]
   PIN din0[493]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1536.605 4.2375 1536.74 4.3725 ;
      END
   END din0[493]
   PIN din0[494]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1539.465 4.2375 1539.6 4.3725 ;
      END
   END din0[494]
   PIN din0[495]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1542.325 4.2375 1542.46 4.3725 ;
      END
   END din0[495]
   PIN din0[496]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1545.185 4.2375 1545.32 4.3725 ;
      END
   END din0[496]
   PIN din0[497]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1548.045 4.2375 1548.18 4.3725 ;
      END
   END din0[497]
   PIN din0[498]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1550.905 4.2375 1551.04 4.3725 ;
      END
   END din0[498]
   PIN din0[499]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1553.765 4.2375 1553.9 4.3725 ;
      END
   END din0[499]
   PIN din0[500]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1556.625 4.2375 1556.76 4.3725 ;
      END
   END din0[500]
   PIN din0[501]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1559.485 4.2375 1559.62 4.3725 ;
      END
   END din0[501]
   PIN din0[502]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1562.345 4.2375 1562.48 4.3725 ;
      END
   END din0[502]
   PIN din0[503]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1565.205 4.2375 1565.34 4.3725 ;
      END
   END din0[503]
   PIN din0[504]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1568.065 4.2375 1568.2 4.3725 ;
      END
   END din0[504]
   PIN din0[505]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1570.925 4.2375 1571.06 4.3725 ;
      END
   END din0[505]
   PIN din0[506]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1573.785 4.2375 1573.92 4.3725 ;
      END
   END din0[506]
   PIN din0[507]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1576.645 4.2375 1576.78 4.3725 ;
      END
   END din0[507]
   PIN din0[508]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1579.505 4.2375 1579.64 4.3725 ;
      END
   END din0[508]
   PIN din0[509]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1582.365 4.2375 1582.5 4.3725 ;
      END
   END din0[509]
   PIN din0[510]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1585.225 4.2375 1585.36 4.3725 ;
      END
   END din0[510]
   PIN din0[511]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1588.085 4.2375 1588.22 4.3725 ;
      END
   END din0[511]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.905 148.7225 121.04 148.8575 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.905 151.4525 121.04 151.5875 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.905 153.6625 121.04 153.7975 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.905 156.3925 121.04 156.5275 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.905 158.6025 121.04 158.7375 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.905 161.3325 121.04 161.4675 ;
      END
   END addr0[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  3.39 104.0025 3.525 104.1375 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  3.39 106.7325 3.525 106.8675 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  9.6325 104.0875 9.7675 104.2225 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.3925 115.65 163.5275 115.785 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.0975 115.65 164.2325 115.785 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.8025 115.65 164.9375 115.785 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.5075 115.65 165.6425 115.785 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.2125 115.65 166.3475 115.785 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.9175 115.65 167.0525 115.785 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.6225 115.65 167.7575 115.785 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.3275 115.65 168.4625 115.785 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.0325 115.65 169.1675 115.785 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.7375 115.65 169.8725 115.785 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.4425 115.65 170.5775 115.785 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.1475 115.65 171.2825 115.785 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.8525 115.65 171.9875 115.785 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.5575 115.65 172.6925 115.785 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.2625 115.65 173.3975 115.785 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.9675 115.65 174.1025 115.785 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.6725 115.65 174.8075 115.785 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.3775 115.65 175.5125 115.785 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.0825 115.65 176.2175 115.785 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.7875 115.65 176.9225 115.785 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.4925 115.65 177.6275 115.785 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.1975 115.65 178.3325 115.785 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.9025 115.65 179.0375 115.785 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.6075 115.65 179.7425 115.785 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.3125 115.65 180.4475 115.785 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.0175 115.65 181.1525 115.785 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.7225 115.65 181.8575 115.785 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.4275 115.65 182.5625 115.785 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.1325 115.65 183.2675 115.785 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.8375 115.65 183.9725 115.785 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.5425 115.65 184.6775 115.785 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.2475 115.65 185.3825 115.785 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.9525 115.65 186.0875 115.785 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.6575 115.65 186.7925 115.785 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.3625 115.65 187.4975 115.785 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.0675 115.65 188.2025 115.785 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.7725 115.65 188.9075 115.785 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.4775 115.65 189.6125 115.785 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.1825 115.65 190.3175 115.785 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.8875 115.65 191.0225 115.785 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.5925 115.65 191.7275 115.785 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.2975 115.65 192.4325 115.785 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.0025 115.65 193.1375 115.785 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.7075 115.65 193.8425 115.785 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.4125 115.65 194.5475 115.785 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.1175 115.65 195.2525 115.785 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.8225 115.65 195.9575 115.785 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.5275 115.65 196.6625 115.785 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.2325 115.65 197.3675 115.785 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.9375 115.65 198.0725 115.785 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.6425 115.65 198.7775 115.785 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.3475 115.65 199.4825 115.785 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.0525 115.65 200.1875 115.785 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.7575 115.65 200.8925 115.785 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.4625 115.65 201.5975 115.785 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.1675 115.65 202.3025 115.785 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.8725 115.65 203.0075 115.785 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.5775 115.65 203.7125 115.785 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.2825 115.65 204.4175 115.785 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.9875 115.65 205.1225 115.785 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.6925 115.65 205.8275 115.785 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.3975 115.65 206.5325 115.785 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.1025 115.65 207.2375 115.785 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.8075 115.65 207.9425 115.785 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.5125 115.65 208.6475 115.785 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.2175 115.65 209.3525 115.785 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.9225 115.65 210.0575 115.785 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.6275 115.65 210.7625 115.785 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.3325 115.65 211.4675 115.785 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.0375 115.65 212.1725 115.785 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.7425 115.65 212.8775 115.785 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.4475 115.65 213.5825 115.785 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.1525 115.65 214.2875 115.785 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.8575 115.65 214.9925 115.785 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.5625 115.65 215.6975 115.785 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.2675 115.65 216.4025 115.785 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.9725 115.65 217.1075 115.785 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.6775 115.65 217.8125 115.785 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.3825 115.65 218.5175 115.785 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.0875 115.65 219.2225 115.785 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.7925 115.65 219.9275 115.785 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.4975 115.65 220.6325 115.785 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.2025 115.65 221.3375 115.785 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.9075 115.65 222.0425 115.785 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.6125 115.65 222.7475 115.785 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.3175 115.65 223.4525 115.785 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.0225 115.65 224.1575 115.785 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.7275 115.65 224.8625 115.785 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.4325 115.65 225.5675 115.785 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.1375 115.65 226.2725 115.785 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.8425 115.65 226.9775 115.785 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.5475 115.65 227.6825 115.785 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.2525 115.65 228.3875 115.785 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.9575 115.65 229.0925 115.785 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.6625 115.65 229.7975 115.785 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.3675 115.65 230.5025 115.785 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.0725 115.65 231.2075 115.785 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.7775 115.65 231.9125 115.785 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.4825 115.65 232.6175 115.785 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.1875 115.65 233.3225 115.785 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.8925 115.65 234.0275 115.785 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.5975 115.65 234.7325 115.785 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.3025 115.65 235.4375 115.785 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.0075 115.65 236.1425 115.785 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.7125 115.65 236.8475 115.785 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.4175 115.65 237.5525 115.785 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.1225 115.65 238.2575 115.785 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.8275 115.65 238.9625 115.785 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.5325 115.65 239.6675 115.785 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.2375 115.65 240.3725 115.785 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.9425 115.65 241.0775 115.785 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.6475 115.65 241.7825 115.785 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.3525 115.65 242.4875 115.785 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.0575 115.65 243.1925 115.785 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.7625 115.65 243.8975 115.785 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.4675 115.65 244.6025 115.785 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.1725 115.65 245.3075 115.785 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.8775 115.65 246.0125 115.785 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.5825 115.65 246.7175 115.785 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.2875 115.65 247.4225 115.785 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.9925 115.65 248.1275 115.785 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.6975 115.65 248.8325 115.785 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.4025 115.65 249.5375 115.785 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.1075 115.65 250.2425 115.785 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.8125 115.65 250.9475 115.785 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.5175 115.65 251.6525 115.785 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.2225 115.65 252.3575 115.785 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.9275 115.65 253.0625 115.785 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.6325 115.65 253.7675 115.785 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.3375 115.65 254.4725 115.785 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.0425 115.65 255.1775 115.785 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.7475 115.65 255.8825 115.785 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.4525 115.65 256.5875 115.785 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.1575 115.65 257.2925 115.785 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.8625 115.65 257.9975 115.785 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.5675 115.65 258.7025 115.785 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.2725 115.65 259.4075 115.785 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.9775 115.65 260.1125 115.785 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.6825 115.65 260.8175 115.785 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.3875 115.65 261.5225 115.785 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.0925 115.65 262.2275 115.785 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.7975 115.65 262.9325 115.785 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.5025 115.65 263.6375 115.785 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.2075 115.65 264.3425 115.785 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.9125 115.65 265.0475 115.785 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.6175 115.65 265.7525 115.785 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.3225 115.65 266.4575 115.785 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.0275 115.65 267.1625 115.785 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.7325 115.65 267.8675 115.785 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.4375 115.65 268.5725 115.785 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.1425 115.65 269.2775 115.785 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.8475 115.65 269.9825 115.785 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.5525 115.65 270.6875 115.785 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.2575 115.65 271.3925 115.785 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.9625 115.65 272.0975 115.785 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.6675 115.65 272.8025 115.785 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.3725 115.65 273.5075 115.785 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.0775 115.65 274.2125 115.785 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.7825 115.65 274.9175 115.785 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.4875 115.65 275.6225 115.785 ;
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.1925 115.65 276.3275 115.785 ;
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.8975 115.65 277.0325 115.785 ;
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.6025 115.65 277.7375 115.785 ;
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.3075 115.65 278.4425 115.785 ;
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.0125 115.65 279.1475 115.785 ;
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  279.7175 115.65 279.8525 115.785 ;
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.4225 115.65 280.5575 115.785 ;
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.1275 115.65 281.2625 115.785 ;
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.8325 115.65 281.9675 115.785 ;
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  282.5375 115.65 282.6725 115.785 ;
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.2425 115.65 283.3775 115.785 ;
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.9475 115.65 284.0825 115.785 ;
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.6525 115.65 284.7875 115.785 ;
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  285.3575 115.65 285.4925 115.785 ;
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.0625 115.65 286.1975 115.785 ;
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.7675 115.65 286.9025 115.785 ;
      END
   END dout0[175]
   PIN dout0[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.4725 115.65 287.6075 115.785 ;
      END
   END dout0[176]
   PIN dout0[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.1775 115.65 288.3125 115.785 ;
      END
   END dout0[177]
   PIN dout0[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.8825 115.65 289.0175 115.785 ;
      END
   END dout0[178]
   PIN dout0[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.5875 115.65 289.7225 115.785 ;
      END
   END dout0[179]
   PIN dout0[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.2925 115.65 290.4275 115.785 ;
      END
   END dout0[180]
   PIN dout0[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.9975 115.65 291.1325 115.785 ;
      END
   END dout0[181]
   PIN dout0[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.7025 115.65 291.8375 115.785 ;
      END
   END dout0[182]
   PIN dout0[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.4075 115.65 292.5425 115.785 ;
      END
   END dout0[183]
   PIN dout0[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.1125 115.65 293.2475 115.785 ;
      END
   END dout0[184]
   PIN dout0[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.8175 115.65 293.9525 115.785 ;
      END
   END dout0[185]
   PIN dout0[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.5225 115.65 294.6575 115.785 ;
      END
   END dout0[186]
   PIN dout0[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.2275 115.65 295.3625 115.785 ;
      END
   END dout0[187]
   PIN dout0[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.9325 115.65 296.0675 115.785 ;
      END
   END dout0[188]
   PIN dout0[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.6375 115.65 296.7725 115.785 ;
      END
   END dout0[189]
   PIN dout0[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.3425 115.65 297.4775 115.785 ;
      END
   END dout0[190]
   PIN dout0[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.0475 115.65 298.1825 115.785 ;
      END
   END dout0[191]
   PIN dout0[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.7525 115.65 298.8875 115.785 ;
      END
   END dout0[192]
   PIN dout0[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  299.4575 115.65 299.5925 115.785 ;
      END
   END dout0[193]
   PIN dout0[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.1625 115.65 300.2975 115.785 ;
      END
   END dout0[194]
   PIN dout0[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.8675 115.65 301.0025 115.785 ;
      END
   END dout0[195]
   PIN dout0[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.5725 115.65 301.7075 115.785 ;
      END
   END dout0[196]
   PIN dout0[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  302.2775 115.65 302.4125 115.785 ;
      END
   END dout0[197]
   PIN dout0[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  302.9825 115.65 303.1175 115.785 ;
      END
   END dout0[198]
   PIN dout0[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.6875 115.65 303.8225 115.785 ;
      END
   END dout0[199]
   PIN dout0[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.3925 115.65 304.5275 115.785 ;
      END
   END dout0[200]
   PIN dout0[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.0975 115.65 305.2325 115.785 ;
      END
   END dout0[201]
   PIN dout0[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.8025 115.65 305.9375 115.785 ;
      END
   END dout0[202]
   PIN dout0[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.5075 115.65 306.6425 115.785 ;
      END
   END dout0[203]
   PIN dout0[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.2125 115.65 307.3475 115.785 ;
      END
   END dout0[204]
   PIN dout0[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.9175 115.65 308.0525 115.785 ;
      END
   END dout0[205]
   PIN dout0[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.6225 115.65 308.7575 115.785 ;
      END
   END dout0[206]
   PIN dout0[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.3275 115.65 309.4625 115.785 ;
      END
   END dout0[207]
   PIN dout0[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.0325 115.65 310.1675 115.785 ;
      END
   END dout0[208]
   PIN dout0[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.7375 115.65 310.8725 115.785 ;
      END
   END dout0[209]
   PIN dout0[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.4425 115.65 311.5775 115.785 ;
      END
   END dout0[210]
   PIN dout0[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.1475 115.65 312.2825 115.785 ;
      END
   END dout0[211]
   PIN dout0[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.8525 115.65 312.9875 115.785 ;
      END
   END dout0[212]
   PIN dout0[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.5575 115.65 313.6925 115.785 ;
      END
   END dout0[213]
   PIN dout0[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.2625 115.65 314.3975 115.785 ;
      END
   END dout0[214]
   PIN dout0[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.9675 115.65 315.1025 115.785 ;
      END
   END dout0[215]
   PIN dout0[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.6725 115.65 315.8075 115.785 ;
      END
   END dout0[216]
   PIN dout0[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.3775 115.65 316.5125 115.785 ;
      END
   END dout0[217]
   PIN dout0[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.0825 115.65 317.2175 115.785 ;
      END
   END dout0[218]
   PIN dout0[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.7875 115.65 317.9225 115.785 ;
      END
   END dout0[219]
   PIN dout0[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.4925 115.65 318.6275 115.785 ;
      END
   END dout0[220]
   PIN dout0[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.1975 115.65 319.3325 115.785 ;
      END
   END dout0[221]
   PIN dout0[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.9025 115.65 320.0375 115.785 ;
      END
   END dout0[222]
   PIN dout0[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.6075 115.65 320.7425 115.785 ;
      END
   END dout0[223]
   PIN dout0[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.3125 115.65 321.4475 115.785 ;
      END
   END dout0[224]
   PIN dout0[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  322.0175 115.65 322.1525 115.785 ;
      END
   END dout0[225]
   PIN dout0[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  322.7225 115.65 322.8575 115.785 ;
      END
   END dout0[226]
   PIN dout0[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.4275 115.65 323.5625 115.785 ;
      END
   END dout0[227]
   PIN dout0[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.1325 115.65 324.2675 115.785 ;
      END
   END dout0[228]
   PIN dout0[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.8375 115.65 324.9725 115.785 ;
      END
   END dout0[229]
   PIN dout0[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  325.5425 115.65 325.6775 115.785 ;
      END
   END dout0[230]
   PIN dout0[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.2475 115.65 326.3825 115.785 ;
      END
   END dout0[231]
   PIN dout0[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.9525 115.65 327.0875 115.785 ;
      END
   END dout0[232]
   PIN dout0[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.6575 115.65 327.7925 115.785 ;
      END
   END dout0[233]
   PIN dout0[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.3625 115.65 328.4975 115.785 ;
      END
   END dout0[234]
   PIN dout0[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.0675 115.65 329.2025 115.785 ;
      END
   END dout0[235]
   PIN dout0[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.7725 115.65 329.9075 115.785 ;
      END
   END dout0[236]
   PIN dout0[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.4775 115.65 330.6125 115.785 ;
      END
   END dout0[237]
   PIN dout0[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.1825 115.65 331.3175 115.785 ;
      END
   END dout0[238]
   PIN dout0[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.8875 115.65 332.0225 115.785 ;
      END
   END dout0[239]
   PIN dout0[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.5925 115.65 332.7275 115.785 ;
      END
   END dout0[240]
   PIN dout0[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.2975 115.65 333.4325 115.785 ;
      END
   END dout0[241]
   PIN dout0[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.0025 115.65 334.1375 115.785 ;
      END
   END dout0[242]
   PIN dout0[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.7075 115.65 334.8425 115.785 ;
      END
   END dout0[243]
   PIN dout0[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.4125 115.65 335.5475 115.785 ;
      END
   END dout0[244]
   PIN dout0[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.1175 115.65 336.2525 115.785 ;
      END
   END dout0[245]
   PIN dout0[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.8225 115.65 336.9575 115.785 ;
      END
   END dout0[246]
   PIN dout0[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.5275 115.65 337.6625 115.785 ;
      END
   END dout0[247]
   PIN dout0[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.2325 115.65 338.3675 115.785 ;
      END
   END dout0[248]
   PIN dout0[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.9375 115.65 339.0725 115.785 ;
      END
   END dout0[249]
   PIN dout0[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.6425 115.65 339.7775 115.785 ;
      END
   END dout0[250]
   PIN dout0[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.3475 115.65 340.4825 115.785 ;
      END
   END dout0[251]
   PIN dout0[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.0525 115.65 341.1875 115.785 ;
      END
   END dout0[252]
   PIN dout0[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.7575 115.65 341.8925 115.785 ;
      END
   END dout0[253]
   PIN dout0[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  342.4625 115.65 342.5975 115.785 ;
      END
   END dout0[254]
   PIN dout0[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.1675 115.65 343.3025 115.785 ;
      END
   END dout0[255]
   PIN dout0[256]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.8725 115.65 344.0075 115.785 ;
      END
   END dout0[256]
   PIN dout0[257]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.5775 115.65 344.7125 115.785 ;
      END
   END dout0[257]
   PIN dout0[258]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.2825 115.65 345.4175 115.785 ;
      END
   END dout0[258]
   PIN dout0[259]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  345.9875 115.65 346.1225 115.785 ;
      END
   END dout0[259]
   PIN dout0[260]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.6925 115.65 346.8275 115.785 ;
      END
   END dout0[260]
   PIN dout0[261]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.3975 115.65 347.5325 115.785 ;
      END
   END dout0[261]
   PIN dout0[262]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.1025 115.65 348.2375 115.785 ;
      END
   END dout0[262]
   PIN dout0[263]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.8075 115.65 348.9425 115.785 ;
      END
   END dout0[263]
   PIN dout0[264]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.5125 115.65 349.6475 115.785 ;
      END
   END dout0[264]
   PIN dout0[265]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.2175 115.65 350.3525 115.785 ;
      END
   END dout0[265]
   PIN dout0[266]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.9225 115.65 351.0575 115.785 ;
      END
   END dout0[266]
   PIN dout0[267]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  351.6275 115.65 351.7625 115.785 ;
      END
   END dout0[267]
   PIN dout0[268]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.3325 115.65 352.4675 115.785 ;
      END
   END dout0[268]
   PIN dout0[269]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.0375 115.65 353.1725 115.785 ;
      END
   END dout0[269]
   PIN dout0[270]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.7425 115.65 353.8775 115.785 ;
      END
   END dout0[270]
   PIN dout0[271]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.4475 115.65 354.5825 115.785 ;
      END
   END dout0[271]
   PIN dout0[272]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.1525 115.65 355.2875 115.785 ;
      END
   END dout0[272]
   PIN dout0[273]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.8575 115.65 355.9925 115.785 ;
      END
   END dout0[273]
   PIN dout0[274]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.5625 115.65 356.6975 115.785 ;
      END
   END dout0[274]
   PIN dout0[275]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.2675 115.65 357.4025 115.785 ;
      END
   END dout0[275]
   PIN dout0[276]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.9725 115.65 358.1075 115.785 ;
      END
   END dout0[276]
   PIN dout0[277]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.6775 115.65 358.8125 115.785 ;
      END
   END dout0[277]
   PIN dout0[278]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.3825 115.65 359.5175 115.785 ;
      END
   END dout0[278]
   PIN dout0[279]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.0875 115.65 360.2225 115.785 ;
      END
   END dout0[279]
   PIN dout0[280]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.7925 115.65 360.9275 115.785 ;
      END
   END dout0[280]
   PIN dout0[281]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.4975 115.65 361.6325 115.785 ;
      END
   END dout0[281]
   PIN dout0[282]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.2025 115.65 362.3375 115.785 ;
      END
   END dout0[282]
   PIN dout0[283]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  362.9075 115.65 363.0425 115.785 ;
      END
   END dout0[283]
   PIN dout0[284]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.6125 115.65 363.7475 115.785 ;
      END
   END dout0[284]
   PIN dout0[285]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.3175 115.65 364.4525 115.785 ;
      END
   END dout0[285]
   PIN dout0[286]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.0225 115.65 365.1575 115.785 ;
      END
   END dout0[286]
   PIN dout0[287]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.7275 115.65 365.8625 115.785 ;
      END
   END dout0[287]
   PIN dout0[288]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.4325 115.65 366.5675 115.785 ;
      END
   END dout0[288]
   PIN dout0[289]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.1375 115.65 367.2725 115.785 ;
      END
   END dout0[289]
   PIN dout0[290]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.8425 115.65 367.9775 115.785 ;
      END
   END dout0[290]
   PIN dout0[291]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.5475 115.65 368.6825 115.785 ;
      END
   END dout0[291]
   PIN dout0[292]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.2525 115.65 369.3875 115.785 ;
      END
   END dout0[292]
   PIN dout0[293]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.9575 115.65 370.0925 115.785 ;
      END
   END dout0[293]
   PIN dout0[294]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.6625 115.65 370.7975 115.785 ;
      END
   END dout0[294]
   PIN dout0[295]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  371.3675 115.65 371.5025 115.785 ;
      END
   END dout0[295]
   PIN dout0[296]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.0725 115.65 372.2075 115.785 ;
      END
   END dout0[296]
   PIN dout0[297]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.7775 115.65 372.9125 115.785 ;
      END
   END dout0[297]
   PIN dout0[298]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.4825 115.65 373.6175 115.785 ;
      END
   END dout0[298]
   PIN dout0[299]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.1875 115.65 374.3225 115.785 ;
      END
   END dout0[299]
   PIN dout0[300]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.8925 115.65 375.0275 115.785 ;
      END
   END dout0[300]
   PIN dout0[301]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.5975 115.65 375.7325 115.785 ;
      END
   END dout0[301]
   PIN dout0[302]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  376.3025 115.65 376.4375 115.785 ;
      END
   END dout0[302]
   PIN dout0[303]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.0075 115.65 377.1425 115.785 ;
      END
   END dout0[303]
   PIN dout0[304]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.7125 115.65 377.8475 115.785 ;
      END
   END dout0[304]
   PIN dout0[305]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.4175 115.65 378.5525 115.785 ;
      END
   END dout0[305]
   PIN dout0[306]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  379.1225 115.65 379.2575 115.785 ;
      END
   END dout0[306]
   PIN dout0[307]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  379.8275 115.65 379.9625 115.785 ;
      END
   END dout0[307]
   PIN dout0[308]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.5325 115.65 380.6675 115.785 ;
      END
   END dout0[308]
   PIN dout0[309]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.2375 115.65 381.3725 115.785 ;
      END
   END dout0[309]
   PIN dout0[310]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.9425 115.65 382.0775 115.785 ;
      END
   END dout0[310]
   PIN dout0[311]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  382.6475 115.65 382.7825 115.785 ;
      END
   END dout0[311]
   PIN dout0[312]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.3525 115.65 383.4875 115.785 ;
      END
   END dout0[312]
   PIN dout0[313]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.0575 115.65 384.1925 115.785 ;
      END
   END dout0[313]
   PIN dout0[314]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.7625 115.65 384.8975 115.785 ;
      END
   END dout0[314]
   PIN dout0[315]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  385.4675 115.65 385.6025 115.785 ;
      END
   END dout0[315]
   PIN dout0[316]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.1725 115.65 386.3075 115.785 ;
      END
   END dout0[316]
   PIN dout0[317]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.8775 115.65 387.0125 115.785 ;
      END
   END dout0[317]
   PIN dout0[318]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  387.5825 115.65 387.7175 115.785 ;
      END
   END dout0[318]
   PIN dout0[319]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  388.2875 115.65 388.4225 115.785 ;
      END
   END dout0[319]
   PIN dout0[320]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  388.9925 115.65 389.1275 115.785 ;
      END
   END dout0[320]
   PIN dout0[321]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.6975 115.65 389.8325 115.785 ;
      END
   END dout0[321]
   PIN dout0[322]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  390.4025 115.65 390.5375 115.785 ;
      END
   END dout0[322]
   PIN dout0[323]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  391.1075 115.65 391.2425 115.785 ;
      END
   END dout0[323]
   PIN dout0[324]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  391.8125 115.65 391.9475 115.785 ;
      END
   END dout0[324]
   PIN dout0[325]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.5175 115.65 392.6525 115.785 ;
      END
   END dout0[325]
   PIN dout0[326]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.2225 115.65 393.3575 115.785 ;
      END
   END dout0[326]
   PIN dout0[327]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.9275 115.65 394.0625 115.785 ;
      END
   END dout0[327]
   PIN dout0[328]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.6325 115.65 394.7675 115.785 ;
      END
   END dout0[328]
   PIN dout0[329]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.3375 115.65 395.4725 115.785 ;
      END
   END dout0[329]
   PIN dout0[330]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.0425 115.65 396.1775 115.785 ;
      END
   END dout0[330]
   PIN dout0[331]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.7475 115.65 396.8825 115.785 ;
      END
   END dout0[331]
   PIN dout0[332]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.4525 115.65 397.5875 115.785 ;
      END
   END dout0[332]
   PIN dout0[333]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.1575 115.65 398.2925 115.785 ;
      END
   END dout0[333]
   PIN dout0[334]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.8625 115.65 398.9975 115.785 ;
      END
   END dout0[334]
   PIN dout0[335]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.5675 115.65 399.7025 115.785 ;
      END
   END dout0[335]
   PIN dout0[336]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.2725 115.65 400.4075 115.785 ;
      END
   END dout0[336]
   PIN dout0[337]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.9775 115.65 401.1125 115.785 ;
      END
   END dout0[337]
   PIN dout0[338]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.6825 115.65 401.8175 115.785 ;
      END
   END dout0[338]
   PIN dout0[339]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  402.3875 115.65 402.5225 115.785 ;
      END
   END dout0[339]
   PIN dout0[340]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.0925 115.65 403.2275 115.785 ;
      END
   END dout0[340]
   PIN dout0[341]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.7975 115.65 403.9325 115.785 ;
      END
   END dout0[341]
   PIN dout0[342]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.5025 115.65 404.6375 115.785 ;
      END
   END dout0[342]
   PIN dout0[343]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  405.2075 115.65 405.3425 115.785 ;
      END
   END dout0[343]
   PIN dout0[344]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  405.9125 115.65 406.0475 115.785 ;
      END
   END dout0[344]
   PIN dout0[345]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.6175 115.65 406.7525 115.785 ;
      END
   END dout0[345]
   PIN dout0[346]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.3225 115.65 407.4575 115.785 ;
      END
   END dout0[346]
   PIN dout0[347]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  408.0275 115.65 408.1625 115.785 ;
      END
   END dout0[347]
   PIN dout0[348]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  408.7325 115.65 408.8675 115.785 ;
      END
   END dout0[348]
   PIN dout0[349]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.4375 115.65 409.5725 115.785 ;
      END
   END dout0[349]
   PIN dout0[350]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.1425 115.65 410.2775 115.785 ;
      END
   END dout0[350]
   PIN dout0[351]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.8475 115.65 410.9825 115.785 ;
      END
   END dout0[351]
   PIN dout0[352]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  411.5525 115.65 411.6875 115.785 ;
      END
   END dout0[352]
   PIN dout0[353]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.2575 115.65 412.3925 115.785 ;
      END
   END dout0[353]
   PIN dout0[354]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.9625 115.65 413.0975 115.785 ;
      END
   END dout0[354]
   PIN dout0[355]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  413.6675 115.65 413.8025 115.785 ;
      END
   END dout0[355]
   PIN dout0[356]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  414.3725 115.65 414.5075 115.785 ;
      END
   END dout0[356]
   PIN dout0[357]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.0775 115.65 415.2125 115.785 ;
      END
   END dout0[357]
   PIN dout0[358]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.7825 115.65 415.9175 115.785 ;
      END
   END dout0[358]
   PIN dout0[359]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  416.4875 115.65 416.6225 115.785 ;
      END
   END dout0[359]
   PIN dout0[360]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.1925 115.65 417.3275 115.785 ;
      END
   END dout0[360]
   PIN dout0[361]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.8975 115.65 418.0325 115.785 ;
      END
   END dout0[361]
   PIN dout0[362]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.6025 115.65 418.7375 115.785 ;
      END
   END dout0[362]
   PIN dout0[363]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  419.3075 115.65 419.4425 115.785 ;
      END
   END dout0[363]
   PIN dout0[364]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.0125 115.65 420.1475 115.785 ;
      END
   END dout0[364]
   PIN dout0[365]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.7175 115.65 420.8525 115.785 ;
      END
   END dout0[365]
   PIN dout0[366]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.4225 115.65 421.5575 115.785 ;
      END
   END dout0[366]
   PIN dout0[367]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  422.1275 115.65 422.2625 115.785 ;
      END
   END dout0[367]
   PIN dout0[368]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  422.8325 115.65 422.9675 115.785 ;
      END
   END dout0[368]
   PIN dout0[369]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.5375 115.65 423.6725 115.785 ;
      END
   END dout0[369]
   PIN dout0[370]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.2425 115.65 424.3775 115.785 ;
      END
   END dout0[370]
   PIN dout0[371]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.9475 115.65 425.0825 115.785 ;
      END
   END dout0[371]
   PIN dout0[372]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  425.6525 115.65 425.7875 115.785 ;
      END
   END dout0[372]
   PIN dout0[373]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.3575 115.65 426.4925 115.785 ;
      END
   END dout0[373]
   PIN dout0[374]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.0625 115.65 427.1975 115.785 ;
      END
   END dout0[374]
   PIN dout0[375]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.7675 115.65 427.9025 115.785 ;
      END
   END dout0[375]
   PIN dout0[376]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  428.4725 115.65 428.6075 115.785 ;
      END
   END dout0[376]
   PIN dout0[377]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.1775 115.65 429.3125 115.785 ;
      END
   END dout0[377]
   PIN dout0[378]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.8825 115.65 430.0175 115.785 ;
      END
   END dout0[378]
   PIN dout0[379]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  430.5875 115.65 430.7225 115.785 ;
      END
   END dout0[379]
   PIN dout0[380]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  431.2925 115.65 431.4275 115.785 ;
      END
   END dout0[380]
   PIN dout0[381]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  431.9975 115.65 432.1325 115.785 ;
      END
   END dout0[381]
   PIN dout0[382]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.7025 115.65 432.8375 115.785 ;
      END
   END dout0[382]
   PIN dout0[383]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  433.4075 115.65 433.5425 115.785 ;
      END
   END dout0[383]
   PIN dout0[384]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  434.1125 115.65 434.2475 115.785 ;
      END
   END dout0[384]
   PIN dout0[385]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  434.8175 115.65 434.9525 115.785 ;
      END
   END dout0[385]
   PIN dout0[386]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.5225 115.65 435.6575 115.785 ;
      END
   END dout0[386]
   PIN dout0[387]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  436.2275 115.65 436.3625 115.785 ;
      END
   END dout0[387]
   PIN dout0[388]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  436.9325 115.65 437.0675 115.785 ;
      END
   END dout0[388]
   PIN dout0[389]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  437.6375 115.65 437.7725 115.785 ;
      END
   END dout0[389]
   PIN dout0[390]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.3425 115.65 438.4775 115.785 ;
      END
   END dout0[390]
   PIN dout0[391]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  439.0475 115.65 439.1825 115.785 ;
      END
   END dout0[391]
   PIN dout0[392]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  439.7525 115.65 439.8875 115.785 ;
      END
   END dout0[392]
   PIN dout0[393]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.4575 115.65 440.5925 115.785 ;
      END
   END dout0[393]
   PIN dout0[394]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.1625 115.65 441.2975 115.785 ;
      END
   END dout0[394]
   PIN dout0[395]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.8675 115.65 442.0025 115.785 ;
      END
   END dout0[395]
   PIN dout0[396]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  442.5725 115.65 442.7075 115.785 ;
      END
   END dout0[396]
   PIN dout0[397]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.2775 115.65 443.4125 115.785 ;
      END
   END dout0[397]
   PIN dout0[398]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.9825 115.65 444.1175 115.785 ;
      END
   END dout0[398]
   PIN dout0[399]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.6875 115.65 444.8225 115.785 ;
      END
   END dout0[399]
   PIN dout0[400]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  445.3925 115.65 445.5275 115.785 ;
      END
   END dout0[400]
   PIN dout0[401]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.0975 115.65 446.2325 115.785 ;
      END
   END dout0[401]
   PIN dout0[402]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.8025 115.65 446.9375 115.785 ;
      END
   END dout0[402]
   PIN dout0[403]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.5075 115.65 447.6425 115.785 ;
      END
   END dout0[403]
   PIN dout0[404]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  448.2125 115.65 448.3475 115.785 ;
      END
   END dout0[404]
   PIN dout0[405]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  448.9175 115.65 449.0525 115.785 ;
      END
   END dout0[405]
   PIN dout0[406]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.6225 115.65 449.7575 115.785 ;
      END
   END dout0[406]
   PIN dout0[407]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  450.3275 115.65 450.4625 115.785 ;
      END
   END dout0[407]
   PIN dout0[408]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  451.0325 115.65 451.1675 115.785 ;
      END
   END dout0[408]
   PIN dout0[409]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  451.7375 115.65 451.8725 115.785 ;
      END
   END dout0[409]
   PIN dout0[410]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.4425 115.65 452.5775 115.785 ;
      END
   END dout0[410]
   PIN dout0[411]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.1475 115.65 453.2825 115.785 ;
      END
   END dout0[411]
   PIN dout0[412]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.8525 115.65 453.9875 115.785 ;
      END
   END dout0[412]
   PIN dout0[413]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  454.5575 115.65 454.6925 115.785 ;
      END
   END dout0[413]
   PIN dout0[414]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.2625 115.65 455.3975 115.785 ;
      END
   END dout0[414]
   PIN dout0[415]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.9675 115.65 456.1025 115.785 ;
      END
   END dout0[415]
   PIN dout0[416]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  456.6725 115.65 456.8075 115.785 ;
      END
   END dout0[416]
   PIN dout0[417]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  457.3775 115.65 457.5125 115.785 ;
      END
   END dout0[417]
   PIN dout0[418]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.0825 115.65 458.2175 115.785 ;
      END
   END dout0[418]
   PIN dout0[419]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.7875 115.65 458.9225 115.785 ;
      END
   END dout0[419]
   PIN dout0[420]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  459.4925 115.65 459.6275 115.785 ;
      END
   END dout0[420]
   PIN dout0[421]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  460.1975 115.65 460.3325 115.785 ;
      END
   END dout0[421]
   PIN dout0[422]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  460.9025 115.65 461.0375 115.785 ;
      END
   END dout0[422]
   PIN dout0[423]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.6075 115.65 461.7425 115.785 ;
      END
   END dout0[423]
   PIN dout0[424]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  462.3125 115.65 462.4475 115.785 ;
      END
   END dout0[424]
   PIN dout0[425]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  463.0175 115.65 463.1525 115.785 ;
      END
   END dout0[425]
   PIN dout0[426]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  463.7225 115.65 463.8575 115.785 ;
      END
   END dout0[426]
   PIN dout0[427]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.4275 115.65 464.5625 115.785 ;
      END
   END dout0[427]
   PIN dout0[428]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  465.1325 115.65 465.2675 115.785 ;
      END
   END dout0[428]
   PIN dout0[429]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  465.8375 115.65 465.9725 115.785 ;
      END
   END dout0[429]
   PIN dout0[430]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  466.5425 115.65 466.6775 115.785 ;
      END
   END dout0[430]
   PIN dout0[431]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.2475 115.65 467.3825 115.785 ;
      END
   END dout0[431]
   PIN dout0[432]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.9525 115.65 468.0875 115.785 ;
      END
   END dout0[432]
   PIN dout0[433]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  468.6575 115.65 468.7925 115.785 ;
      END
   END dout0[433]
   PIN dout0[434]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  469.3625 115.65 469.4975 115.785 ;
      END
   END dout0[434]
   PIN dout0[435]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.0675 115.65 470.2025 115.785 ;
      END
   END dout0[435]
   PIN dout0[436]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.7725 115.65 470.9075 115.785 ;
      END
   END dout0[436]
   PIN dout0[437]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  471.4775 115.65 471.6125 115.785 ;
      END
   END dout0[437]
   PIN dout0[438]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.1825 115.65 472.3175 115.785 ;
      END
   END dout0[438]
   PIN dout0[439]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.8875 115.65 473.0225 115.785 ;
      END
   END dout0[439]
   PIN dout0[440]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  473.5925 115.65 473.7275 115.785 ;
      END
   END dout0[440]
   PIN dout0[441]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  474.2975 115.65 474.4325 115.785 ;
      END
   END dout0[441]
   PIN dout0[442]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.0025 115.65 475.1375 115.785 ;
      END
   END dout0[442]
   PIN dout0[443]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.7075 115.65 475.8425 115.785 ;
      END
   END dout0[443]
   PIN dout0[444]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  476.4125 115.65 476.5475 115.785 ;
      END
   END dout0[444]
   PIN dout0[445]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  477.1175 115.65 477.2525 115.785 ;
      END
   END dout0[445]
   PIN dout0[446]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  477.8225 115.65 477.9575 115.785 ;
      END
   END dout0[446]
   PIN dout0[447]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.5275 115.65 478.6625 115.785 ;
      END
   END dout0[447]
   PIN dout0[448]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  479.2325 115.65 479.3675 115.785 ;
      END
   END dout0[448]
   PIN dout0[449]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  479.9375 115.65 480.0725 115.785 ;
      END
   END dout0[449]
   PIN dout0[450]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  480.6425 115.65 480.7775 115.785 ;
      END
   END dout0[450]
   PIN dout0[451]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.3475 115.65 481.4825 115.785 ;
      END
   END dout0[451]
   PIN dout0[452]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.0525 115.65 482.1875 115.785 ;
      END
   END dout0[452]
   PIN dout0[453]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.7575 115.65 482.8925 115.785 ;
      END
   END dout0[453]
   PIN dout0[454]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  483.4625 115.65 483.5975 115.785 ;
      END
   END dout0[454]
   PIN dout0[455]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.1675 115.65 484.3025 115.785 ;
      END
   END dout0[455]
   PIN dout0[456]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.8725 115.65 485.0075 115.785 ;
      END
   END dout0[456]
   PIN dout0[457]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  485.5775 115.65 485.7125 115.785 ;
      END
   END dout0[457]
   PIN dout0[458]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.2825 115.65 486.4175 115.785 ;
      END
   END dout0[458]
   PIN dout0[459]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  486.9875 115.65 487.1225 115.785 ;
      END
   END dout0[459]
   PIN dout0[460]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.6925 115.65 487.8275 115.785 ;
      END
   END dout0[460]
   PIN dout0[461]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  488.3975 115.65 488.5325 115.785 ;
      END
   END dout0[461]
   PIN dout0[462]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.1025 115.65 489.2375 115.785 ;
      END
   END dout0[462]
   PIN dout0[463]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  489.8075 115.65 489.9425 115.785 ;
      END
   END dout0[463]
   PIN dout0[464]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  490.5125 115.65 490.6475 115.785 ;
      END
   END dout0[464]
   PIN dout0[465]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  491.2175 115.65 491.3525 115.785 ;
      END
   END dout0[465]
   PIN dout0[466]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  491.9225 115.65 492.0575 115.785 ;
      END
   END dout0[466]
   PIN dout0[467]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  492.6275 115.65 492.7625 115.785 ;
      END
   END dout0[467]
   PIN dout0[468]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  493.3325 115.65 493.4675 115.785 ;
      END
   END dout0[468]
   PIN dout0[469]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  494.0375 115.65 494.1725 115.785 ;
      END
   END dout0[469]
   PIN dout0[470]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  494.7425 115.65 494.8775 115.785 ;
      END
   END dout0[470]
   PIN dout0[471]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  495.4475 115.65 495.5825 115.785 ;
      END
   END dout0[471]
   PIN dout0[472]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  496.1525 115.65 496.2875 115.785 ;
      END
   END dout0[472]
   PIN dout0[473]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  496.8575 115.65 496.9925 115.785 ;
      END
   END dout0[473]
   PIN dout0[474]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  497.5625 115.65 497.6975 115.785 ;
      END
   END dout0[474]
   PIN dout0[475]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.2675 115.65 498.4025 115.785 ;
      END
   END dout0[475]
   PIN dout0[476]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.9725 115.65 499.1075 115.785 ;
      END
   END dout0[476]
   PIN dout0[477]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  499.6775 115.65 499.8125 115.785 ;
      END
   END dout0[477]
   PIN dout0[478]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  500.3825 115.65 500.5175 115.785 ;
      END
   END dout0[478]
   PIN dout0[479]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.0875 115.65 501.2225 115.785 ;
      END
   END dout0[479]
   PIN dout0[480]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.7925 115.65 501.9275 115.785 ;
      END
   END dout0[480]
   PIN dout0[481]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  502.4975 115.65 502.6325 115.785 ;
      END
   END dout0[481]
   PIN dout0[482]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  503.2025 115.65 503.3375 115.785 ;
      END
   END dout0[482]
   PIN dout0[483]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  503.9075 115.65 504.0425 115.785 ;
      END
   END dout0[483]
   PIN dout0[484]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.6125 115.65 504.7475 115.785 ;
      END
   END dout0[484]
   PIN dout0[485]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  505.3175 115.65 505.4525 115.785 ;
      END
   END dout0[485]
   PIN dout0[486]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  506.0225 115.65 506.1575 115.785 ;
      END
   END dout0[486]
   PIN dout0[487]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  506.7275 115.65 506.8625 115.785 ;
      END
   END dout0[487]
   PIN dout0[488]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.4325 115.65 507.5675 115.785 ;
      END
   END dout0[488]
   PIN dout0[489]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  508.1375 115.65 508.2725 115.785 ;
      END
   END dout0[489]
   PIN dout0[490]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  508.8425 115.65 508.9775 115.785 ;
      END
   END dout0[490]
   PIN dout0[491]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  509.5475 115.65 509.6825 115.785 ;
      END
   END dout0[491]
   PIN dout0[492]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.2525 115.65 510.3875 115.785 ;
      END
   END dout0[492]
   PIN dout0[493]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.9575 115.65 511.0925 115.785 ;
      END
   END dout0[493]
   PIN dout0[494]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  511.6625 115.65 511.7975 115.785 ;
      END
   END dout0[494]
   PIN dout0[495]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  512.3675 115.65 512.5025 115.785 ;
      END
   END dout0[495]
   PIN dout0[496]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  513.0725 115.65 513.2075 115.785 ;
      END
   END dout0[496]
   PIN dout0[497]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  513.7775 115.65 513.9125 115.785 ;
      END
   END dout0[497]
   PIN dout0[498]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.4825 115.65 514.6175 115.785 ;
      END
   END dout0[498]
   PIN dout0[499]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.1875 115.65 515.3225 115.785 ;
      END
   END dout0[499]
   PIN dout0[500]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  515.8925 115.65 516.0275 115.785 ;
      END
   END dout0[500]
   PIN dout0[501]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  516.5975 115.65 516.7325 115.785 ;
      END
   END dout0[501]
   PIN dout0[502]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  517.3025 115.65 517.4375 115.785 ;
      END
   END dout0[502]
   PIN dout0[503]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.0075 115.65 518.1425 115.785 ;
      END
   END dout0[503]
   PIN dout0[504]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.7125 115.65 518.8475 115.785 ;
      END
   END dout0[504]
   PIN dout0[505]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  519.4175 115.65 519.5525 115.785 ;
      END
   END dout0[505]
   PIN dout0[506]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  520.1225 115.65 520.2575 115.785 ;
      END
   END dout0[506]
   PIN dout0[507]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  520.8275 115.65 520.9625 115.785 ;
      END
   END dout0[507]
   PIN dout0[508]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.5325 115.65 521.6675 115.785 ;
      END
   END dout0[508]
   PIN dout0[509]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  522.2375 115.65 522.3725 115.785 ;
      END
   END dout0[509]
   PIN dout0[510]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  522.9425 115.65 523.0775 115.785 ;
      END
   END dout0[510]
   PIN dout0[511]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  523.6475 115.65 523.7825 115.785 ;
      END
   END dout0[511]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  1.4 216.72 1592.5 217.42 ;
         LAYER metal3 ;
         RECT  1.4 1.4 1592.5 2.1 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 217.42 ;
         LAYER metal4 ;
         RECT  1591.8 1.4 1592.5 217.42 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  1593.2 0.0 1593.9 218.82 ;
         LAYER metal3 ;
         RECT  0.0 218.12 1593.9 218.82 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 218.82 ;
         LAYER metal3 ;
         RECT  0.0 0.0 1593.9 0.7 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 1593.76 218.68 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 1593.76 218.68 ;
   LAYER  metal3 ;
      RECT  0.14 4.0975 126.485 4.5125 ;
      RECT  126.9 4.0975 129.345 4.5125 ;
      RECT  129.76 4.0975 132.205 4.5125 ;
      RECT  132.62 4.0975 135.065 4.5125 ;
      RECT  135.48 4.0975 137.925 4.5125 ;
      RECT  138.34 4.0975 140.785 4.5125 ;
      RECT  141.2 4.0975 143.645 4.5125 ;
      RECT  144.06 4.0975 146.505 4.5125 ;
      RECT  146.92 4.0975 149.365 4.5125 ;
      RECT  149.78 4.0975 152.225 4.5125 ;
      RECT  152.64 4.0975 155.085 4.5125 ;
      RECT  155.5 4.0975 157.945 4.5125 ;
      RECT  158.36 4.0975 160.805 4.5125 ;
      RECT  161.22 4.0975 163.665 4.5125 ;
      RECT  164.08 4.0975 166.525 4.5125 ;
      RECT  166.94 4.0975 169.385 4.5125 ;
      RECT  169.8 4.0975 172.245 4.5125 ;
      RECT  172.66 4.0975 175.105 4.5125 ;
      RECT  175.52 4.0975 177.965 4.5125 ;
      RECT  178.38 4.0975 180.825 4.5125 ;
      RECT  181.24 4.0975 183.685 4.5125 ;
      RECT  184.1 4.0975 186.545 4.5125 ;
      RECT  186.96 4.0975 189.405 4.5125 ;
      RECT  189.82 4.0975 192.265 4.5125 ;
      RECT  192.68 4.0975 195.125 4.5125 ;
      RECT  195.54 4.0975 197.985 4.5125 ;
      RECT  198.4 4.0975 200.845 4.5125 ;
      RECT  201.26 4.0975 203.705 4.5125 ;
      RECT  204.12 4.0975 206.565 4.5125 ;
      RECT  206.98 4.0975 209.425 4.5125 ;
      RECT  209.84 4.0975 212.285 4.5125 ;
      RECT  212.7 4.0975 215.145 4.5125 ;
      RECT  215.56 4.0975 218.005 4.5125 ;
      RECT  218.42 4.0975 220.865 4.5125 ;
      RECT  221.28 4.0975 223.725 4.5125 ;
      RECT  224.14 4.0975 226.585 4.5125 ;
      RECT  227.0 4.0975 229.445 4.5125 ;
      RECT  229.86 4.0975 232.305 4.5125 ;
      RECT  232.72 4.0975 235.165 4.5125 ;
      RECT  235.58 4.0975 238.025 4.5125 ;
      RECT  238.44 4.0975 240.885 4.5125 ;
      RECT  241.3 4.0975 243.745 4.5125 ;
      RECT  244.16 4.0975 246.605 4.5125 ;
      RECT  247.02 4.0975 249.465 4.5125 ;
      RECT  249.88 4.0975 252.325 4.5125 ;
      RECT  252.74 4.0975 255.185 4.5125 ;
      RECT  255.6 4.0975 258.045 4.5125 ;
      RECT  258.46 4.0975 260.905 4.5125 ;
      RECT  261.32 4.0975 263.765 4.5125 ;
      RECT  264.18 4.0975 266.625 4.5125 ;
      RECT  267.04 4.0975 269.485 4.5125 ;
      RECT  269.9 4.0975 272.345 4.5125 ;
      RECT  272.76 4.0975 275.205 4.5125 ;
      RECT  275.62 4.0975 278.065 4.5125 ;
      RECT  278.48 4.0975 280.925 4.5125 ;
      RECT  281.34 4.0975 283.785 4.5125 ;
      RECT  284.2 4.0975 286.645 4.5125 ;
      RECT  287.06 4.0975 289.505 4.5125 ;
      RECT  289.92 4.0975 292.365 4.5125 ;
      RECT  292.78 4.0975 295.225 4.5125 ;
      RECT  295.64 4.0975 298.085 4.5125 ;
      RECT  298.5 4.0975 300.945 4.5125 ;
      RECT  301.36 4.0975 303.805 4.5125 ;
      RECT  304.22 4.0975 306.665 4.5125 ;
      RECT  307.08 4.0975 309.525 4.5125 ;
      RECT  309.94 4.0975 312.385 4.5125 ;
      RECT  312.8 4.0975 315.245 4.5125 ;
      RECT  315.66 4.0975 318.105 4.5125 ;
      RECT  318.52 4.0975 320.965 4.5125 ;
      RECT  321.38 4.0975 323.825 4.5125 ;
      RECT  324.24 4.0975 326.685 4.5125 ;
      RECT  327.1 4.0975 329.545 4.5125 ;
      RECT  329.96 4.0975 332.405 4.5125 ;
      RECT  332.82 4.0975 335.265 4.5125 ;
      RECT  335.68 4.0975 338.125 4.5125 ;
      RECT  338.54 4.0975 340.985 4.5125 ;
      RECT  341.4 4.0975 343.845 4.5125 ;
      RECT  344.26 4.0975 346.705 4.5125 ;
      RECT  347.12 4.0975 349.565 4.5125 ;
      RECT  349.98 4.0975 352.425 4.5125 ;
      RECT  352.84 4.0975 355.285 4.5125 ;
      RECT  355.7 4.0975 358.145 4.5125 ;
      RECT  358.56 4.0975 361.005 4.5125 ;
      RECT  361.42 4.0975 363.865 4.5125 ;
      RECT  364.28 4.0975 366.725 4.5125 ;
      RECT  367.14 4.0975 369.585 4.5125 ;
      RECT  370.0 4.0975 372.445 4.5125 ;
      RECT  372.86 4.0975 375.305 4.5125 ;
      RECT  375.72 4.0975 378.165 4.5125 ;
      RECT  378.58 4.0975 381.025 4.5125 ;
      RECT  381.44 4.0975 383.885 4.5125 ;
      RECT  384.3 4.0975 386.745 4.5125 ;
      RECT  387.16 4.0975 389.605 4.5125 ;
      RECT  390.02 4.0975 392.465 4.5125 ;
      RECT  392.88 4.0975 395.325 4.5125 ;
      RECT  395.74 4.0975 398.185 4.5125 ;
      RECT  398.6 4.0975 401.045 4.5125 ;
      RECT  401.46 4.0975 403.905 4.5125 ;
      RECT  404.32 4.0975 406.765 4.5125 ;
      RECT  407.18 4.0975 409.625 4.5125 ;
      RECT  410.04 4.0975 412.485 4.5125 ;
      RECT  412.9 4.0975 415.345 4.5125 ;
      RECT  415.76 4.0975 418.205 4.5125 ;
      RECT  418.62 4.0975 421.065 4.5125 ;
      RECT  421.48 4.0975 423.925 4.5125 ;
      RECT  424.34 4.0975 426.785 4.5125 ;
      RECT  427.2 4.0975 429.645 4.5125 ;
      RECT  430.06 4.0975 432.505 4.5125 ;
      RECT  432.92 4.0975 435.365 4.5125 ;
      RECT  435.78 4.0975 438.225 4.5125 ;
      RECT  438.64 4.0975 441.085 4.5125 ;
      RECT  441.5 4.0975 443.945 4.5125 ;
      RECT  444.36 4.0975 446.805 4.5125 ;
      RECT  447.22 4.0975 449.665 4.5125 ;
      RECT  450.08 4.0975 452.525 4.5125 ;
      RECT  452.94 4.0975 455.385 4.5125 ;
      RECT  455.8 4.0975 458.245 4.5125 ;
      RECT  458.66 4.0975 461.105 4.5125 ;
      RECT  461.52 4.0975 463.965 4.5125 ;
      RECT  464.38 4.0975 466.825 4.5125 ;
      RECT  467.24 4.0975 469.685 4.5125 ;
      RECT  470.1 4.0975 472.545 4.5125 ;
      RECT  472.96 4.0975 475.405 4.5125 ;
      RECT  475.82 4.0975 478.265 4.5125 ;
      RECT  478.68 4.0975 481.125 4.5125 ;
      RECT  481.54 4.0975 483.985 4.5125 ;
      RECT  484.4 4.0975 486.845 4.5125 ;
      RECT  487.26 4.0975 489.705 4.5125 ;
      RECT  490.12 4.0975 492.565 4.5125 ;
      RECT  492.98 4.0975 495.425 4.5125 ;
      RECT  495.84 4.0975 498.285 4.5125 ;
      RECT  498.7 4.0975 501.145 4.5125 ;
      RECT  501.56 4.0975 504.005 4.5125 ;
      RECT  504.42 4.0975 506.865 4.5125 ;
      RECT  507.28 4.0975 509.725 4.5125 ;
      RECT  510.14 4.0975 512.585 4.5125 ;
      RECT  513.0 4.0975 515.445 4.5125 ;
      RECT  515.86 4.0975 518.305 4.5125 ;
      RECT  518.72 4.0975 521.165 4.5125 ;
      RECT  521.58 4.0975 524.025 4.5125 ;
      RECT  524.44 4.0975 526.885 4.5125 ;
      RECT  527.3 4.0975 529.745 4.5125 ;
      RECT  530.16 4.0975 532.605 4.5125 ;
      RECT  533.02 4.0975 535.465 4.5125 ;
      RECT  535.88 4.0975 538.325 4.5125 ;
      RECT  538.74 4.0975 541.185 4.5125 ;
      RECT  541.6 4.0975 544.045 4.5125 ;
      RECT  544.46 4.0975 546.905 4.5125 ;
      RECT  547.32 4.0975 549.765 4.5125 ;
      RECT  550.18 4.0975 552.625 4.5125 ;
      RECT  553.04 4.0975 555.485 4.5125 ;
      RECT  555.9 4.0975 558.345 4.5125 ;
      RECT  558.76 4.0975 561.205 4.5125 ;
      RECT  561.62 4.0975 564.065 4.5125 ;
      RECT  564.48 4.0975 566.925 4.5125 ;
      RECT  567.34 4.0975 569.785 4.5125 ;
      RECT  570.2 4.0975 572.645 4.5125 ;
      RECT  573.06 4.0975 575.505 4.5125 ;
      RECT  575.92 4.0975 578.365 4.5125 ;
      RECT  578.78 4.0975 581.225 4.5125 ;
      RECT  581.64 4.0975 584.085 4.5125 ;
      RECT  584.5 4.0975 586.945 4.5125 ;
      RECT  587.36 4.0975 589.805 4.5125 ;
      RECT  590.22 4.0975 592.665 4.5125 ;
      RECT  593.08 4.0975 595.525 4.5125 ;
      RECT  595.94 4.0975 598.385 4.5125 ;
      RECT  598.8 4.0975 601.245 4.5125 ;
      RECT  601.66 4.0975 604.105 4.5125 ;
      RECT  604.52 4.0975 606.965 4.5125 ;
      RECT  607.38 4.0975 609.825 4.5125 ;
      RECT  610.24 4.0975 612.685 4.5125 ;
      RECT  613.1 4.0975 615.545 4.5125 ;
      RECT  615.96 4.0975 618.405 4.5125 ;
      RECT  618.82 4.0975 621.265 4.5125 ;
      RECT  621.68 4.0975 624.125 4.5125 ;
      RECT  624.54 4.0975 626.985 4.5125 ;
      RECT  627.4 4.0975 629.845 4.5125 ;
      RECT  630.26 4.0975 632.705 4.5125 ;
      RECT  633.12 4.0975 635.565 4.5125 ;
      RECT  635.98 4.0975 638.425 4.5125 ;
      RECT  638.84 4.0975 641.285 4.5125 ;
      RECT  641.7 4.0975 644.145 4.5125 ;
      RECT  644.56 4.0975 647.005 4.5125 ;
      RECT  647.42 4.0975 649.865 4.5125 ;
      RECT  650.28 4.0975 652.725 4.5125 ;
      RECT  653.14 4.0975 655.585 4.5125 ;
      RECT  656.0 4.0975 658.445 4.5125 ;
      RECT  658.86 4.0975 661.305 4.5125 ;
      RECT  661.72 4.0975 664.165 4.5125 ;
      RECT  664.58 4.0975 667.025 4.5125 ;
      RECT  667.44 4.0975 669.885 4.5125 ;
      RECT  670.3 4.0975 672.745 4.5125 ;
      RECT  673.16 4.0975 675.605 4.5125 ;
      RECT  676.02 4.0975 678.465 4.5125 ;
      RECT  678.88 4.0975 681.325 4.5125 ;
      RECT  681.74 4.0975 684.185 4.5125 ;
      RECT  684.6 4.0975 687.045 4.5125 ;
      RECT  687.46 4.0975 689.905 4.5125 ;
      RECT  690.32 4.0975 692.765 4.5125 ;
      RECT  693.18 4.0975 695.625 4.5125 ;
      RECT  696.04 4.0975 698.485 4.5125 ;
      RECT  698.9 4.0975 701.345 4.5125 ;
      RECT  701.76 4.0975 704.205 4.5125 ;
      RECT  704.62 4.0975 707.065 4.5125 ;
      RECT  707.48 4.0975 709.925 4.5125 ;
      RECT  710.34 4.0975 712.785 4.5125 ;
      RECT  713.2 4.0975 715.645 4.5125 ;
      RECT  716.06 4.0975 718.505 4.5125 ;
      RECT  718.92 4.0975 721.365 4.5125 ;
      RECT  721.78 4.0975 724.225 4.5125 ;
      RECT  724.64 4.0975 727.085 4.5125 ;
      RECT  727.5 4.0975 729.945 4.5125 ;
      RECT  730.36 4.0975 732.805 4.5125 ;
      RECT  733.22 4.0975 735.665 4.5125 ;
      RECT  736.08 4.0975 738.525 4.5125 ;
      RECT  738.94 4.0975 741.385 4.5125 ;
      RECT  741.8 4.0975 744.245 4.5125 ;
      RECT  744.66 4.0975 747.105 4.5125 ;
      RECT  747.52 4.0975 749.965 4.5125 ;
      RECT  750.38 4.0975 752.825 4.5125 ;
      RECT  753.24 4.0975 755.685 4.5125 ;
      RECT  756.1 4.0975 758.545 4.5125 ;
      RECT  758.96 4.0975 761.405 4.5125 ;
      RECT  761.82 4.0975 764.265 4.5125 ;
      RECT  764.68 4.0975 767.125 4.5125 ;
      RECT  767.54 4.0975 769.985 4.5125 ;
      RECT  770.4 4.0975 772.845 4.5125 ;
      RECT  773.26 4.0975 775.705 4.5125 ;
      RECT  776.12 4.0975 778.565 4.5125 ;
      RECT  778.98 4.0975 781.425 4.5125 ;
      RECT  781.84 4.0975 784.285 4.5125 ;
      RECT  784.7 4.0975 787.145 4.5125 ;
      RECT  787.56 4.0975 790.005 4.5125 ;
      RECT  790.42 4.0975 792.865 4.5125 ;
      RECT  793.28 4.0975 795.725 4.5125 ;
      RECT  796.14 4.0975 798.585 4.5125 ;
      RECT  799.0 4.0975 801.445 4.5125 ;
      RECT  801.86 4.0975 804.305 4.5125 ;
      RECT  804.72 4.0975 807.165 4.5125 ;
      RECT  807.58 4.0975 810.025 4.5125 ;
      RECT  810.44 4.0975 812.885 4.5125 ;
      RECT  813.3 4.0975 815.745 4.5125 ;
      RECT  816.16 4.0975 818.605 4.5125 ;
      RECT  819.02 4.0975 821.465 4.5125 ;
      RECT  821.88 4.0975 824.325 4.5125 ;
      RECT  824.74 4.0975 827.185 4.5125 ;
      RECT  827.6 4.0975 830.045 4.5125 ;
      RECT  830.46 4.0975 832.905 4.5125 ;
      RECT  833.32 4.0975 835.765 4.5125 ;
      RECT  836.18 4.0975 838.625 4.5125 ;
      RECT  839.04 4.0975 841.485 4.5125 ;
      RECT  841.9 4.0975 844.345 4.5125 ;
      RECT  844.76 4.0975 847.205 4.5125 ;
      RECT  847.62 4.0975 850.065 4.5125 ;
      RECT  850.48 4.0975 852.925 4.5125 ;
      RECT  853.34 4.0975 855.785 4.5125 ;
      RECT  856.2 4.0975 858.645 4.5125 ;
      RECT  859.06 4.0975 861.505 4.5125 ;
      RECT  861.92 4.0975 864.365 4.5125 ;
      RECT  864.78 4.0975 867.225 4.5125 ;
      RECT  867.64 4.0975 870.085 4.5125 ;
      RECT  870.5 4.0975 872.945 4.5125 ;
      RECT  873.36 4.0975 875.805 4.5125 ;
      RECT  876.22 4.0975 878.665 4.5125 ;
      RECT  879.08 4.0975 881.525 4.5125 ;
      RECT  881.94 4.0975 884.385 4.5125 ;
      RECT  884.8 4.0975 887.245 4.5125 ;
      RECT  887.66 4.0975 890.105 4.5125 ;
      RECT  890.52 4.0975 892.965 4.5125 ;
      RECT  893.38 4.0975 895.825 4.5125 ;
      RECT  896.24 4.0975 898.685 4.5125 ;
      RECT  899.1 4.0975 901.545 4.5125 ;
      RECT  901.96 4.0975 904.405 4.5125 ;
      RECT  904.82 4.0975 907.265 4.5125 ;
      RECT  907.68 4.0975 910.125 4.5125 ;
      RECT  910.54 4.0975 912.985 4.5125 ;
      RECT  913.4 4.0975 915.845 4.5125 ;
      RECT  916.26 4.0975 918.705 4.5125 ;
      RECT  919.12 4.0975 921.565 4.5125 ;
      RECT  921.98 4.0975 924.425 4.5125 ;
      RECT  924.84 4.0975 927.285 4.5125 ;
      RECT  927.7 4.0975 930.145 4.5125 ;
      RECT  930.56 4.0975 933.005 4.5125 ;
      RECT  933.42 4.0975 935.865 4.5125 ;
      RECT  936.28 4.0975 938.725 4.5125 ;
      RECT  939.14 4.0975 941.585 4.5125 ;
      RECT  942.0 4.0975 944.445 4.5125 ;
      RECT  944.86 4.0975 947.305 4.5125 ;
      RECT  947.72 4.0975 950.165 4.5125 ;
      RECT  950.58 4.0975 953.025 4.5125 ;
      RECT  953.44 4.0975 955.885 4.5125 ;
      RECT  956.3 4.0975 958.745 4.5125 ;
      RECT  959.16 4.0975 961.605 4.5125 ;
      RECT  962.02 4.0975 964.465 4.5125 ;
      RECT  964.88 4.0975 967.325 4.5125 ;
      RECT  967.74 4.0975 970.185 4.5125 ;
      RECT  970.6 4.0975 973.045 4.5125 ;
      RECT  973.46 4.0975 975.905 4.5125 ;
      RECT  976.32 4.0975 978.765 4.5125 ;
      RECT  979.18 4.0975 981.625 4.5125 ;
      RECT  982.04 4.0975 984.485 4.5125 ;
      RECT  984.9 4.0975 987.345 4.5125 ;
      RECT  987.76 4.0975 990.205 4.5125 ;
      RECT  990.62 4.0975 993.065 4.5125 ;
      RECT  993.48 4.0975 995.925 4.5125 ;
      RECT  996.34 4.0975 998.785 4.5125 ;
      RECT  999.2 4.0975 1001.645 4.5125 ;
      RECT  1002.06 4.0975 1004.505 4.5125 ;
      RECT  1004.92 4.0975 1007.365 4.5125 ;
      RECT  1007.78 4.0975 1010.225 4.5125 ;
      RECT  1010.64 4.0975 1013.085 4.5125 ;
      RECT  1013.5 4.0975 1015.945 4.5125 ;
      RECT  1016.36 4.0975 1018.805 4.5125 ;
      RECT  1019.22 4.0975 1021.665 4.5125 ;
      RECT  1022.08 4.0975 1024.525 4.5125 ;
      RECT  1024.94 4.0975 1027.385 4.5125 ;
      RECT  1027.8 4.0975 1030.245 4.5125 ;
      RECT  1030.66 4.0975 1033.105 4.5125 ;
      RECT  1033.52 4.0975 1035.965 4.5125 ;
      RECT  1036.38 4.0975 1038.825 4.5125 ;
      RECT  1039.24 4.0975 1041.685 4.5125 ;
      RECT  1042.1 4.0975 1044.545 4.5125 ;
      RECT  1044.96 4.0975 1047.405 4.5125 ;
      RECT  1047.82 4.0975 1050.265 4.5125 ;
      RECT  1050.68 4.0975 1053.125 4.5125 ;
      RECT  1053.54 4.0975 1055.985 4.5125 ;
      RECT  1056.4 4.0975 1058.845 4.5125 ;
      RECT  1059.26 4.0975 1061.705 4.5125 ;
      RECT  1062.12 4.0975 1064.565 4.5125 ;
      RECT  1064.98 4.0975 1067.425 4.5125 ;
      RECT  1067.84 4.0975 1070.285 4.5125 ;
      RECT  1070.7 4.0975 1073.145 4.5125 ;
      RECT  1073.56 4.0975 1076.005 4.5125 ;
      RECT  1076.42 4.0975 1078.865 4.5125 ;
      RECT  1079.28 4.0975 1081.725 4.5125 ;
      RECT  1082.14 4.0975 1084.585 4.5125 ;
      RECT  1085.0 4.0975 1087.445 4.5125 ;
      RECT  1087.86 4.0975 1090.305 4.5125 ;
      RECT  1090.72 4.0975 1093.165 4.5125 ;
      RECT  1093.58 4.0975 1096.025 4.5125 ;
      RECT  1096.44 4.0975 1098.885 4.5125 ;
      RECT  1099.3 4.0975 1101.745 4.5125 ;
      RECT  1102.16 4.0975 1104.605 4.5125 ;
      RECT  1105.02 4.0975 1107.465 4.5125 ;
      RECT  1107.88 4.0975 1110.325 4.5125 ;
      RECT  1110.74 4.0975 1113.185 4.5125 ;
      RECT  1113.6 4.0975 1116.045 4.5125 ;
      RECT  1116.46 4.0975 1118.905 4.5125 ;
      RECT  1119.32 4.0975 1121.765 4.5125 ;
      RECT  1122.18 4.0975 1124.625 4.5125 ;
      RECT  1125.04 4.0975 1127.485 4.5125 ;
      RECT  1127.9 4.0975 1130.345 4.5125 ;
      RECT  1130.76 4.0975 1133.205 4.5125 ;
      RECT  1133.62 4.0975 1136.065 4.5125 ;
      RECT  1136.48 4.0975 1138.925 4.5125 ;
      RECT  1139.34 4.0975 1141.785 4.5125 ;
      RECT  1142.2 4.0975 1144.645 4.5125 ;
      RECT  1145.06 4.0975 1147.505 4.5125 ;
      RECT  1147.92 4.0975 1150.365 4.5125 ;
      RECT  1150.78 4.0975 1153.225 4.5125 ;
      RECT  1153.64 4.0975 1156.085 4.5125 ;
      RECT  1156.5 4.0975 1158.945 4.5125 ;
      RECT  1159.36 4.0975 1161.805 4.5125 ;
      RECT  1162.22 4.0975 1164.665 4.5125 ;
      RECT  1165.08 4.0975 1167.525 4.5125 ;
      RECT  1167.94 4.0975 1170.385 4.5125 ;
      RECT  1170.8 4.0975 1173.245 4.5125 ;
      RECT  1173.66 4.0975 1176.105 4.5125 ;
      RECT  1176.52 4.0975 1178.965 4.5125 ;
      RECT  1179.38 4.0975 1181.825 4.5125 ;
      RECT  1182.24 4.0975 1184.685 4.5125 ;
      RECT  1185.1 4.0975 1187.545 4.5125 ;
      RECT  1187.96 4.0975 1190.405 4.5125 ;
      RECT  1190.82 4.0975 1193.265 4.5125 ;
      RECT  1193.68 4.0975 1196.125 4.5125 ;
      RECT  1196.54 4.0975 1198.985 4.5125 ;
      RECT  1199.4 4.0975 1201.845 4.5125 ;
      RECT  1202.26 4.0975 1204.705 4.5125 ;
      RECT  1205.12 4.0975 1207.565 4.5125 ;
      RECT  1207.98 4.0975 1210.425 4.5125 ;
      RECT  1210.84 4.0975 1213.285 4.5125 ;
      RECT  1213.7 4.0975 1216.145 4.5125 ;
      RECT  1216.56 4.0975 1219.005 4.5125 ;
      RECT  1219.42 4.0975 1221.865 4.5125 ;
      RECT  1222.28 4.0975 1224.725 4.5125 ;
      RECT  1225.14 4.0975 1227.585 4.5125 ;
      RECT  1228.0 4.0975 1230.445 4.5125 ;
      RECT  1230.86 4.0975 1233.305 4.5125 ;
      RECT  1233.72 4.0975 1236.165 4.5125 ;
      RECT  1236.58 4.0975 1239.025 4.5125 ;
      RECT  1239.44 4.0975 1241.885 4.5125 ;
      RECT  1242.3 4.0975 1244.745 4.5125 ;
      RECT  1245.16 4.0975 1247.605 4.5125 ;
      RECT  1248.02 4.0975 1250.465 4.5125 ;
      RECT  1250.88 4.0975 1253.325 4.5125 ;
      RECT  1253.74 4.0975 1256.185 4.5125 ;
      RECT  1256.6 4.0975 1259.045 4.5125 ;
      RECT  1259.46 4.0975 1261.905 4.5125 ;
      RECT  1262.32 4.0975 1264.765 4.5125 ;
      RECT  1265.18 4.0975 1267.625 4.5125 ;
      RECT  1268.04 4.0975 1270.485 4.5125 ;
      RECT  1270.9 4.0975 1273.345 4.5125 ;
      RECT  1273.76 4.0975 1276.205 4.5125 ;
      RECT  1276.62 4.0975 1279.065 4.5125 ;
      RECT  1279.48 4.0975 1281.925 4.5125 ;
      RECT  1282.34 4.0975 1284.785 4.5125 ;
      RECT  1285.2 4.0975 1287.645 4.5125 ;
      RECT  1288.06 4.0975 1290.505 4.5125 ;
      RECT  1290.92 4.0975 1293.365 4.5125 ;
      RECT  1293.78 4.0975 1296.225 4.5125 ;
      RECT  1296.64 4.0975 1299.085 4.5125 ;
      RECT  1299.5 4.0975 1301.945 4.5125 ;
      RECT  1302.36 4.0975 1304.805 4.5125 ;
      RECT  1305.22 4.0975 1307.665 4.5125 ;
      RECT  1308.08 4.0975 1310.525 4.5125 ;
      RECT  1310.94 4.0975 1313.385 4.5125 ;
      RECT  1313.8 4.0975 1316.245 4.5125 ;
      RECT  1316.66 4.0975 1319.105 4.5125 ;
      RECT  1319.52 4.0975 1321.965 4.5125 ;
      RECT  1322.38 4.0975 1324.825 4.5125 ;
      RECT  1325.24 4.0975 1327.685 4.5125 ;
      RECT  1328.1 4.0975 1330.545 4.5125 ;
      RECT  1330.96 4.0975 1333.405 4.5125 ;
      RECT  1333.82 4.0975 1336.265 4.5125 ;
      RECT  1336.68 4.0975 1339.125 4.5125 ;
      RECT  1339.54 4.0975 1341.985 4.5125 ;
      RECT  1342.4 4.0975 1344.845 4.5125 ;
      RECT  1345.26 4.0975 1347.705 4.5125 ;
      RECT  1348.12 4.0975 1350.565 4.5125 ;
      RECT  1350.98 4.0975 1353.425 4.5125 ;
      RECT  1353.84 4.0975 1356.285 4.5125 ;
      RECT  1356.7 4.0975 1359.145 4.5125 ;
      RECT  1359.56 4.0975 1362.005 4.5125 ;
      RECT  1362.42 4.0975 1364.865 4.5125 ;
      RECT  1365.28 4.0975 1367.725 4.5125 ;
      RECT  1368.14 4.0975 1370.585 4.5125 ;
      RECT  1371.0 4.0975 1373.445 4.5125 ;
      RECT  1373.86 4.0975 1376.305 4.5125 ;
      RECT  1376.72 4.0975 1379.165 4.5125 ;
      RECT  1379.58 4.0975 1382.025 4.5125 ;
      RECT  1382.44 4.0975 1384.885 4.5125 ;
      RECT  1385.3 4.0975 1387.745 4.5125 ;
      RECT  1388.16 4.0975 1390.605 4.5125 ;
      RECT  1391.02 4.0975 1393.465 4.5125 ;
      RECT  1393.88 4.0975 1396.325 4.5125 ;
      RECT  1396.74 4.0975 1399.185 4.5125 ;
      RECT  1399.6 4.0975 1402.045 4.5125 ;
      RECT  1402.46 4.0975 1404.905 4.5125 ;
      RECT  1405.32 4.0975 1407.765 4.5125 ;
      RECT  1408.18 4.0975 1410.625 4.5125 ;
      RECT  1411.04 4.0975 1413.485 4.5125 ;
      RECT  1413.9 4.0975 1416.345 4.5125 ;
      RECT  1416.76 4.0975 1419.205 4.5125 ;
      RECT  1419.62 4.0975 1422.065 4.5125 ;
      RECT  1422.48 4.0975 1424.925 4.5125 ;
      RECT  1425.34 4.0975 1427.785 4.5125 ;
      RECT  1428.2 4.0975 1430.645 4.5125 ;
      RECT  1431.06 4.0975 1433.505 4.5125 ;
      RECT  1433.92 4.0975 1436.365 4.5125 ;
      RECT  1436.78 4.0975 1439.225 4.5125 ;
      RECT  1439.64 4.0975 1442.085 4.5125 ;
      RECT  1442.5 4.0975 1444.945 4.5125 ;
      RECT  1445.36 4.0975 1447.805 4.5125 ;
      RECT  1448.22 4.0975 1450.665 4.5125 ;
      RECT  1451.08 4.0975 1453.525 4.5125 ;
      RECT  1453.94 4.0975 1456.385 4.5125 ;
      RECT  1456.8 4.0975 1459.245 4.5125 ;
      RECT  1459.66 4.0975 1462.105 4.5125 ;
      RECT  1462.52 4.0975 1464.965 4.5125 ;
      RECT  1465.38 4.0975 1467.825 4.5125 ;
      RECT  1468.24 4.0975 1470.685 4.5125 ;
      RECT  1471.1 4.0975 1473.545 4.5125 ;
      RECT  1473.96 4.0975 1476.405 4.5125 ;
      RECT  1476.82 4.0975 1479.265 4.5125 ;
      RECT  1479.68 4.0975 1482.125 4.5125 ;
      RECT  1482.54 4.0975 1484.985 4.5125 ;
      RECT  1485.4 4.0975 1487.845 4.5125 ;
      RECT  1488.26 4.0975 1490.705 4.5125 ;
      RECT  1491.12 4.0975 1493.565 4.5125 ;
      RECT  1493.98 4.0975 1496.425 4.5125 ;
      RECT  1496.84 4.0975 1499.285 4.5125 ;
      RECT  1499.7 4.0975 1502.145 4.5125 ;
      RECT  1502.56 4.0975 1505.005 4.5125 ;
      RECT  1505.42 4.0975 1507.865 4.5125 ;
      RECT  1508.28 4.0975 1510.725 4.5125 ;
      RECT  1511.14 4.0975 1513.585 4.5125 ;
      RECT  1514.0 4.0975 1516.445 4.5125 ;
      RECT  1516.86 4.0975 1519.305 4.5125 ;
      RECT  1519.72 4.0975 1522.165 4.5125 ;
      RECT  1522.58 4.0975 1525.025 4.5125 ;
      RECT  1525.44 4.0975 1527.885 4.5125 ;
      RECT  1528.3 4.0975 1530.745 4.5125 ;
      RECT  1531.16 4.0975 1533.605 4.5125 ;
      RECT  1534.02 4.0975 1536.465 4.5125 ;
      RECT  1536.88 4.0975 1539.325 4.5125 ;
      RECT  1539.74 4.0975 1542.185 4.5125 ;
      RECT  1542.6 4.0975 1545.045 4.5125 ;
      RECT  1545.46 4.0975 1547.905 4.5125 ;
      RECT  1548.32 4.0975 1550.765 4.5125 ;
      RECT  1551.18 4.0975 1553.625 4.5125 ;
      RECT  1554.04 4.0975 1556.485 4.5125 ;
      RECT  1556.9 4.0975 1559.345 4.5125 ;
      RECT  1559.76 4.0975 1562.205 4.5125 ;
      RECT  1562.62 4.0975 1565.065 4.5125 ;
      RECT  1565.48 4.0975 1567.925 4.5125 ;
      RECT  1568.34 4.0975 1570.785 4.5125 ;
      RECT  1571.2 4.0975 1573.645 4.5125 ;
      RECT  1574.06 4.0975 1576.505 4.5125 ;
      RECT  1576.92 4.0975 1579.365 4.5125 ;
      RECT  1579.78 4.0975 1582.225 4.5125 ;
      RECT  1582.64 4.0975 1585.085 4.5125 ;
      RECT  1585.5 4.0975 1587.945 4.5125 ;
      RECT  1588.36 4.0975 1593.76 4.5125 ;
      RECT  0.14 148.5825 120.765 148.9975 ;
      RECT  120.765 4.5125 121.18 148.5825 ;
      RECT  121.18 4.5125 126.485 148.5825 ;
      RECT  121.18 148.5825 126.485 148.9975 ;
      RECT  120.765 148.9975 121.18 151.3125 ;
      RECT  120.765 151.7275 121.18 153.5225 ;
      RECT  120.765 153.9375 121.18 156.2525 ;
      RECT  120.765 156.6675 121.18 158.4625 ;
      RECT  120.765 158.8775 121.18 161.1925 ;
      RECT  0.14 4.5125 3.25 103.8625 ;
      RECT  0.14 103.8625 3.25 104.2775 ;
      RECT  0.14 104.2775 3.25 148.5825 ;
      RECT  3.25 4.5125 3.665 103.8625 ;
      RECT  3.665 4.5125 120.765 103.8625 ;
      RECT  3.25 104.2775 3.665 106.5925 ;
      RECT  3.25 107.0075 3.665 148.5825 ;
      RECT  3.665 103.8625 9.4925 103.9475 ;
      RECT  3.665 103.9475 9.4925 104.2775 ;
      RECT  9.4925 103.8625 9.9075 103.9475 ;
      RECT  9.9075 103.8625 120.765 103.9475 ;
      RECT  9.9075 103.9475 120.765 104.2775 ;
      RECT  3.665 104.2775 9.4925 104.3625 ;
      RECT  3.665 104.3625 9.4925 148.5825 ;
      RECT  9.4925 104.3625 9.9075 148.5825 ;
      RECT  9.9075 104.2775 120.765 104.3625 ;
      RECT  9.9075 104.3625 120.765 148.5825 ;
      RECT  126.9 4.5125 163.2525 115.51 ;
      RECT  126.9 115.51 163.2525 115.925 ;
      RECT  163.2525 4.5125 163.6675 115.51 ;
      RECT  163.6675 4.5125 1593.76 115.51 ;
      RECT  163.6675 115.51 163.9575 115.925 ;
      RECT  164.3725 115.51 164.6625 115.925 ;
      RECT  165.0775 115.51 165.3675 115.925 ;
      RECT  165.7825 115.51 166.0725 115.925 ;
      RECT  166.4875 115.51 166.7775 115.925 ;
      RECT  167.1925 115.51 167.4825 115.925 ;
      RECT  167.8975 115.51 168.1875 115.925 ;
      RECT  168.6025 115.51 168.8925 115.925 ;
      RECT  169.3075 115.51 169.5975 115.925 ;
      RECT  170.0125 115.51 170.3025 115.925 ;
      RECT  170.7175 115.51 171.0075 115.925 ;
      RECT  171.4225 115.51 171.7125 115.925 ;
      RECT  172.1275 115.51 172.4175 115.925 ;
      RECT  172.8325 115.51 173.1225 115.925 ;
      RECT  173.5375 115.51 173.8275 115.925 ;
      RECT  174.2425 115.51 174.5325 115.925 ;
      RECT  174.9475 115.51 175.2375 115.925 ;
      RECT  175.6525 115.51 175.9425 115.925 ;
      RECT  176.3575 115.51 176.6475 115.925 ;
      RECT  177.0625 115.51 177.3525 115.925 ;
      RECT  177.7675 115.51 178.0575 115.925 ;
      RECT  178.4725 115.51 178.7625 115.925 ;
      RECT  179.1775 115.51 179.4675 115.925 ;
      RECT  179.8825 115.51 180.1725 115.925 ;
      RECT  180.5875 115.51 180.8775 115.925 ;
      RECT  181.2925 115.51 181.5825 115.925 ;
      RECT  181.9975 115.51 182.2875 115.925 ;
      RECT  182.7025 115.51 182.9925 115.925 ;
      RECT  183.4075 115.51 183.6975 115.925 ;
      RECT  184.1125 115.51 184.4025 115.925 ;
      RECT  184.8175 115.51 185.1075 115.925 ;
      RECT  185.5225 115.51 185.8125 115.925 ;
      RECT  186.2275 115.51 186.5175 115.925 ;
      RECT  186.9325 115.51 187.2225 115.925 ;
      RECT  187.6375 115.51 187.9275 115.925 ;
      RECT  188.3425 115.51 188.6325 115.925 ;
      RECT  189.0475 115.51 189.3375 115.925 ;
      RECT  189.7525 115.51 190.0425 115.925 ;
      RECT  190.4575 115.51 190.7475 115.925 ;
      RECT  191.1625 115.51 191.4525 115.925 ;
      RECT  191.8675 115.51 192.1575 115.925 ;
      RECT  192.5725 115.51 192.8625 115.925 ;
      RECT  193.2775 115.51 193.5675 115.925 ;
      RECT  193.9825 115.51 194.2725 115.925 ;
      RECT  194.6875 115.51 194.9775 115.925 ;
      RECT  195.3925 115.51 195.6825 115.925 ;
      RECT  196.0975 115.51 196.3875 115.925 ;
      RECT  196.8025 115.51 197.0925 115.925 ;
      RECT  197.5075 115.51 197.7975 115.925 ;
      RECT  198.2125 115.51 198.5025 115.925 ;
      RECT  198.9175 115.51 199.2075 115.925 ;
      RECT  199.6225 115.51 199.9125 115.925 ;
      RECT  200.3275 115.51 200.6175 115.925 ;
      RECT  201.0325 115.51 201.3225 115.925 ;
      RECT  201.7375 115.51 202.0275 115.925 ;
      RECT  202.4425 115.51 202.7325 115.925 ;
      RECT  203.1475 115.51 203.4375 115.925 ;
      RECT  203.8525 115.51 204.1425 115.925 ;
      RECT  204.5575 115.51 204.8475 115.925 ;
      RECT  205.2625 115.51 205.5525 115.925 ;
      RECT  205.9675 115.51 206.2575 115.925 ;
      RECT  206.6725 115.51 206.9625 115.925 ;
      RECT  207.3775 115.51 207.6675 115.925 ;
      RECT  208.0825 115.51 208.3725 115.925 ;
      RECT  208.7875 115.51 209.0775 115.925 ;
      RECT  209.4925 115.51 209.7825 115.925 ;
      RECT  210.1975 115.51 210.4875 115.925 ;
      RECT  210.9025 115.51 211.1925 115.925 ;
      RECT  211.6075 115.51 211.8975 115.925 ;
      RECT  212.3125 115.51 212.6025 115.925 ;
      RECT  213.0175 115.51 213.3075 115.925 ;
      RECT  213.7225 115.51 214.0125 115.925 ;
      RECT  214.4275 115.51 214.7175 115.925 ;
      RECT  215.1325 115.51 215.4225 115.925 ;
      RECT  215.8375 115.51 216.1275 115.925 ;
      RECT  216.5425 115.51 216.8325 115.925 ;
      RECT  217.2475 115.51 217.5375 115.925 ;
      RECT  217.9525 115.51 218.2425 115.925 ;
      RECT  218.6575 115.51 218.9475 115.925 ;
      RECT  219.3625 115.51 219.6525 115.925 ;
      RECT  220.0675 115.51 220.3575 115.925 ;
      RECT  220.7725 115.51 221.0625 115.925 ;
      RECT  221.4775 115.51 221.7675 115.925 ;
      RECT  222.1825 115.51 222.4725 115.925 ;
      RECT  222.8875 115.51 223.1775 115.925 ;
      RECT  223.5925 115.51 223.8825 115.925 ;
      RECT  224.2975 115.51 224.5875 115.925 ;
      RECT  225.0025 115.51 225.2925 115.925 ;
      RECT  225.7075 115.51 225.9975 115.925 ;
      RECT  226.4125 115.51 226.7025 115.925 ;
      RECT  227.1175 115.51 227.4075 115.925 ;
      RECT  227.8225 115.51 228.1125 115.925 ;
      RECT  228.5275 115.51 228.8175 115.925 ;
      RECT  229.2325 115.51 229.5225 115.925 ;
      RECT  229.9375 115.51 230.2275 115.925 ;
      RECT  230.6425 115.51 230.9325 115.925 ;
      RECT  231.3475 115.51 231.6375 115.925 ;
      RECT  232.0525 115.51 232.3425 115.925 ;
      RECT  232.7575 115.51 233.0475 115.925 ;
      RECT  233.4625 115.51 233.7525 115.925 ;
      RECT  234.1675 115.51 234.4575 115.925 ;
      RECT  234.8725 115.51 235.1625 115.925 ;
      RECT  235.5775 115.51 235.8675 115.925 ;
      RECT  236.2825 115.51 236.5725 115.925 ;
      RECT  236.9875 115.51 237.2775 115.925 ;
      RECT  237.6925 115.51 237.9825 115.925 ;
      RECT  238.3975 115.51 238.6875 115.925 ;
      RECT  239.1025 115.51 239.3925 115.925 ;
      RECT  239.8075 115.51 240.0975 115.925 ;
      RECT  240.5125 115.51 240.8025 115.925 ;
      RECT  241.2175 115.51 241.5075 115.925 ;
      RECT  241.9225 115.51 242.2125 115.925 ;
      RECT  242.6275 115.51 242.9175 115.925 ;
      RECT  243.3325 115.51 243.6225 115.925 ;
      RECT  244.0375 115.51 244.3275 115.925 ;
      RECT  244.7425 115.51 245.0325 115.925 ;
      RECT  245.4475 115.51 245.7375 115.925 ;
      RECT  246.1525 115.51 246.4425 115.925 ;
      RECT  246.8575 115.51 247.1475 115.925 ;
      RECT  247.5625 115.51 247.8525 115.925 ;
      RECT  248.2675 115.51 248.5575 115.925 ;
      RECT  248.9725 115.51 249.2625 115.925 ;
      RECT  249.6775 115.51 249.9675 115.925 ;
      RECT  250.3825 115.51 250.6725 115.925 ;
      RECT  251.0875 115.51 251.3775 115.925 ;
      RECT  251.7925 115.51 252.0825 115.925 ;
      RECT  252.4975 115.51 252.7875 115.925 ;
      RECT  253.2025 115.51 253.4925 115.925 ;
      RECT  253.9075 115.51 254.1975 115.925 ;
      RECT  254.6125 115.51 254.9025 115.925 ;
      RECT  255.3175 115.51 255.6075 115.925 ;
      RECT  256.0225 115.51 256.3125 115.925 ;
      RECT  256.7275 115.51 257.0175 115.925 ;
      RECT  257.4325 115.51 257.7225 115.925 ;
      RECT  258.1375 115.51 258.4275 115.925 ;
      RECT  258.8425 115.51 259.1325 115.925 ;
      RECT  259.5475 115.51 259.8375 115.925 ;
      RECT  260.2525 115.51 260.5425 115.925 ;
      RECT  260.9575 115.51 261.2475 115.925 ;
      RECT  261.6625 115.51 261.9525 115.925 ;
      RECT  262.3675 115.51 262.6575 115.925 ;
      RECT  263.0725 115.51 263.3625 115.925 ;
      RECT  263.7775 115.51 264.0675 115.925 ;
      RECT  264.4825 115.51 264.7725 115.925 ;
      RECT  265.1875 115.51 265.4775 115.925 ;
      RECT  265.8925 115.51 266.1825 115.925 ;
      RECT  266.5975 115.51 266.8875 115.925 ;
      RECT  267.3025 115.51 267.5925 115.925 ;
      RECT  268.0075 115.51 268.2975 115.925 ;
      RECT  268.7125 115.51 269.0025 115.925 ;
      RECT  269.4175 115.51 269.7075 115.925 ;
      RECT  270.1225 115.51 270.4125 115.925 ;
      RECT  270.8275 115.51 271.1175 115.925 ;
      RECT  271.5325 115.51 271.8225 115.925 ;
      RECT  272.2375 115.51 272.5275 115.925 ;
      RECT  272.9425 115.51 273.2325 115.925 ;
      RECT  273.6475 115.51 273.9375 115.925 ;
      RECT  274.3525 115.51 274.6425 115.925 ;
      RECT  275.0575 115.51 275.3475 115.925 ;
      RECT  275.7625 115.51 276.0525 115.925 ;
      RECT  276.4675 115.51 276.7575 115.925 ;
      RECT  277.1725 115.51 277.4625 115.925 ;
      RECT  277.8775 115.51 278.1675 115.925 ;
      RECT  278.5825 115.51 278.8725 115.925 ;
      RECT  279.2875 115.51 279.5775 115.925 ;
      RECT  279.9925 115.51 280.2825 115.925 ;
      RECT  280.6975 115.51 280.9875 115.925 ;
      RECT  281.4025 115.51 281.6925 115.925 ;
      RECT  282.1075 115.51 282.3975 115.925 ;
      RECT  282.8125 115.51 283.1025 115.925 ;
      RECT  283.5175 115.51 283.8075 115.925 ;
      RECT  284.2225 115.51 284.5125 115.925 ;
      RECT  284.9275 115.51 285.2175 115.925 ;
      RECT  285.6325 115.51 285.9225 115.925 ;
      RECT  286.3375 115.51 286.6275 115.925 ;
      RECT  287.0425 115.51 287.3325 115.925 ;
      RECT  287.7475 115.51 288.0375 115.925 ;
      RECT  288.4525 115.51 288.7425 115.925 ;
      RECT  289.1575 115.51 289.4475 115.925 ;
      RECT  289.8625 115.51 290.1525 115.925 ;
      RECT  290.5675 115.51 290.8575 115.925 ;
      RECT  291.2725 115.51 291.5625 115.925 ;
      RECT  291.9775 115.51 292.2675 115.925 ;
      RECT  292.6825 115.51 292.9725 115.925 ;
      RECT  293.3875 115.51 293.6775 115.925 ;
      RECT  294.0925 115.51 294.3825 115.925 ;
      RECT  294.7975 115.51 295.0875 115.925 ;
      RECT  295.5025 115.51 295.7925 115.925 ;
      RECT  296.2075 115.51 296.4975 115.925 ;
      RECT  296.9125 115.51 297.2025 115.925 ;
      RECT  297.6175 115.51 297.9075 115.925 ;
      RECT  298.3225 115.51 298.6125 115.925 ;
      RECT  299.0275 115.51 299.3175 115.925 ;
      RECT  299.7325 115.51 300.0225 115.925 ;
      RECT  300.4375 115.51 300.7275 115.925 ;
      RECT  301.1425 115.51 301.4325 115.925 ;
      RECT  301.8475 115.51 302.1375 115.925 ;
      RECT  302.5525 115.51 302.8425 115.925 ;
      RECT  303.2575 115.51 303.5475 115.925 ;
      RECT  303.9625 115.51 304.2525 115.925 ;
      RECT  304.6675 115.51 304.9575 115.925 ;
      RECT  305.3725 115.51 305.6625 115.925 ;
      RECT  306.0775 115.51 306.3675 115.925 ;
      RECT  306.7825 115.51 307.0725 115.925 ;
      RECT  307.4875 115.51 307.7775 115.925 ;
      RECT  308.1925 115.51 308.4825 115.925 ;
      RECT  308.8975 115.51 309.1875 115.925 ;
      RECT  309.6025 115.51 309.8925 115.925 ;
      RECT  310.3075 115.51 310.5975 115.925 ;
      RECT  311.0125 115.51 311.3025 115.925 ;
      RECT  311.7175 115.51 312.0075 115.925 ;
      RECT  312.4225 115.51 312.7125 115.925 ;
      RECT  313.1275 115.51 313.4175 115.925 ;
      RECT  313.8325 115.51 314.1225 115.925 ;
      RECT  314.5375 115.51 314.8275 115.925 ;
      RECT  315.2425 115.51 315.5325 115.925 ;
      RECT  315.9475 115.51 316.2375 115.925 ;
      RECT  316.6525 115.51 316.9425 115.925 ;
      RECT  317.3575 115.51 317.6475 115.925 ;
      RECT  318.0625 115.51 318.3525 115.925 ;
      RECT  318.7675 115.51 319.0575 115.925 ;
      RECT  319.4725 115.51 319.7625 115.925 ;
      RECT  320.1775 115.51 320.4675 115.925 ;
      RECT  320.8825 115.51 321.1725 115.925 ;
      RECT  321.5875 115.51 321.8775 115.925 ;
      RECT  322.2925 115.51 322.5825 115.925 ;
      RECT  322.9975 115.51 323.2875 115.925 ;
      RECT  323.7025 115.51 323.9925 115.925 ;
      RECT  324.4075 115.51 324.6975 115.925 ;
      RECT  325.1125 115.51 325.4025 115.925 ;
      RECT  325.8175 115.51 326.1075 115.925 ;
      RECT  326.5225 115.51 326.8125 115.925 ;
      RECT  327.2275 115.51 327.5175 115.925 ;
      RECT  327.9325 115.51 328.2225 115.925 ;
      RECT  328.6375 115.51 328.9275 115.925 ;
      RECT  329.3425 115.51 329.6325 115.925 ;
      RECT  330.0475 115.51 330.3375 115.925 ;
      RECT  330.7525 115.51 331.0425 115.925 ;
      RECT  331.4575 115.51 331.7475 115.925 ;
      RECT  332.1625 115.51 332.4525 115.925 ;
      RECT  332.8675 115.51 333.1575 115.925 ;
      RECT  333.5725 115.51 333.8625 115.925 ;
      RECT  334.2775 115.51 334.5675 115.925 ;
      RECT  334.9825 115.51 335.2725 115.925 ;
      RECT  335.6875 115.51 335.9775 115.925 ;
      RECT  336.3925 115.51 336.6825 115.925 ;
      RECT  337.0975 115.51 337.3875 115.925 ;
      RECT  337.8025 115.51 338.0925 115.925 ;
      RECT  338.5075 115.51 338.7975 115.925 ;
      RECT  339.2125 115.51 339.5025 115.925 ;
      RECT  339.9175 115.51 340.2075 115.925 ;
      RECT  340.6225 115.51 340.9125 115.925 ;
      RECT  341.3275 115.51 341.6175 115.925 ;
      RECT  342.0325 115.51 342.3225 115.925 ;
      RECT  342.7375 115.51 343.0275 115.925 ;
      RECT  343.4425 115.51 343.7325 115.925 ;
      RECT  344.1475 115.51 344.4375 115.925 ;
      RECT  344.8525 115.51 345.1425 115.925 ;
      RECT  345.5575 115.51 345.8475 115.925 ;
      RECT  346.2625 115.51 346.5525 115.925 ;
      RECT  346.9675 115.51 347.2575 115.925 ;
      RECT  347.6725 115.51 347.9625 115.925 ;
      RECT  348.3775 115.51 348.6675 115.925 ;
      RECT  349.0825 115.51 349.3725 115.925 ;
      RECT  349.7875 115.51 350.0775 115.925 ;
      RECT  350.4925 115.51 350.7825 115.925 ;
      RECT  351.1975 115.51 351.4875 115.925 ;
      RECT  351.9025 115.51 352.1925 115.925 ;
      RECT  352.6075 115.51 352.8975 115.925 ;
      RECT  353.3125 115.51 353.6025 115.925 ;
      RECT  354.0175 115.51 354.3075 115.925 ;
      RECT  354.7225 115.51 355.0125 115.925 ;
      RECT  355.4275 115.51 355.7175 115.925 ;
      RECT  356.1325 115.51 356.4225 115.925 ;
      RECT  356.8375 115.51 357.1275 115.925 ;
      RECT  357.5425 115.51 357.8325 115.925 ;
      RECT  358.2475 115.51 358.5375 115.925 ;
      RECT  358.9525 115.51 359.2425 115.925 ;
      RECT  359.6575 115.51 359.9475 115.925 ;
      RECT  360.3625 115.51 360.6525 115.925 ;
      RECT  361.0675 115.51 361.3575 115.925 ;
      RECT  361.7725 115.51 362.0625 115.925 ;
      RECT  362.4775 115.51 362.7675 115.925 ;
      RECT  363.1825 115.51 363.4725 115.925 ;
      RECT  363.8875 115.51 364.1775 115.925 ;
      RECT  364.5925 115.51 364.8825 115.925 ;
      RECT  365.2975 115.51 365.5875 115.925 ;
      RECT  366.0025 115.51 366.2925 115.925 ;
      RECT  366.7075 115.51 366.9975 115.925 ;
      RECT  367.4125 115.51 367.7025 115.925 ;
      RECT  368.1175 115.51 368.4075 115.925 ;
      RECT  368.8225 115.51 369.1125 115.925 ;
      RECT  369.5275 115.51 369.8175 115.925 ;
      RECT  370.2325 115.51 370.5225 115.925 ;
      RECT  370.9375 115.51 371.2275 115.925 ;
      RECT  371.6425 115.51 371.9325 115.925 ;
      RECT  372.3475 115.51 372.6375 115.925 ;
      RECT  373.0525 115.51 373.3425 115.925 ;
      RECT  373.7575 115.51 374.0475 115.925 ;
      RECT  374.4625 115.51 374.7525 115.925 ;
      RECT  375.1675 115.51 375.4575 115.925 ;
      RECT  375.8725 115.51 376.1625 115.925 ;
      RECT  376.5775 115.51 376.8675 115.925 ;
      RECT  377.2825 115.51 377.5725 115.925 ;
      RECT  377.9875 115.51 378.2775 115.925 ;
      RECT  378.6925 115.51 378.9825 115.925 ;
      RECT  379.3975 115.51 379.6875 115.925 ;
      RECT  380.1025 115.51 380.3925 115.925 ;
      RECT  380.8075 115.51 381.0975 115.925 ;
      RECT  381.5125 115.51 381.8025 115.925 ;
      RECT  382.2175 115.51 382.5075 115.925 ;
      RECT  382.9225 115.51 383.2125 115.925 ;
      RECT  383.6275 115.51 383.9175 115.925 ;
      RECT  384.3325 115.51 384.6225 115.925 ;
      RECT  385.0375 115.51 385.3275 115.925 ;
      RECT  385.7425 115.51 386.0325 115.925 ;
      RECT  386.4475 115.51 386.7375 115.925 ;
      RECT  387.1525 115.51 387.4425 115.925 ;
      RECT  387.8575 115.51 388.1475 115.925 ;
      RECT  388.5625 115.51 388.8525 115.925 ;
      RECT  389.2675 115.51 389.5575 115.925 ;
      RECT  389.9725 115.51 390.2625 115.925 ;
      RECT  390.6775 115.51 390.9675 115.925 ;
      RECT  391.3825 115.51 391.6725 115.925 ;
      RECT  392.0875 115.51 392.3775 115.925 ;
      RECT  392.7925 115.51 393.0825 115.925 ;
      RECT  393.4975 115.51 393.7875 115.925 ;
      RECT  394.2025 115.51 394.4925 115.925 ;
      RECT  394.9075 115.51 395.1975 115.925 ;
      RECT  395.6125 115.51 395.9025 115.925 ;
      RECT  396.3175 115.51 396.6075 115.925 ;
      RECT  397.0225 115.51 397.3125 115.925 ;
      RECT  397.7275 115.51 398.0175 115.925 ;
      RECT  398.4325 115.51 398.7225 115.925 ;
      RECT  399.1375 115.51 399.4275 115.925 ;
      RECT  399.8425 115.51 400.1325 115.925 ;
      RECT  400.5475 115.51 400.8375 115.925 ;
      RECT  401.2525 115.51 401.5425 115.925 ;
      RECT  401.9575 115.51 402.2475 115.925 ;
      RECT  402.6625 115.51 402.9525 115.925 ;
      RECT  403.3675 115.51 403.6575 115.925 ;
      RECT  404.0725 115.51 404.3625 115.925 ;
      RECT  404.7775 115.51 405.0675 115.925 ;
      RECT  405.4825 115.51 405.7725 115.925 ;
      RECT  406.1875 115.51 406.4775 115.925 ;
      RECT  406.8925 115.51 407.1825 115.925 ;
      RECT  407.5975 115.51 407.8875 115.925 ;
      RECT  408.3025 115.51 408.5925 115.925 ;
      RECT  409.0075 115.51 409.2975 115.925 ;
      RECT  409.7125 115.51 410.0025 115.925 ;
      RECT  410.4175 115.51 410.7075 115.925 ;
      RECT  411.1225 115.51 411.4125 115.925 ;
      RECT  411.8275 115.51 412.1175 115.925 ;
      RECT  412.5325 115.51 412.8225 115.925 ;
      RECT  413.2375 115.51 413.5275 115.925 ;
      RECT  413.9425 115.51 414.2325 115.925 ;
      RECT  414.6475 115.51 414.9375 115.925 ;
      RECT  415.3525 115.51 415.6425 115.925 ;
      RECT  416.0575 115.51 416.3475 115.925 ;
      RECT  416.7625 115.51 417.0525 115.925 ;
      RECT  417.4675 115.51 417.7575 115.925 ;
      RECT  418.1725 115.51 418.4625 115.925 ;
      RECT  418.8775 115.51 419.1675 115.925 ;
      RECT  419.5825 115.51 419.8725 115.925 ;
      RECT  420.2875 115.51 420.5775 115.925 ;
      RECT  420.9925 115.51 421.2825 115.925 ;
      RECT  421.6975 115.51 421.9875 115.925 ;
      RECT  422.4025 115.51 422.6925 115.925 ;
      RECT  423.1075 115.51 423.3975 115.925 ;
      RECT  423.8125 115.51 424.1025 115.925 ;
      RECT  424.5175 115.51 424.8075 115.925 ;
      RECT  425.2225 115.51 425.5125 115.925 ;
      RECT  425.9275 115.51 426.2175 115.925 ;
      RECT  426.6325 115.51 426.9225 115.925 ;
      RECT  427.3375 115.51 427.6275 115.925 ;
      RECT  428.0425 115.51 428.3325 115.925 ;
      RECT  428.7475 115.51 429.0375 115.925 ;
      RECT  429.4525 115.51 429.7425 115.925 ;
      RECT  430.1575 115.51 430.4475 115.925 ;
      RECT  430.8625 115.51 431.1525 115.925 ;
      RECT  431.5675 115.51 431.8575 115.925 ;
      RECT  432.2725 115.51 432.5625 115.925 ;
      RECT  432.9775 115.51 433.2675 115.925 ;
      RECT  433.6825 115.51 433.9725 115.925 ;
      RECT  434.3875 115.51 434.6775 115.925 ;
      RECT  435.0925 115.51 435.3825 115.925 ;
      RECT  435.7975 115.51 436.0875 115.925 ;
      RECT  436.5025 115.51 436.7925 115.925 ;
      RECT  437.2075 115.51 437.4975 115.925 ;
      RECT  437.9125 115.51 438.2025 115.925 ;
      RECT  438.6175 115.51 438.9075 115.925 ;
      RECT  439.3225 115.51 439.6125 115.925 ;
      RECT  440.0275 115.51 440.3175 115.925 ;
      RECT  440.7325 115.51 441.0225 115.925 ;
      RECT  441.4375 115.51 441.7275 115.925 ;
      RECT  442.1425 115.51 442.4325 115.925 ;
      RECT  442.8475 115.51 443.1375 115.925 ;
      RECT  443.5525 115.51 443.8425 115.925 ;
      RECT  444.2575 115.51 444.5475 115.925 ;
      RECT  444.9625 115.51 445.2525 115.925 ;
      RECT  445.6675 115.51 445.9575 115.925 ;
      RECT  446.3725 115.51 446.6625 115.925 ;
      RECT  447.0775 115.51 447.3675 115.925 ;
      RECT  447.7825 115.51 448.0725 115.925 ;
      RECT  448.4875 115.51 448.7775 115.925 ;
      RECT  449.1925 115.51 449.4825 115.925 ;
      RECT  449.8975 115.51 450.1875 115.925 ;
      RECT  450.6025 115.51 450.8925 115.925 ;
      RECT  451.3075 115.51 451.5975 115.925 ;
      RECT  452.0125 115.51 452.3025 115.925 ;
      RECT  452.7175 115.51 453.0075 115.925 ;
      RECT  453.4225 115.51 453.7125 115.925 ;
      RECT  454.1275 115.51 454.4175 115.925 ;
      RECT  454.8325 115.51 455.1225 115.925 ;
      RECT  455.5375 115.51 455.8275 115.925 ;
      RECT  456.2425 115.51 456.5325 115.925 ;
      RECT  456.9475 115.51 457.2375 115.925 ;
      RECT  457.6525 115.51 457.9425 115.925 ;
      RECT  458.3575 115.51 458.6475 115.925 ;
      RECT  459.0625 115.51 459.3525 115.925 ;
      RECT  459.7675 115.51 460.0575 115.925 ;
      RECT  460.4725 115.51 460.7625 115.925 ;
      RECT  461.1775 115.51 461.4675 115.925 ;
      RECT  461.8825 115.51 462.1725 115.925 ;
      RECT  462.5875 115.51 462.8775 115.925 ;
      RECT  463.2925 115.51 463.5825 115.925 ;
      RECT  463.9975 115.51 464.2875 115.925 ;
      RECT  464.7025 115.51 464.9925 115.925 ;
      RECT  465.4075 115.51 465.6975 115.925 ;
      RECT  466.1125 115.51 466.4025 115.925 ;
      RECT  466.8175 115.51 467.1075 115.925 ;
      RECT  467.5225 115.51 467.8125 115.925 ;
      RECT  468.2275 115.51 468.5175 115.925 ;
      RECT  468.9325 115.51 469.2225 115.925 ;
      RECT  469.6375 115.51 469.9275 115.925 ;
      RECT  470.3425 115.51 470.6325 115.925 ;
      RECT  471.0475 115.51 471.3375 115.925 ;
      RECT  471.7525 115.51 472.0425 115.925 ;
      RECT  472.4575 115.51 472.7475 115.925 ;
      RECT  473.1625 115.51 473.4525 115.925 ;
      RECT  473.8675 115.51 474.1575 115.925 ;
      RECT  474.5725 115.51 474.8625 115.925 ;
      RECT  475.2775 115.51 475.5675 115.925 ;
      RECT  475.9825 115.51 476.2725 115.925 ;
      RECT  476.6875 115.51 476.9775 115.925 ;
      RECT  477.3925 115.51 477.6825 115.925 ;
      RECT  478.0975 115.51 478.3875 115.925 ;
      RECT  478.8025 115.51 479.0925 115.925 ;
      RECT  479.5075 115.51 479.7975 115.925 ;
      RECT  480.2125 115.51 480.5025 115.925 ;
      RECT  480.9175 115.51 481.2075 115.925 ;
      RECT  481.6225 115.51 481.9125 115.925 ;
      RECT  482.3275 115.51 482.6175 115.925 ;
      RECT  483.0325 115.51 483.3225 115.925 ;
      RECT  483.7375 115.51 484.0275 115.925 ;
      RECT  484.4425 115.51 484.7325 115.925 ;
      RECT  485.1475 115.51 485.4375 115.925 ;
      RECT  485.8525 115.51 486.1425 115.925 ;
      RECT  486.5575 115.51 486.8475 115.925 ;
      RECT  487.2625 115.51 487.5525 115.925 ;
      RECT  487.9675 115.51 488.2575 115.925 ;
      RECT  488.6725 115.51 488.9625 115.925 ;
      RECT  489.3775 115.51 489.6675 115.925 ;
      RECT  490.0825 115.51 490.3725 115.925 ;
      RECT  490.7875 115.51 491.0775 115.925 ;
      RECT  491.4925 115.51 491.7825 115.925 ;
      RECT  492.1975 115.51 492.4875 115.925 ;
      RECT  492.9025 115.51 493.1925 115.925 ;
      RECT  493.6075 115.51 493.8975 115.925 ;
      RECT  494.3125 115.51 494.6025 115.925 ;
      RECT  495.0175 115.51 495.3075 115.925 ;
      RECT  495.7225 115.51 496.0125 115.925 ;
      RECT  496.4275 115.51 496.7175 115.925 ;
      RECT  497.1325 115.51 497.4225 115.925 ;
      RECT  497.8375 115.51 498.1275 115.925 ;
      RECT  498.5425 115.51 498.8325 115.925 ;
      RECT  499.2475 115.51 499.5375 115.925 ;
      RECT  499.9525 115.51 500.2425 115.925 ;
      RECT  500.6575 115.51 500.9475 115.925 ;
      RECT  501.3625 115.51 501.6525 115.925 ;
      RECT  502.0675 115.51 502.3575 115.925 ;
      RECT  502.7725 115.51 503.0625 115.925 ;
      RECT  503.4775 115.51 503.7675 115.925 ;
      RECT  504.1825 115.51 504.4725 115.925 ;
      RECT  504.8875 115.51 505.1775 115.925 ;
      RECT  505.5925 115.51 505.8825 115.925 ;
      RECT  506.2975 115.51 506.5875 115.925 ;
      RECT  507.0025 115.51 507.2925 115.925 ;
      RECT  507.7075 115.51 507.9975 115.925 ;
      RECT  508.4125 115.51 508.7025 115.925 ;
      RECT  509.1175 115.51 509.4075 115.925 ;
      RECT  509.8225 115.51 510.1125 115.925 ;
      RECT  510.5275 115.51 510.8175 115.925 ;
      RECT  511.2325 115.51 511.5225 115.925 ;
      RECT  511.9375 115.51 512.2275 115.925 ;
      RECT  512.6425 115.51 512.9325 115.925 ;
      RECT  513.3475 115.51 513.6375 115.925 ;
      RECT  514.0525 115.51 514.3425 115.925 ;
      RECT  514.7575 115.51 515.0475 115.925 ;
      RECT  515.4625 115.51 515.7525 115.925 ;
      RECT  516.1675 115.51 516.4575 115.925 ;
      RECT  516.8725 115.51 517.1625 115.925 ;
      RECT  517.5775 115.51 517.8675 115.925 ;
      RECT  518.2825 115.51 518.5725 115.925 ;
      RECT  518.9875 115.51 519.2775 115.925 ;
      RECT  519.6925 115.51 519.9825 115.925 ;
      RECT  520.3975 115.51 520.6875 115.925 ;
      RECT  521.1025 115.51 521.3925 115.925 ;
      RECT  521.8075 115.51 522.0975 115.925 ;
      RECT  522.5125 115.51 522.8025 115.925 ;
      RECT  523.2175 115.51 523.5075 115.925 ;
      RECT  523.9225 115.51 1593.76 115.925 ;
      RECT  126.485 4.5125 126.9 216.58 ;
      RECT  0.14 148.9975 1.26 216.58 ;
      RECT  0.14 216.58 1.26 217.56 ;
      RECT  1.26 148.9975 120.765 216.58 ;
      RECT  121.18 148.9975 126.485 216.58 ;
      RECT  120.765 161.6075 121.18 216.58 ;
      RECT  126.9 115.925 163.2525 216.58 ;
      RECT  163.2525 115.925 163.6675 216.58 ;
      RECT  163.6675 115.925 1592.64 216.58 ;
      RECT  1592.64 115.925 1593.76 216.58 ;
      RECT  1592.64 216.58 1593.76 217.56 ;
      RECT  0.14 1.26 1.26 2.24 ;
      RECT  0.14 2.24 1.26 4.0975 ;
      RECT  1.26 2.24 126.485 4.0975 ;
      RECT  126.485 2.24 126.9 4.0975 ;
      RECT  126.9 2.24 1592.64 4.0975 ;
      RECT  1592.64 1.26 1593.76 2.24 ;
      RECT  1592.64 2.24 1593.76 4.0975 ;
      RECT  126.485 217.56 126.9 217.98 ;
      RECT  0.14 217.56 1.26 217.98 ;
      RECT  1.26 217.56 120.765 217.98 ;
      RECT  121.18 217.56 126.485 217.98 ;
      RECT  120.765 217.56 121.18 217.98 ;
      RECT  126.9 217.56 163.2525 217.98 ;
      RECT  163.2525 217.56 163.6675 217.98 ;
      RECT  163.6675 217.56 1592.64 217.98 ;
      RECT  1592.64 217.56 1593.76 217.98 ;
      RECT  0.14 0.84 1.26 1.26 ;
      RECT  1.26 0.84 126.485 1.26 ;
      RECT  126.485 0.84 126.9 1.26 ;
      RECT  126.9 0.84 1592.64 1.26 ;
      RECT  1592.64 0.84 1593.76 1.26 ;
   LAYER  metal4 ;
      RECT  1.12 0.14 2.38 1.12 ;
      RECT  1.12 217.7 2.38 218.68 ;
      RECT  2.38 1.12 1591.52 217.7 ;
      RECT  2.38 0.14 1592.92 1.12 ;
      RECT  2.38 217.7 1592.92 218.68 ;
      RECT  1592.78 1.12 1592.92 217.7 ;
      RECT  0.98 0.14 1.12 1.12 ;
      RECT  0.98 1.12 1.12 217.7 ;
      RECT  0.98 217.7 1.12 218.68 ;
   END
END    freepdk45_sram_1rw0r_64x512
END    LIBRARY
