VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_128x40
   CLASS BLOCK ;
   SIZE 170.995 BY 134.51 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  25.725 1.1075 25.86 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.585 1.1075 28.72 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.445 1.1075 31.58 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.305 1.1075 34.44 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.165 1.1075 37.3 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.025 1.1075 40.16 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.885 1.1075 43.02 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.745 1.1075 45.88 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.605 1.1075 48.74 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.465 1.1075 51.6 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.325 1.1075 54.46 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.185 1.1075 57.32 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.045 1.1075 60.18 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.905 1.1075 63.04 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.765 1.1075 65.9 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.625 1.1075 68.76 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.485 1.1075 71.62 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.345 1.1075 74.48 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.205 1.1075 77.34 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.065 1.1075 80.2 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.925 1.1075 83.06 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.785 1.1075 85.92 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.645 1.1075 88.78 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.505 1.1075 91.64 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.365 1.1075 94.5 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.225 1.1075 97.36 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.085 1.1075 100.22 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.945 1.1075 103.08 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.805 1.1075 105.94 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.665 1.1075 108.8 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.525 1.1075 111.66 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.385 1.1075 114.52 1.2425 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.245 1.1075 117.38 1.2425 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.105 1.1075 120.24 1.2425 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.965 1.1075 123.1 1.2425 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.825 1.1075 125.96 1.2425 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.685 1.1075 128.82 1.2425 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.545 1.1075 131.68 1.2425 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.405 1.1075 134.54 1.2425 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.265 1.1075 137.4 1.2425 ;
      END
   END din0[39]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  22.865 1.1075 23.0 1.2425 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.145 45.6975 17.28 45.8325 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.145 48.4275 17.28 48.5625 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.145 50.6375 17.28 50.7725 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.145 53.3675 17.28 53.5025 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.145 55.5775 17.28 55.7125 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.145 58.3075 17.28 58.4425 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.995 132.0025 145.13 132.1375 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.575 19.5675 153.71 19.7025 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.575 16.8375 153.71 16.9725 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.575 14.6275 153.71 14.7625 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.575 11.8975 153.71 12.0325 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.575 9.6875 153.71 9.8225 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.575 6.9575 153.71 7.0925 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.575 133.2675 170.71 133.4025 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.4725 133.1825 164.6075 133.3175 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.2975 129.515 38.4325 129.65 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.6475 129.515 40.7825 129.65 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.9975 129.515 43.1325 129.65 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.3475 129.515 45.4825 129.65 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.6975 129.515 47.8325 129.65 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.0475 129.515 50.1825 129.65 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.3975 129.515 52.5325 129.65 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.7475 129.515 54.8825 129.65 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.0975 129.515 57.2325 129.65 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.4475 129.515 59.5825 129.65 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.7975 129.515 61.9325 129.65 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.1475 129.515 64.2825 129.65 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.4975 129.515 66.6325 129.65 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.8475 129.515 68.9825 129.65 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.1975 129.515 71.3325 129.65 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.5475 129.515 73.6825 129.65 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.8975 129.515 76.0325 129.65 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.2475 129.515 78.3825 129.65 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.5975 129.515 80.7325 129.65 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.9475 129.515 83.0825 129.65 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.2975 129.515 85.4325 129.65 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.6475 129.515 87.7825 129.65 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.9975 129.515 90.1325 129.65 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.3475 129.515 92.4825 129.65 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.6975 129.515 94.8325 129.65 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.0475 129.515 97.1825 129.65 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.3975 129.515 99.5325 129.65 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.7475 129.515 101.8825 129.65 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.0975 129.515 104.2325 129.65 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.4475 129.515 106.5825 129.65 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.7975 129.515 108.9325 129.65 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.1475 129.515 111.2825 129.65 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.4975 129.515 113.6325 129.65 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.8475 129.515 115.9825 129.65 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.1975 129.515 118.3325 129.65 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.5475 129.515 120.6825 129.65 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.8975 129.515 123.0325 129.65 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.2475 129.515 125.3825 129.65 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.5975 129.515 127.7325 129.65 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.9475 129.515 130.0825 129.65 ;
      END
   END dout1[39]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  142.005 20.67 142.145 116.56 ;
         LAYER metal4 ;
         RECT  170.1675 102.26 170.3075 124.6625 ;
         LAYER metal4 ;
         RECT  35.045 17.5 35.185 119.41 ;
         LAYER metal3 ;
         RECT  82.6425 2.4725 82.7775 2.6075 ;
         LAYER metal3 ;
         RECT  71.2025 2.4725 71.3375 2.6075 ;
         LAYER metal4 ;
         RECT  16.86 44.59 17.0 59.55 ;
         LAYER metal3 ;
         RECT  29.135 19.965 29.27 20.1 ;
         LAYER metal4 ;
         RECT  135.475 17.5 135.615 119.41 ;
         LAYER metal3 ;
         RECT  22.9625 31.1375 23.0975 31.2725 ;
         LAYER metal3 ;
         RECT  35.1125 8.415 130.7525 8.485 ;
         LAYER metal3 ;
         RECT  147.5625 25.1575 147.6975 25.2925 ;
         LAYER metal4 ;
         RECT  136.555 20.67 136.695 116.49 ;
         LAYER metal3 ;
         RECT  116.9625 2.4725 117.0975 2.6075 ;
         LAYER metal3 ;
         RECT  147.5625 43.0975 147.6975 43.2325 ;
         LAYER metal4 ;
         RECT  19.58 2.47 19.72 17.43 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal3 ;
         RECT  22.9625 22.1675 23.0975 22.3025 ;
         LAYER metal3 ;
         RECT  22.9625 43.0975 23.0975 43.2325 ;
         LAYER metal3 ;
         RECT  27.225 11.9075 27.36 12.0425 ;
         LAYER metal3 ;
         RECT  35.1125 126.9575 130.7525 127.0275 ;
         LAYER metal3 ;
         RECT  22.9625 34.1275 23.0975 34.2625 ;
         LAYER metal3 ;
         RECT  141.39 117.06 141.525 117.195 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
         LAYER metal4 ;
         RECT  151.135 122.02 151.275 132.04 ;
         LAYER metal4 ;
         RECT  28.515 20.67 28.655 116.56 ;
         LAYER metal3 ;
         RECT  35.1125 120.105 133.5725 120.175 ;
         LAYER metal3 ;
         RECT  22.5825 2.4725 22.7175 2.6075 ;
         LAYER metal3 ;
         RECT  168.435 131.9025 168.57 132.0375 ;
         LAYER metal3 ;
         RECT  145.2775 130.6375 145.4125 130.7725 ;
         LAYER metal3 ;
         RECT  25.4425 2.4725 25.5775 2.6075 ;
         LAYER metal4 ;
         RECT  153.855 5.85 153.995 20.81 ;
         LAYER metal3 ;
         RECT  147.5625 22.1675 147.6975 22.3025 ;
         LAYER metal3 ;
         RECT  33.9675 19.1775 34.1025 19.3125 ;
         LAYER metal4 ;
         RECT  33.965 20.67 34.105 116.49 ;
         LAYER metal3 ;
         RECT  94.0825 2.4725 94.2175 2.6075 ;
         LAYER metal3 ;
         RECT  22.9625 25.1575 23.0975 25.2925 ;
         LAYER metal3 ;
         RECT  147.5625 40.1075 147.6975 40.2425 ;
         LAYER metal3 ;
         RECT  48.3225 2.4725 48.4575 2.6075 ;
         LAYER metal3 ;
         RECT  22.9625 40.1075 23.0975 40.2425 ;
         LAYER metal3 ;
         RECT  147.5625 34.1275 147.6975 34.2625 ;
         LAYER metal3 ;
         RECT  59.7625 2.4725 59.8975 2.6075 ;
         LAYER metal3 ;
         RECT  128.4025 2.4725 128.5375 2.6075 ;
         LAYER metal3 ;
         RECT  36.8825 2.4725 37.0175 2.6075 ;
         LAYER metal3 ;
         RECT  147.5625 31.1375 147.6975 31.2725 ;
         LAYER metal3 ;
         RECT  143.3 124.9375 143.435 125.0725 ;
         LAYER metal3 ;
         RECT  105.5225 2.4725 105.6575 2.6075 ;
         LAYER metal3 ;
         RECT  35.1125 16.805 132.3975 16.875 ;
         LAYER metal3 ;
         RECT  136.5575 117.8475 136.6925 117.9825 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  21.435 35.6225 21.57 35.7575 ;
         LAYER metal3 ;
         RECT  149.09 32.6325 149.225 32.7675 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal4 ;
         RECT  150.995 5.785 151.135 20.875 ;
         LAYER metal4 ;
         RECT  141.445 20.6375 141.585 116.5225 ;
         LAYER metal4 ;
         RECT  19.72 44.525 19.86 59.615 ;
         LAYER metal4 ;
         RECT  29.075 20.6375 29.215 116.5225 ;
         LAYER metal3 ;
         RECT  143.3 127.4075 143.435 127.5425 ;
         LAYER metal3 ;
         RECT  149.09 26.6525 149.225 26.7875 ;
         LAYER metal3 ;
         RECT  51.1825 0.0025 51.3175 0.1375 ;
         LAYER metal3 ;
         RECT  21.435 20.6725 21.57 20.8075 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal4 ;
         RECT  26.58 20.6375 26.72 116.56 ;
         LAYER metal3 ;
         RECT  85.5025 0.0025 85.6375 0.1375 ;
         LAYER metal3 ;
         RECT  149.09 38.6125 149.225 38.7475 ;
         LAYER metal3 ;
         RECT  21.435 26.6525 21.57 26.7875 ;
         LAYER metal3 ;
         RECT  27.225 9.4375 27.36 9.5725 ;
         LAYER metal4 ;
         RECT  35.505 17.5 35.645 119.41 ;
         LAYER metal3 ;
         RECT  28.3025 0.0025 28.4375 0.1375 ;
         LAYER metal3 ;
         RECT  35.1125 125.065 130.7875 125.135 ;
         LAYER metal3 ;
         RECT  149.09 29.6425 149.225 29.7775 ;
         LAYER metal3 ;
         RECT  35.1125 10.465 130.7525 10.535 ;
         LAYER metal3 ;
         RECT  143.3 122.4675 143.435 122.6025 ;
         LAYER metal3 ;
         RECT  35.1125 14.185 132.43 14.255 ;
         LAYER metal4 ;
         RECT  168.105 102.2275 168.245 124.63 ;
         LAYER metal3 ;
         RECT  27.225 14.3775 27.36 14.5125 ;
         LAYER metal3 ;
         RECT  149.09 20.6725 149.225 20.8075 ;
         LAYER metal3 ;
         RECT  21.435 44.5925 21.57 44.7275 ;
         LAYER metal4 ;
         RECT  135.015 17.5 135.155 119.41 ;
         LAYER metal3 ;
         RECT  168.435 134.3725 168.57 134.5075 ;
         LAYER metal3 ;
         RECT  142.4175 133.1075 142.5525 133.2425 ;
         LAYER metal3 ;
         RECT  21.435 38.6125 21.57 38.7475 ;
         LAYER metal3 ;
         RECT  119.8225 0.0025 119.9575 0.1375 ;
         LAYER metal3 ;
         RECT  149.09 23.6625 149.225 23.7975 ;
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal4 ;
         RECT  164.61 119.55 164.75 134.51 ;
         LAYER metal3 ;
         RECT  149.09 44.5925 149.225 44.7275 ;
         LAYER metal4 ;
         RECT  143.94 20.6375 144.08 116.56 ;
         LAYER metal3 ;
         RECT  62.6225 0.0025 62.7575 0.1375 ;
         LAYER metal3 ;
         RECT  21.435 29.6425 21.57 29.7775 ;
         LAYER metal3 ;
         RECT  149.09 35.6225 149.225 35.7575 ;
         LAYER metal3 ;
         RECT  35.1125 122.725 132.43 122.795 ;
         LAYER metal3 ;
         RECT  39.7425 0.0025 39.8775 0.1375 ;
         LAYER metal3 ;
         RECT  74.0625 0.0025 74.1975 0.1375 ;
         LAYER metal3 ;
         RECT  21.435 32.6325 21.57 32.7675 ;
         LAYER metal3 ;
         RECT  25.4425 0.0025 25.5775 0.1375 ;
         LAYER metal3 ;
         RECT  96.9425 0.0025 97.0775 0.1375 ;
         LAYER metal3 ;
         RECT  21.435 41.6025 21.57 41.7375 ;
         LAYER metal3 ;
         RECT  131.2625 0.0025 131.3975 0.1375 ;
         LAYER metal3 ;
         RECT  21.435 23.6625 21.57 23.7975 ;
         LAYER metal3 ;
         RECT  108.3825 0.0025 108.5175 0.1375 ;
         LAYER metal3 ;
         RECT  149.09 41.6025 149.225 41.7375 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 170.855 134.37 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 170.855 134.37 ;
   LAYER  metal3 ;
      RECT  26.0 0.9675 28.445 1.3825 ;
      RECT  28.86 0.9675 31.305 1.3825 ;
      RECT  31.72 0.9675 34.165 1.3825 ;
      RECT  34.58 0.9675 37.025 1.3825 ;
      RECT  37.44 0.9675 39.885 1.3825 ;
      RECT  40.3 0.9675 42.745 1.3825 ;
      RECT  43.16 0.9675 45.605 1.3825 ;
      RECT  46.02 0.9675 48.465 1.3825 ;
      RECT  48.88 0.9675 51.325 1.3825 ;
      RECT  51.74 0.9675 54.185 1.3825 ;
      RECT  54.6 0.9675 57.045 1.3825 ;
      RECT  57.46 0.9675 59.905 1.3825 ;
      RECT  60.32 0.9675 62.765 1.3825 ;
      RECT  63.18 0.9675 65.625 1.3825 ;
      RECT  66.04 0.9675 68.485 1.3825 ;
      RECT  68.9 0.9675 71.345 1.3825 ;
      RECT  71.76 0.9675 74.205 1.3825 ;
      RECT  74.62 0.9675 77.065 1.3825 ;
      RECT  77.48 0.9675 79.925 1.3825 ;
      RECT  80.34 0.9675 82.785 1.3825 ;
      RECT  83.2 0.9675 85.645 1.3825 ;
      RECT  86.06 0.9675 88.505 1.3825 ;
      RECT  88.92 0.9675 91.365 1.3825 ;
      RECT  91.78 0.9675 94.225 1.3825 ;
      RECT  94.64 0.9675 97.085 1.3825 ;
      RECT  97.5 0.9675 99.945 1.3825 ;
      RECT  100.36 0.9675 102.805 1.3825 ;
      RECT  103.22 0.9675 105.665 1.3825 ;
      RECT  106.08 0.9675 108.525 1.3825 ;
      RECT  108.94 0.9675 111.385 1.3825 ;
      RECT  111.8 0.9675 114.245 1.3825 ;
      RECT  114.66 0.9675 117.105 1.3825 ;
      RECT  117.52 0.9675 119.965 1.3825 ;
      RECT  120.38 0.9675 122.825 1.3825 ;
      RECT  123.24 0.9675 125.685 1.3825 ;
      RECT  126.1 0.9675 128.545 1.3825 ;
      RECT  128.96 0.9675 131.405 1.3825 ;
      RECT  131.82 0.9675 134.265 1.3825 ;
      RECT  134.68 0.9675 137.125 1.3825 ;
      RECT  137.54 0.9675 170.855 1.3825 ;
      RECT  23.14 0.9675 25.585 1.3825 ;
      RECT  0.14 45.5575 17.005 45.9725 ;
      RECT  0.14 45.9725 17.005 134.37 ;
      RECT  17.005 1.3825 17.42 45.5575 ;
      RECT  17.42 45.5575 25.585 45.9725 ;
      RECT  17.42 45.9725 25.585 134.37 ;
      RECT  17.005 45.9725 17.42 48.2875 ;
      RECT  17.005 48.7025 17.42 50.4975 ;
      RECT  17.005 50.9125 17.42 53.2275 ;
      RECT  17.005 53.6425 17.42 55.4375 ;
      RECT  17.005 55.8525 17.42 58.1675 ;
      RECT  17.005 58.5825 17.42 134.37 ;
      RECT  26.0 131.8625 144.855 132.2775 ;
      RECT  144.855 132.2775 145.27 134.37 ;
      RECT  145.27 1.3825 153.435 19.4275 ;
      RECT  145.27 19.4275 153.435 19.8425 ;
      RECT  153.435 19.8425 153.85 131.8625 ;
      RECT  153.85 1.3825 170.855 19.4275 ;
      RECT  153.85 19.4275 170.855 19.8425 ;
      RECT  153.435 17.1125 153.85 19.4275 ;
      RECT  153.435 14.9025 153.85 16.6975 ;
      RECT  153.435 12.1725 153.85 14.4875 ;
      RECT  153.435 9.9625 153.85 11.7575 ;
      RECT  153.435 1.3825 153.85 6.8175 ;
      RECT  153.435 7.2325 153.85 9.5475 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  170.435 132.2775 170.85 133.1275 ;
      RECT  170.435 133.5425 170.85 134.37 ;
      RECT  170.85 132.2775 170.855 133.1275 ;
      RECT  170.85 133.1275 170.855 133.5425 ;
      RECT  170.85 133.5425 170.855 134.37 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 45.5575 ;
      RECT  6.5225 1.3825 17.005 1.4675 ;
      RECT  6.5225 1.4675 17.005 45.5575 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 22.725 1.0525 ;
      RECT  6.5225 1.0525 22.725 1.3825 ;
      RECT  145.27 132.2775 164.3325 133.0425 ;
      RECT  145.27 133.0425 164.3325 133.1275 ;
      RECT  164.3325 132.2775 164.7475 133.0425 ;
      RECT  164.7475 132.2775 170.435 133.0425 ;
      RECT  164.7475 133.0425 170.435 133.1275 ;
      RECT  145.27 133.1275 164.3325 133.4575 ;
      RECT  145.27 133.4575 164.3325 133.5425 ;
      RECT  164.3325 133.4575 164.7475 133.5425 ;
      RECT  164.7475 133.1275 170.435 133.4575 ;
      RECT  164.7475 133.4575 170.435 133.5425 ;
      RECT  26.0 129.375 38.1575 129.79 ;
      RECT  26.0 129.79 38.1575 131.8625 ;
      RECT  38.1575 129.79 38.5725 131.8625 ;
      RECT  38.5725 129.79 144.855 131.8625 ;
      RECT  38.5725 129.375 40.5075 129.79 ;
      RECT  40.9225 129.375 42.8575 129.79 ;
      RECT  43.2725 129.375 45.2075 129.79 ;
      RECT  45.6225 129.375 47.5575 129.79 ;
      RECT  47.9725 129.375 49.9075 129.79 ;
      RECT  50.3225 129.375 52.2575 129.79 ;
      RECT  52.6725 129.375 54.6075 129.79 ;
      RECT  55.0225 129.375 56.9575 129.79 ;
      RECT  57.3725 129.375 59.3075 129.79 ;
      RECT  59.7225 129.375 61.6575 129.79 ;
      RECT  62.0725 129.375 64.0075 129.79 ;
      RECT  64.4225 129.375 66.3575 129.79 ;
      RECT  66.7725 129.375 68.7075 129.79 ;
      RECT  69.1225 129.375 71.0575 129.79 ;
      RECT  71.4725 129.375 73.4075 129.79 ;
      RECT  73.8225 129.375 75.7575 129.79 ;
      RECT  76.1725 129.375 78.1075 129.79 ;
      RECT  78.5225 129.375 80.4575 129.79 ;
      RECT  80.8725 129.375 82.8075 129.79 ;
      RECT  83.2225 129.375 85.1575 129.79 ;
      RECT  85.5725 129.375 87.5075 129.79 ;
      RECT  87.9225 129.375 89.8575 129.79 ;
      RECT  90.2725 129.375 92.2075 129.79 ;
      RECT  92.6225 129.375 94.5575 129.79 ;
      RECT  94.9725 129.375 96.9075 129.79 ;
      RECT  97.3225 129.375 99.2575 129.79 ;
      RECT  99.6725 129.375 101.6075 129.79 ;
      RECT  102.0225 129.375 103.9575 129.79 ;
      RECT  104.3725 129.375 106.3075 129.79 ;
      RECT  106.7225 129.375 108.6575 129.79 ;
      RECT  109.0725 129.375 111.0075 129.79 ;
      RECT  111.4225 129.375 113.3575 129.79 ;
      RECT  113.7725 129.375 115.7075 129.79 ;
      RECT  116.1225 129.375 118.0575 129.79 ;
      RECT  118.4725 129.375 120.4075 129.79 ;
      RECT  120.8225 129.375 122.7575 129.79 ;
      RECT  123.1725 129.375 125.1075 129.79 ;
      RECT  125.5225 129.375 127.4575 129.79 ;
      RECT  127.8725 129.375 129.8075 129.79 ;
      RECT  130.2225 129.375 144.855 129.79 ;
      RECT  38.5725 1.3825 82.5025 2.3325 ;
      RECT  82.5025 1.3825 82.9175 2.3325 ;
      RECT  82.9175 1.3825 144.855 2.3325 ;
      RECT  71.4775 2.3325 82.5025 2.7475 ;
      RECT  26.0 19.825 28.995 20.24 ;
      RECT  26.0 20.24 28.995 129.375 ;
      RECT  28.995 1.3825 29.41 19.825 ;
      RECT  28.995 20.24 29.41 129.375 ;
      RECT  29.41 19.825 38.1575 20.24 ;
      RECT  17.42 30.9975 22.8225 31.4125 ;
      RECT  23.2375 30.9975 25.585 31.4125 ;
      RECT  23.2375 31.4125 25.585 45.5575 ;
      RECT  38.1575 1.3825 38.5725 8.275 ;
      RECT  38.5725 2.7475 82.5025 8.275 ;
      RECT  82.5025 2.7475 82.9175 8.275 ;
      RECT  82.9175 2.7475 130.8925 8.275 ;
      RECT  130.8925 2.7475 144.855 8.275 ;
      RECT  130.8925 8.275 144.855 8.625 ;
      RECT  29.41 1.3825 34.9725 8.275 ;
      RECT  29.41 8.275 34.9725 8.625 ;
      RECT  145.27 19.8425 147.4225 25.0175 ;
      RECT  145.27 25.0175 147.4225 25.4325 ;
      RECT  147.8375 25.0175 153.435 25.4325 ;
      RECT  147.4225 43.3725 147.8375 131.8625 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 45.5575 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 45.5575 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 45.5575 ;
      RECT  22.8225 43.3725 23.2375 45.5575 ;
      RECT  26.0 1.3825 27.085 11.7675 ;
      RECT  26.0 11.7675 27.085 12.1825 ;
      RECT  26.0 12.1825 27.085 19.825 ;
      RECT  27.5 1.3825 28.995 11.7675 ;
      RECT  27.5 11.7675 28.995 12.1825 ;
      RECT  27.5 12.1825 28.995 19.825 ;
      RECT  29.41 20.24 34.9725 126.8175 ;
      RECT  29.41 126.8175 34.9725 127.1675 ;
      RECT  29.41 127.1675 34.9725 129.375 ;
      RECT  34.9725 127.1675 38.1575 129.375 ;
      RECT  38.1575 127.1675 38.5725 129.375 ;
      RECT  38.5725 127.1675 82.5025 129.375 ;
      RECT  82.5025 127.1675 82.9175 129.375 ;
      RECT  82.9175 127.1675 130.8925 129.375 ;
      RECT  22.8225 31.4125 23.2375 33.9875 ;
      RECT  130.8925 116.92 141.25 117.335 ;
      RECT  141.25 8.625 141.665 116.92 ;
      RECT  141.25 117.335 141.665 129.375 ;
      RECT  141.665 8.625 144.855 116.92 ;
      RECT  141.665 116.92 144.855 117.335 ;
      RECT  34.9725 20.24 38.1575 119.965 ;
      RECT  130.8925 117.335 133.7125 119.965 ;
      RECT  133.7125 119.965 141.25 120.315 ;
      RECT  133.7125 120.315 141.25 129.375 ;
      RECT  17.42 1.3825 22.4425 2.3325 ;
      RECT  17.42 2.3325 22.4425 2.7475 ;
      RECT  22.4425 1.3825 22.8225 2.3325 ;
      RECT  22.4425 2.7475 22.8225 30.9975 ;
      RECT  22.8225 1.3825 22.8575 2.3325 ;
      RECT  22.8225 2.7475 22.8575 22.0275 ;
      RECT  22.8575 1.3825 23.2375 2.3325 ;
      RECT  22.8575 2.3325 23.2375 2.7475 ;
      RECT  22.8575 2.7475 23.2375 22.0275 ;
      RECT  145.27 131.8625 168.295 132.1775 ;
      RECT  145.27 132.1775 168.295 132.2775 ;
      RECT  168.295 132.1775 168.71 132.2775 ;
      RECT  168.71 131.8625 170.855 132.1775 ;
      RECT  168.71 132.1775 170.855 132.2775 ;
      RECT  153.85 19.8425 168.295 131.7625 ;
      RECT  153.85 131.7625 168.295 131.8625 ;
      RECT  168.295 19.8425 168.71 131.7625 ;
      RECT  168.71 19.8425 170.855 131.7625 ;
      RECT  168.71 131.7625 170.855 131.8625 ;
      RECT  144.855 1.3825 145.1375 130.4975 ;
      RECT  144.855 130.4975 145.1375 130.9125 ;
      RECT  144.855 130.9125 145.1375 131.8625 ;
      RECT  145.1375 1.3825 145.27 130.4975 ;
      RECT  145.1375 130.9125 145.27 131.8625 ;
      RECT  145.27 25.4325 145.5525 130.4975 ;
      RECT  145.27 130.9125 145.5525 131.8625 ;
      RECT  145.5525 25.4325 147.4225 130.4975 ;
      RECT  145.5525 130.4975 147.4225 130.9125 ;
      RECT  145.5525 130.9125 147.4225 131.8625 ;
      RECT  25.585 1.3825 25.7175 2.3325 ;
      RECT  25.585 2.7475 25.7175 134.37 ;
      RECT  25.7175 1.3825 26.0 2.3325 ;
      RECT  25.7175 2.3325 26.0 2.7475 ;
      RECT  25.7175 2.7475 26.0 134.37 ;
      RECT  23.2375 1.3825 25.3025 2.3325 ;
      RECT  23.2375 2.3325 25.3025 2.7475 ;
      RECT  23.2375 2.7475 25.3025 30.9975 ;
      RECT  25.3025 1.3825 25.585 2.3325 ;
      RECT  25.3025 2.7475 25.585 30.9975 ;
      RECT  147.4225 19.8425 147.8375 22.0275 ;
      RECT  147.4225 22.4425 147.8375 25.0175 ;
      RECT  29.41 8.625 33.8275 19.0375 ;
      RECT  29.41 19.0375 33.8275 19.4525 ;
      RECT  29.41 19.4525 33.8275 19.825 ;
      RECT  33.8275 8.625 34.2425 19.0375 ;
      RECT  33.8275 19.4525 34.2425 19.825 ;
      RECT  34.2425 8.625 34.9725 19.0375 ;
      RECT  34.2425 19.0375 34.9725 19.4525 ;
      RECT  34.2425 19.4525 34.9725 19.825 ;
      RECT  82.9175 2.3325 93.9425 2.7475 ;
      RECT  22.8225 22.4425 23.2375 25.0175 ;
      RECT  22.8225 25.4325 23.2375 30.9975 ;
      RECT  147.4225 40.3825 147.8375 42.9575 ;
      RECT  38.5725 2.3325 48.1825 2.7475 ;
      RECT  22.8225 34.4025 23.2375 39.9675 ;
      RECT  22.8225 40.3825 23.2375 42.9575 ;
      RECT  147.4225 34.4025 147.8375 39.9675 ;
      RECT  48.5975 2.3325 59.6225 2.7475 ;
      RECT  60.0375 2.3325 71.0625 2.7475 ;
      RECT  117.2375 2.3325 128.2625 2.7475 ;
      RECT  128.6775 2.3325 144.855 2.7475 ;
      RECT  34.9725 1.3825 36.7425 2.3325 ;
      RECT  34.9725 2.3325 36.7425 2.7475 ;
      RECT  34.9725 2.7475 36.7425 8.275 ;
      RECT  36.7425 1.3825 37.1575 2.3325 ;
      RECT  36.7425 2.7475 37.1575 8.275 ;
      RECT  37.1575 1.3825 38.1575 2.3325 ;
      RECT  37.1575 2.3325 38.1575 2.7475 ;
      RECT  37.1575 2.7475 38.1575 8.275 ;
      RECT  147.4225 25.4325 147.8375 30.9975 ;
      RECT  147.4225 31.4125 147.8375 33.9875 ;
      RECT  141.665 117.335 143.16 124.7975 ;
      RECT  141.665 124.7975 143.16 125.2125 ;
      RECT  141.665 125.2125 143.16 129.375 ;
      RECT  143.575 117.335 144.855 124.7975 ;
      RECT  143.575 124.7975 144.855 125.2125 ;
      RECT  143.575 125.2125 144.855 129.375 ;
      RECT  94.3575 2.3325 105.3825 2.7475 ;
      RECT  105.7975 2.3325 116.8225 2.7475 ;
      RECT  34.9725 17.015 38.1575 19.825 ;
      RECT  130.8925 17.015 132.5375 116.92 ;
      RECT  132.5375 16.665 141.25 17.015 ;
      RECT  132.5375 17.015 141.25 116.92 ;
      RECT  38.1575 17.015 38.5725 119.965 ;
      RECT  38.5725 17.015 82.5025 119.965 ;
      RECT  82.5025 17.015 82.9175 119.965 ;
      RECT  82.9175 17.015 130.8925 119.965 ;
      RECT  133.7125 117.335 136.4175 117.7075 ;
      RECT  133.7125 117.7075 136.4175 118.1225 ;
      RECT  133.7125 118.1225 136.4175 119.965 ;
      RECT  136.4175 117.335 136.8325 117.7075 ;
      RECT  136.4175 118.1225 136.8325 119.965 ;
      RECT  136.8325 117.335 141.25 117.7075 ;
      RECT  136.8325 117.7075 141.25 118.1225 ;
      RECT  136.8325 118.1225 141.25 119.965 ;
      RECT  17.42 31.4125 21.295 35.4825 ;
      RECT  17.42 35.4825 21.295 35.8975 ;
      RECT  17.42 35.8975 21.295 45.5575 ;
      RECT  21.71 31.4125 22.8225 35.4825 ;
      RECT  21.71 35.4825 22.8225 35.8975 ;
      RECT  21.71 35.8975 22.8225 45.5575 ;
      RECT  147.8375 25.4325 148.95 32.4925 ;
      RECT  147.8375 32.4925 148.95 32.9075 ;
      RECT  147.8375 32.9075 148.95 131.8625 ;
      RECT  149.365 25.4325 153.435 32.4925 ;
      RECT  149.365 32.4925 153.435 32.9075 ;
      RECT  149.365 32.9075 153.435 131.8625 ;
      RECT  143.16 125.2125 143.575 127.2675 ;
      RECT  143.16 127.6825 143.575 129.375 ;
      RECT  148.95 25.4325 149.365 26.5125 ;
      RECT  26.0 0.2775 51.0425 0.9675 ;
      RECT  51.0425 0.2775 51.4575 0.9675 ;
      RECT  51.4575 0.2775 170.855 0.9675 ;
      RECT  17.42 2.7475 21.295 20.5325 ;
      RECT  17.42 20.5325 21.295 20.9475 ;
      RECT  17.42 20.9475 21.295 30.9975 ;
      RECT  21.295 2.7475 21.71 20.5325 ;
      RECT  21.71 2.7475 22.4425 20.5325 ;
      RECT  21.71 20.5325 22.4425 20.9475 ;
      RECT  21.71 20.9475 22.4425 30.9975 ;
      RECT  27.085 1.3825 27.5 9.2975 ;
      RECT  27.085 9.7125 27.5 11.7675 ;
      RECT  26.0 0.14 28.1625 0.2775 ;
      RECT  34.9725 125.275 38.1575 126.8175 ;
      RECT  38.1575 125.275 38.5725 126.8175 ;
      RECT  38.5725 125.275 82.5025 126.8175 ;
      RECT  82.5025 125.275 82.9175 126.8175 ;
      RECT  82.9175 125.275 130.8925 126.8175 ;
      RECT  130.8925 125.275 130.9275 129.375 ;
      RECT  130.9275 124.925 133.7125 125.275 ;
      RECT  130.9275 125.275 133.7125 129.375 ;
      RECT  148.95 26.9275 149.365 29.5025 ;
      RECT  148.95 29.9175 149.365 32.4925 ;
      RECT  34.9725 8.625 38.1575 10.325 ;
      RECT  38.1575 8.625 38.5725 10.325 ;
      RECT  38.5725 8.625 82.5025 10.325 ;
      RECT  82.5025 8.625 82.9175 10.325 ;
      RECT  82.9175 8.625 130.8925 10.325 ;
      RECT  143.16 117.335 143.575 122.3275 ;
      RECT  143.16 122.7425 143.575 124.7975 ;
      RECT  130.8925 8.625 132.5375 14.045 ;
      RECT  130.8925 14.395 132.5375 16.665 ;
      RECT  132.5375 8.625 132.57 14.045 ;
      RECT  132.5375 14.395 132.57 16.665 ;
      RECT  132.57 8.625 141.25 14.045 ;
      RECT  132.57 14.045 141.25 14.395 ;
      RECT  132.57 14.395 141.25 16.665 ;
      RECT  34.9725 10.675 38.1575 14.045 ;
      RECT  34.9725 14.395 38.1575 16.665 ;
      RECT  38.1575 10.675 38.5725 14.045 ;
      RECT  38.1575 14.395 38.5725 16.665 ;
      RECT  38.5725 10.675 82.5025 14.045 ;
      RECT  38.5725 14.395 82.5025 16.665 ;
      RECT  82.5025 10.675 82.9175 14.045 ;
      RECT  82.5025 14.395 82.9175 16.665 ;
      RECT  82.9175 10.675 130.8925 14.045 ;
      RECT  82.9175 14.395 130.8925 16.665 ;
      RECT  27.085 12.1825 27.5 14.2375 ;
      RECT  27.085 14.6525 27.5 19.825 ;
      RECT  147.8375 19.8425 148.95 20.5325 ;
      RECT  147.8375 20.5325 148.95 20.9475 ;
      RECT  147.8375 20.9475 148.95 25.0175 ;
      RECT  148.95 19.8425 149.365 20.5325 ;
      RECT  149.365 19.8425 153.435 20.5325 ;
      RECT  149.365 20.5325 153.435 20.9475 ;
      RECT  149.365 20.9475 153.435 25.0175 ;
      RECT  21.295 44.8675 21.71 45.5575 ;
      RECT  145.27 133.5425 168.295 134.2325 ;
      RECT  145.27 134.2325 168.295 134.37 ;
      RECT  168.295 133.5425 168.71 134.2325 ;
      RECT  168.71 133.5425 170.435 134.2325 ;
      RECT  168.71 134.2325 170.435 134.37 ;
      RECT  26.0 132.2775 142.2775 132.9675 ;
      RECT  26.0 132.9675 142.2775 133.3825 ;
      RECT  26.0 133.3825 142.2775 134.37 ;
      RECT  142.2775 132.2775 142.6925 132.9675 ;
      RECT  142.2775 133.3825 142.6925 134.37 ;
      RECT  142.6925 132.2775 144.855 132.9675 ;
      RECT  142.6925 132.9675 144.855 133.3825 ;
      RECT  142.6925 133.3825 144.855 134.37 ;
      RECT  21.295 35.8975 21.71 38.4725 ;
      RECT  148.95 20.9475 149.365 23.5225 ;
      RECT  148.95 23.9375 149.365 25.0175 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  0.14 0.2775 2.285 0.9675 ;
      RECT  2.285 0.2775 2.7 0.9675 ;
      RECT  2.7 0.2775 25.585 0.9675 ;
      RECT  148.95 44.8675 149.365 131.8625 ;
      RECT  51.4575 0.14 62.4825 0.2775 ;
      RECT  21.295 26.9275 21.71 29.5025 ;
      RECT  21.295 29.9175 21.71 30.9975 ;
      RECT  148.95 32.9075 149.365 35.4825 ;
      RECT  148.95 35.8975 149.365 38.4725 ;
      RECT  34.9725 120.315 38.1575 122.585 ;
      RECT  34.9725 122.935 38.1575 124.925 ;
      RECT  38.1575 120.315 38.5725 122.585 ;
      RECT  38.1575 122.935 38.5725 124.925 ;
      RECT  38.5725 120.315 82.5025 122.585 ;
      RECT  38.5725 122.935 82.5025 124.925 ;
      RECT  82.5025 120.315 82.9175 122.585 ;
      RECT  82.5025 122.935 82.9175 124.925 ;
      RECT  82.9175 120.315 130.8925 122.585 ;
      RECT  82.9175 122.935 130.8925 124.925 ;
      RECT  130.8925 120.315 130.9275 122.585 ;
      RECT  130.8925 122.935 130.9275 124.925 ;
      RECT  130.9275 120.315 132.57 122.585 ;
      RECT  130.9275 122.935 132.57 124.925 ;
      RECT  132.57 120.315 133.7125 122.585 ;
      RECT  132.57 122.585 133.7125 122.935 ;
      RECT  132.57 122.935 133.7125 124.925 ;
      RECT  28.5775 0.14 39.6025 0.2775 ;
      RECT  40.0175 0.14 51.0425 0.2775 ;
      RECT  62.8975 0.14 73.9225 0.2775 ;
      RECT  74.3375 0.14 85.3625 0.2775 ;
      RECT  21.295 31.4125 21.71 32.4925 ;
      RECT  21.295 32.9075 21.71 35.4825 ;
      RECT  25.585 0.2775 25.7175 0.9675 ;
      RECT  25.7175 0.14 26.0 0.2775 ;
      RECT  25.7175 0.2775 26.0 0.9675 ;
      RECT  2.7 0.14 25.3025 0.2775 ;
      RECT  85.7775 0.14 96.8025 0.2775 ;
      RECT  21.295 38.8875 21.71 41.4625 ;
      RECT  21.295 41.8775 21.71 44.4525 ;
      RECT  120.0975 0.14 131.1225 0.2775 ;
      RECT  131.5375 0.14 170.855 0.2775 ;
      RECT  21.295 20.9475 21.71 23.5225 ;
      RECT  21.295 23.9375 21.71 26.5125 ;
      RECT  97.2175 0.14 108.2425 0.2775 ;
      RECT  108.6575 0.14 119.6825 0.2775 ;
      RECT  148.95 38.8875 149.365 41.4625 ;
      RECT  148.95 41.8775 149.365 44.4525 ;
   LAYER  metal4 ;
      RECT  141.725 116.84 142.425 134.37 ;
      RECT  169.8875 20.39 170.5875 101.98 ;
      RECT  170.5875 20.39 170.855 101.98 ;
      RECT  170.5875 101.98 170.855 116.84 ;
      RECT  169.8875 124.9425 170.5875 134.37 ;
      RECT  170.5875 116.84 170.855 124.9425 ;
      RECT  170.5875 124.9425 170.855 134.37 ;
      RECT  34.765 0.14 35.465 17.22 ;
      RECT  35.465 0.14 141.725 17.22 ;
      RECT  0.14 116.84 34.765 119.69 ;
      RECT  0.14 119.69 34.765 134.37 ;
      RECT  34.765 119.69 35.465 134.37 ;
      RECT  35.465 119.69 141.725 134.37 ;
      RECT  0.14 44.31 16.58 59.83 ;
      RECT  0.14 59.83 16.58 116.84 ;
      RECT  16.58 20.39 17.28 44.31 ;
      RECT  16.58 59.83 17.28 116.84 ;
      RECT  135.895 116.84 141.725 119.69 ;
      RECT  135.895 20.39 136.275 116.77 ;
      RECT  135.895 116.77 136.275 116.84 ;
      RECT  136.275 116.77 136.975 116.84 ;
      RECT  19.3 0.14 20.0 2.19 ;
      RECT  20.0 0.14 34.765 2.19 ;
      RECT  20.0 2.19 34.765 17.22 ;
      RECT  19.3 17.71 20.0 20.39 ;
      RECT  20.0 17.22 34.765 17.71 ;
      RECT  0.14 20.39 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 44.31 ;
      RECT  0.4075 32.53 1.1075 44.31 ;
      RECT  0.14 2.19 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 17.22 ;
      RECT  0.4075 2.19 1.1075 9.5675 ;
      RECT  0.14 17.22 0.4075 17.71 ;
      RECT  0.14 17.71 0.4075 20.39 ;
      RECT  142.425 116.84 150.855 121.74 ;
      RECT  142.425 121.74 150.855 124.9425 ;
      RECT  150.855 116.84 151.555 121.74 ;
      RECT  142.425 124.9425 150.855 132.32 ;
      RECT  142.425 132.32 150.855 134.37 ;
      RECT  150.855 132.32 151.555 134.37 ;
      RECT  153.575 0.14 154.275 5.57 ;
      RECT  154.275 0.14 170.855 5.57 ;
      RECT  154.275 5.57 170.855 20.39 ;
      RECT  153.575 21.09 154.275 101.98 ;
      RECT  154.275 20.39 169.8875 21.09 ;
      RECT  34.385 20.39 34.765 44.31 ;
      RECT  34.385 44.31 34.765 59.83 ;
      RECT  33.685 116.77 34.385 116.84 ;
      RECT  34.385 59.83 34.765 116.77 ;
      RECT  34.385 116.77 34.765 116.84 ;
      RECT  0.14 0.14 5.825 2.19 ;
      RECT  6.525 0.14 19.3 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 19.3 9.5675 ;
      RECT  5.825 15.24 6.525 17.22 ;
      RECT  6.525 9.5675 19.3 15.24 ;
      RECT  6.525 15.24 19.3 17.22 ;
      RECT  142.425 0.14 150.715 5.505 ;
      RECT  142.425 5.505 150.715 5.57 ;
      RECT  150.715 0.14 151.415 5.505 ;
      RECT  151.415 0.14 153.575 5.505 ;
      RECT  151.415 5.505 153.575 5.57 ;
      RECT  151.415 5.57 153.575 20.39 ;
      RECT  151.415 20.39 153.575 21.09 ;
      RECT  150.715 21.155 151.415 101.98 ;
      RECT  151.415 21.09 153.575 21.155 ;
      RECT  151.415 21.155 153.575 101.98 ;
      RECT  141.725 0.14 141.865 20.3575 ;
      RECT  141.865 0.14 142.425 20.3575 ;
      RECT  141.865 20.3575 142.425 20.39 ;
      RECT  135.895 17.22 141.165 20.3575 ;
      RECT  135.895 20.3575 141.165 20.39 ;
      RECT  141.165 17.22 141.725 20.3575 ;
      RECT  136.975 20.39 141.165 116.77 ;
      RECT  136.975 116.77 141.165 116.8025 ;
      RECT  136.975 116.8025 141.165 116.84 ;
      RECT  141.165 116.8025 141.725 116.84 ;
      RECT  17.28 20.39 19.44 44.245 ;
      RECT  17.28 44.245 19.44 44.31 ;
      RECT  19.44 20.39 20.14 44.245 ;
      RECT  17.28 44.31 19.44 59.83 ;
      RECT  17.28 59.83 19.44 59.895 ;
      RECT  17.28 59.895 19.44 116.84 ;
      RECT  19.44 59.895 20.14 116.84 ;
      RECT  20.0 17.71 28.795 20.3575 ;
      RECT  28.795 17.71 29.495 20.3575 ;
      RECT  29.495 17.71 34.765 20.3575 ;
      RECT  29.495 20.3575 34.765 20.39 ;
      RECT  29.495 20.39 33.685 44.31 ;
      RECT  29.495 44.31 33.685 59.83 ;
      RECT  29.495 59.83 33.685 116.77 ;
      RECT  28.935 116.8025 29.495 116.84 ;
      RECT  29.495 116.77 33.685 116.8025 ;
      RECT  29.495 116.8025 33.685 116.84 ;
      RECT  1.1075 20.39 2.47 32.53 ;
      RECT  3.17 20.39 16.58 32.53 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 44.31 ;
      RECT  2.47 32.5625 3.17 44.31 ;
      RECT  3.17 32.53 16.58 32.5625 ;
      RECT  3.17 32.5625 16.58 44.31 ;
      RECT  1.1075 17.22 2.47 17.71 ;
      RECT  3.17 17.22 19.3 17.71 ;
      RECT  1.1075 17.71 2.47 20.39 ;
      RECT  3.17 17.71 19.3 20.39 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 15.24 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  1.1075 15.24 2.47 17.22 ;
      RECT  3.17 15.24 5.825 17.22 ;
      RECT  20.14 20.39 26.3 44.245 ;
      RECT  27.0 20.39 28.235 44.245 ;
      RECT  20.14 44.245 26.3 44.31 ;
      RECT  27.0 44.245 28.235 44.31 ;
      RECT  20.14 44.31 26.3 59.83 ;
      RECT  27.0 44.31 28.235 59.83 ;
      RECT  20.14 59.83 26.3 59.895 ;
      RECT  27.0 59.83 28.235 59.895 ;
      RECT  20.14 59.895 26.3 116.84 ;
      RECT  27.0 59.895 28.235 116.84 ;
      RECT  20.0 20.3575 26.3 20.39 ;
      RECT  27.0 20.3575 28.795 20.39 ;
      RECT  168.525 101.98 169.8875 116.84 ;
      RECT  168.525 116.84 169.8875 121.74 ;
      RECT  167.825 124.91 168.525 124.9425 ;
      RECT  168.525 121.74 169.8875 124.91 ;
      RECT  168.525 124.91 169.8875 124.9425 ;
      RECT  154.275 21.09 167.825 101.9475 ;
      RECT  154.275 101.9475 167.825 101.98 ;
      RECT  167.825 21.09 168.525 101.9475 ;
      RECT  168.525 21.09 169.8875 101.9475 ;
      RECT  168.525 101.9475 169.8875 101.98 ;
      RECT  35.925 17.22 134.735 20.39 ;
      RECT  35.925 20.39 134.735 116.84 ;
      RECT  35.925 116.84 134.735 119.69 ;
      RECT  151.555 124.9425 164.33 132.32 ;
      RECT  165.03 124.9425 169.8875 132.32 ;
      RECT  151.555 132.32 164.33 134.37 ;
      RECT  165.03 132.32 169.8875 134.37 ;
      RECT  151.555 116.84 164.33 119.27 ;
      RECT  151.555 119.27 164.33 121.74 ;
      RECT  164.33 116.84 165.03 119.27 ;
      RECT  165.03 116.84 167.825 119.27 ;
      RECT  165.03 119.27 167.825 121.74 ;
      RECT  151.555 121.74 164.33 124.91 ;
      RECT  165.03 121.74 167.825 124.91 ;
      RECT  151.555 124.91 164.33 124.9425 ;
      RECT  165.03 124.91 167.825 124.9425 ;
      RECT  142.425 5.57 143.66 20.3575 ;
      RECT  142.425 20.3575 143.66 20.39 ;
      RECT  143.66 5.57 144.36 20.3575 ;
      RECT  144.36 5.57 150.715 20.3575 ;
      RECT  144.36 20.3575 150.715 20.39 ;
      RECT  142.425 20.39 143.66 21.09 ;
      RECT  144.36 20.39 150.715 21.09 ;
      RECT  142.425 21.09 143.66 21.155 ;
      RECT  144.36 21.09 150.715 21.155 ;
      RECT  142.425 21.155 143.66 101.98 ;
      RECT  144.36 21.155 150.715 101.98 ;
      RECT  142.425 101.98 143.66 116.84 ;
      RECT  144.36 101.98 167.825 116.84 ;
   END
END    freepdk45_sram_1w1r_128x40
END    LIBRARY
