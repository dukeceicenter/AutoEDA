VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_12x256
   CLASS BLOCK ;
   SIZE 120.195 BY 136.265 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.36 1.105 23.495 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.22 1.105 26.355 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.08 1.105 29.215 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.94 1.105 32.075 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.8 1.105 34.935 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.66 1.105 37.795 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.52 1.105 40.655 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.38 1.105 43.515 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.24 1.105 46.375 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.1 1.105 49.235 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.96 1.105 52.095 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.82 1.105 54.955 1.24 ;
      END
   END din0[11]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.64 1.105 17.775 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.5 1.105 20.635 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 46.08 12.055 46.215 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 48.81 12.055 48.945 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 51.02 12.055 51.155 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 53.75 12.055 53.885 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 55.96 12.055 56.095 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 58.69 12.055 58.825 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.42 135.025 99.555 135.16 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.56 135.025 96.695 135.16 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.0 19.95 108.135 20.085 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.0 17.22 108.135 17.355 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.0 15.01 108.135 15.145 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.0 12.28 108.135 12.415 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.0 10.07 108.135 10.205 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.0 7.34 108.135 7.475 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.49 0.42 1.625 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.775 133.65 119.91 133.785 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.575 6.3825 1.71 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.6725 133.565 113.8075 133.7 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.6975 130.1575 31.8325 130.2925 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.3975 130.1575 36.5325 130.2925 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.0975 130.1575 41.2325 130.2925 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.7975 130.1575 45.9325 130.2925 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.4975 130.1575 50.6325 130.2925 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.1975 130.1575 55.3325 130.2925 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.8975 130.1575 60.0325 130.2925 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.5975 130.1575 64.7325 130.2925 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.2975 130.1575 69.4325 130.2925 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.9975 130.1575 74.1325 130.2925 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.6975 130.1575 78.8325 130.2925 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.3975 130.1575 83.5325 130.2925 ;
      END
   END dout1[11]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  92.355 21.0525 92.495 116.8725 ;
         LAYER metal3 ;
         RECT  17.7375 40.49 17.8725 40.625 ;
         LAYER metal4 ;
         RECT  119.3675 102.6425 119.5075 125.045 ;
         LAYER metal3 ;
         RECT  17.3575 2.47 17.4925 2.605 ;
         LAYER metal4 ;
         RECT  21.445 4.845 21.585 14.865 ;
         LAYER metal3 ;
         RECT  101.9875 25.54 102.1225 25.675 ;
         LAYER metal4 ;
         RECT  11.635 44.9725 11.775 59.9325 ;
         LAYER metal3 ;
         RECT  17.7375 43.48 17.8725 43.615 ;
         LAYER metal3 ;
         RECT  23.0775 2.47 23.2125 2.605 ;
         LAYER metal3 ;
         RECT  28.5125 8.5375 84.2025 8.6075 ;
         LAYER metal3 ;
         RECT  101.9875 34.51 102.1225 34.645 ;
         LAYER metal4 ;
         RECT  96.43 21.0525 96.57 116.9425 ;
         LAYER metal3 ;
         RECT  28.5125 127.6 84.2025 127.67 ;
         LAYER metal4 ;
         RECT  91.275 17.8825 91.415 119.7925 ;
         LAYER metal3 ;
         RECT  28.5125 17.1875 88.1975 17.2575 ;
         LAYER metal3 ;
         RECT  95.815 117.4425 95.95 117.5775 ;
         LAYER metal3 ;
         RECT  101.9875 22.55 102.1225 22.685 ;
         LAYER metal3 ;
         RECT  17.7375 22.55 17.8725 22.685 ;
         LAYER metal3 ;
         RECT  17.7375 31.52 17.8725 31.655 ;
         LAYER metal3 ;
         RECT  101.9875 43.48 102.1225 43.615 ;
         LAYER metal3 ;
         RECT  117.635 132.285 117.77 132.42 ;
         LAYER metal3 ;
         RECT  34.5175 2.47 34.6525 2.605 ;
         LAYER metal3 ;
         RECT  28.5125 120.4875 89.3725 120.5575 ;
         LAYER metal4 ;
         RECT  105.56 122.4025 105.7 132.4225 ;
         LAYER metal3 ;
         RECT  101.9875 31.52 102.1225 31.655 ;
         LAYER metal3 ;
         RECT  99.7025 133.66 99.8375 133.795 ;
         LAYER metal4 ;
         RECT  27.365 21.0525 27.505 116.8725 ;
         LAYER metal4 ;
         RECT  98.275 122.88 98.415 132.9 ;
         LAYER metal3 ;
         RECT  23.91 20.3475 24.045 20.4825 ;
         LAYER metal3 ;
         RECT  27.3675 19.56 27.5025 19.695 ;
         LAYER metal4 ;
         RECT  28.445 17.8825 28.585 119.7925 ;
         LAYER metal3 ;
         RECT  2.425 2.855 2.56 2.99 ;
         LAYER metal3 ;
         RECT  45.9575 2.47 46.0925 2.605 ;
         LAYER metal3 ;
         RECT  17.7375 34.51 17.8725 34.645 ;
         LAYER metal3 ;
         RECT  92.3575 118.23 92.4925 118.365 ;
         LAYER metal4 ;
         RECT  0.6875 10.23 0.8275 32.6325 ;
         LAYER metal4 ;
         RECT  108.28 6.2325 108.42 21.1925 ;
         LAYER metal3 ;
         RECT  101.9875 40.49 102.1225 40.625 ;
         LAYER metal3 ;
         RECT  17.7375 25.54 17.8725 25.675 ;
         LAYER metal4 ;
         RECT  14.355 2.8525 14.495 17.8125 ;
         LAYER metal4 ;
         RECT  23.29 21.0525 23.43 116.9425 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  28.5125 14.5675 88.23 14.6375 ;
         LAYER metal3 ;
         RECT  16.21 38.995 16.345 39.13 ;
         LAYER metal4 ;
         RECT  95.87 21.02 96.01 116.905 ;
         LAYER metal3 ;
         RECT  16.21 30.025 16.345 30.16 ;
         LAYER metal4 ;
         RECT  90.815 17.8825 90.955 119.7925 ;
         LAYER metal4 ;
         RECT  2.75 10.2625 2.89 32.665 ;
         LAYER metal3 ;
         RECT  16.21 44.975 16.345 45.11 ;
         LAYER metal3 ;
         RECT  28.5125 125.7075 84.2375 125.7775 ;
         LAYER metal3 ;
         RECT  103.515 21.055 103.65 21.19 ;
         LAYER metal3 ;
         RECT  96.8425 136.13 96.9775 136.265 ;
         LAYER metal3 ;
         RECT  103.515 44.975 103.65 45.11 ;
         LAYER metal3 ;
         RECT  117.635 134.755 117.77 134.89 ;
         LAYER metal3 ;
         RECT  25.9375 0.0 26.0725 0.135 ;
         LAYER metal4 ;
         RECT  6.105 0.3825 6.245 15.3425 ;
         LAYER metal3 ;
         RECT  28.5125 123.1075 88.23 123.1775 ;
         LAYER metal4 ;
         RECT  14.495 44.9075 14.635 59.9975 ;
         LAYER metal4 ;
         RECT  105.42 6.1675 105.56 21.2575 ;
         LAYER metal4 ;
         RECT  98.365 21.02 98.505 116.9425 ;
         LAYER metal4 ;
         RECT  21.355 21.02 21.495 116.9425 ;
         LAYER metal3 ;
         RECT  48.8175 0.0 48.9525 0.135 ;
         LAYER metal4 ;
         RECT  99.9375 122.8125 100.0775 132.9675 ;
         LAYER metal4 ;
         RECT  28.905 17.8825 29.045 119.7925 ;
         LAYER metal3 ;
         RECT  37.3775 0.0 37.5125 0.135 ;
         LAYER metal3 ;
         RECT  28.5125 10.5875 84.2025 10.6575 ;
         LAYER metal3 ;
         RECT  16.21 33.015 16.345 33.15 ;
         LAYER metal3 ;
         RECT  103.515 41.985 103.65 42.12 ;
         LAYER metal3 ;
         RECT  103.515 24.045 103.65 24.18 ;
         LAYER metal3 ;
         RECT  16.21 27.035 16.345 27.17 ;
         LAYER metal4 ;
         RECT  23.85 21.02 23.99 116.905 ;
         LAYER metal3 ;
         RECT  103.515 38.995 103.65 39.13 ;
         LAYER metal3 ;
         RECT  16.21 36.005 16.345 36.14 ;
         LAYER metal3 ;
         RECT  103.515 27.035 103.65 27.17 ;
         LAYER metal3 ;
         RECT  20.2175 0.0 20.3525 0.135 ;
         LAYER metal3 ;
         RECT  103.515 30.025 103.65 30.16 ;
         LAYER metal3 ;
         RECT  2.425 0.385 2.56 0.52 ;
         LAYER metal3 ;
         RECT  103.515 33.015 103.65 33.15 ;
         LAYER metal3 ;
         RECT  16.21 41.985 16.345 42.12 ;
         LAYER metal3 ;
         RECT  103.515 36.005 103.65 36.14 ;
         LAYER metal4 ;
         RECT  19.7825 4.7775 19.9225 14.9325 ;
         LAYER metal4 ;
         RECT  117.305 102.61 117.445 125.0125 ;
         LAYER metal3 ;
         RECT  16.21 24.045 16.345 24.18 ;
         LAYER metal3 ;
         RECT  16.21 21.055 16.345 21.19 ;
         LAYER metal4 ;
         RECT  113.81 119.9325 113.95 134.8925 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 120.055 136.125 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 120.055 136.125 ;
   LAYER  metal3 ;
      RECT  23.22 0.14 23.635 0.965 ;
      RECT  23.635 0.965 26.08 1.38 ;
      RECT  26.495 0.965 28.94 1.38 ;
      RECT  29.355 0.965 31.8 1.38 ;
      RECT  32.215 0.965 34.66 1.38 ;
      RECT  35.075 0.965 37.52 1.38 ;
      RECT  37.935 0.965 40.38 1.38 ;
      RECT  40.795 0.965 43.24 1.38 ;
      RECT  43.655 0.965 46.1 1.38 ;
      RECT  46.515 0.965 48.96 1.38 ;
      RECT  49.375 0.965 51.82 1.38 ;
      RECT  52.235 0.965 54.68 1.38 ;
      RECT  55.095 0.965 120.055 1.38 ;
      RECT  17.915 0.965 20.36 1.38 ;
      RECT  20.775 0.965 23.22 1.38 ;
      RECT  0.14 45.94 11.78 46.355 ;
      RECT  0.14 46.355 11.78 136.125 ;
      RECT  11.78 1.38 12.195 45.94 ;
      RECT  12.195 45.94 23.22 46.355 ;
      RECT  12.195 46.355 23.22 136.125 ;
      RECT  11.78 46.355 12.195 48.67 ;
      RECT  11.78 49.085 12.195 50.88 ;
      RECT  11.78 51.295 12.195 53.61 ;
      RECT  11.78 54.025 12.195 55.82 ;
      RECT  11.78 56.235 12.195 58.55 ;
      RECT  11.78 58.965 12.195 136.125 ;
      RECT  99.28 135.3 99.695 136.125 ;
      RECT  99.695 135.3 120.055 136.125 ;
      RECT  23.635 134.885 96.42 135.3 ;
      RECT  96.835 134.885 99.28 135.3 ;
      RECT  99.695 1.38 107.86 19.81 ;
      RECT  99.695 19.81 107.86 20.225 ;
      RECT  107.86 20.225 108.275 134.885 ;
      RECT  108.275 1.38 120.055 19.81 ;
      RECT  108.275 19.81 120.055 20.225 ;
      RECT  107.86 17.495 108.275 19.81 ;
      RECT  107.86 15.285 108.275 17.08 ;
      RECT  107.86 12.555 108.275 14.87 ;
      RECT  107.86 10.345 108.275 12.14 ;
      RECT  107.86 1.38 108.275 7.2 ;
      RECT  107.86 7.615 108.275 9.93 ;
      RECT  0.14 0.965 0.145 1.35 ;
      RECT  0.14 1.35 0.145 1.38 ;
      RECT  0.145 0.965 0.56 1.35 ;
      RECT  0.56 0.965 17.5 1.35 ;
      RECT  0.56 1.35 17.5 1.38 ;
      RECT  0.14 1.38 0.145 1.765 ;
      RECT  0.14 1.765 0.145 45.94 ;
      RECT  0.145 1.765 0.56 45.94 ;
      RECT  119.635 20.225 120.05 133.51 ;
      RECT  119.635 133.925 120.05 134.885 ;
      RECT  120.05 20.225 120.055 133.51 ;
      RECT  120.05 133.51 120.055 133.925 ;
      RECT  120.05 133.925 120.055 134.885 ;
      RECT  0.56 1.38 6.1075 1.435 ;
      RECT  0.56 1.435 6.1075 1.765 ;
      RECT  6.1075 1.38 6.5225 1.435 ;
      RECT  6.5225 1.38 11.78 1.435 ;
      RECT  6.5225 1.435 11.78 1.765 ;
      RECT  0.56 1.765 6.1075 1.85 ;
      RECT  6.1075 1.85 6.5225 45.94 ;
      RECT  6.5225 1.765 11.78 1.85 ;
      RECT  6.5225 1.85 11.78 45.94 ;
      RECT  108.275 20.225 113.5325 133.425 ;
      RECT  108.275 133.425 113.5325 133.51 ;
      RECT  113.5325 20.225 113.9475 133.425 ;
      RECT  113.9475 133.425 119.635 133.51 ;
      RECT  108.275 133.51 113.5325 133.84 ;
      RECT  108.275 133.84 113.5325 133.925 ;
      RECT  113.5325 133.84 113.9475 133.925 ;
      RECT  113.9475 133.51 119.635 133.84 ;
      RECT  113.9475 133.84 119.635 133.925 ;
      RECT  23.635 130.0175 31.5575 130.4325 ;
      RECT  23.635 130.4325 31.5575 134.885 ;
      RECT  31.5575 130.4325 31.9725 134.885 ;
      RECT  31.9725 130.4325 99.28 134.885 ;
      RECT  31.9725 130.0175 36.2575 130.4325 ;
      RECT  36.6725 130.0175 40.9575 130.4325 ;
      RECT  41.3725 130.0175 45.6575 130.4325 ;
      RECT  46.0725 130.0175 50.3575 130.4325 ;
      RECT  50.7725 130.0175 55.0575 130.4325 ;
      RECT  55.4725 130.0175 59.7575 130.4325 ;
      RECT  60.1725 130.0175 64.4575 130.4325 ;
      RECT  64.8725 130.0175 69.1575 130.4325 ;
      RECT  69.5725 130.0175 73.8575 130.4325 ;
      RECT  74.2725 130.0175 78.5575 130.4325 ;
      RECT  78.9725 130.0175 83.2575 130.4325 ;
      RECT  83.6725 130.0175 99.28 130.4325 ;
      RECT  12.195 40.35 17.5975 40.765 ;
      RECT  18.0125 40.35 23.22 40.765 ;
      RECT  18.0125 40.765 23.22 45.94 ;
      RECT  12.195 1.38 17.2175 2.33 ;
      RECT  12.195 2.33 17.2175 2.745 ;
      RECT  17.2175 1.38 17.5975 2.33 ;
      RECT  17.2175 2.745 17.5975 40.35 ;
      RECT  17.5975 1.38 17.6325 2.33 ;
      RECT  17.6325 1.38 18.0125 2.33 ;
      RECT  17.6325 2.33 18.0125 2.745 ;
      RECT  99.695 20.225 101.8475 25.4 ;
      RECT  99.695 25.4 101.8475 25.815 ;
      RECT  102.2625 25.4 107.86 25.815 ;
      RECT  17.5975 40.765 18.0125 43.34 ;
      RECT  17.5975 43.755 18.0125 45.94 ;
      RECT  23.22 1.38 23.3525 2.33 ;
      RECT  23.22 2.745 23.3525 136.125 ;
      RECT  23.3525 1.38 23.635 2.33 ;
      RECT  23.3525 2.33 23.635 2.745 ;
      RECT  23.3525 2.745 23.635 136.125 ;
      RECT  18.0125 1.38 22.9375 2.33 ;
      RECT  18.0125 2.33 22.9375 2.745 ;
      RECT  18.0125 2.745 22.9375 40.35 ;
      RECT  22.9375 1.38 23.22 2.33 ;
      RECT  22.9375 2.745 23.22 40.35 ;
      RECT  23.635 1.38 28.3725 8.3975 ;
      RECT  23.635 8.3975 28.3725 8.7475 ;
      RECT  28.3725 1.38 31.5575 8.3975 ;
      RECT  31.5575 1.38 31.9725 8.3975 ;
      RECT  84.3425 1.38 99.28 8.3975 ;
      RECT  84.3425 8.3975 99.28 8.7475 ;
      RECT  28.3725 127.81 31.5575 130.0175 ;
      RECT  31.5575 127.81 31.9725 130.0175 ;
      RECT  31.9725 127.81 84.3425 130.0175 ;
      RECT  88.3375 17.0475 99.28 17.3975 ;
      RECT  88.3375 17.3975 95.675 117.3025 ;
      RECT  88.3375 117.3025 95.675 117.7175 ;
      RECT  95.675 17.3975 96.09 117.3025 ;
      RECT  95.675 117.7175 96.09 130.0175 ;
      RECT  96.09 17.3975 99.28 117.3025 ;
      RECT  96.09 117.3025 99.28 117.7175 ;
      RECT  96.09 117.7175 99.28 130.0175 ;
      RECT  101.8475 20.225 102.2625 22.41 ;
      RECT  101.8475 22.825 102.2625 25.4 ;
      RECT  17.5975 2.745 17.6325 22.41 ;
      RECT  17.6325 2.745 18.0125 22.41 ;
      RECT  101.8475 43.755 102.2625 134.885 ;
      RECT  113.9475 20.225 117.495 132.145 ;
      RECT  113.9475 132.145 117.495 132.56 ;
      RECT  113.9475 132.56 117.495 133.425 ;
      RECT  117.495 20.225 117.91 132.145 ;
      RECT  117.495 132.56 117.91 133.425 ;
      RECT  117.91 20.225 119.635 132.145 ;
      RECT  117.91 132.145 119.635 132.56 ;
      RECT  117.91 132.56 119.635 133.425 ;
      RECT  31.9725 1.38 34.3775 2.33 ;
      RECT  31.9725 2.33 34.3775 2.745 ;
      RECT  31.9725 2.745 34.3775 8.3975 ;
      RECT  34.3775 1.38 34.7925 2.33 ;
      RECT  34.3775 2.745 34.7925 8.3975 ;
      RECT  34.7925 1.38 84.3425 2.33 ;
      RECT  34.7925 2.745 84.3425 8.3975 ;
      RECT  84.3425 17.3975 88.3375 120.3475 ;
      RECT  28.3725 17.3975 31.5575 120.3475 ;
      RECT  31.5575 17.3975 31.9725 120.3475 ;
      RECT  31.9725 17.3975 84.3425 120.3475 ;
      RECT  88.3375 117.7175 89.5125 120.3475 ;
      RECT  89.5125 120.3475 95.675 120.6975 ;
      RECT  89.5125 120.6975 95.675 130.0175 ;
      RECT  101.8475 25.815 102.2625 31.38 ;
      RECT  101.8475 31.795 102.2625 34.37 ;
      RECT  99.28 1.38 99.5625 133.52 ;
      RECT  99.28 133.52 99.5625 133.935 ;
      RECT  99.28 133.935 99.5625 134.885 ;
      RECT  99.5625 1.38 99.695 133.52 ;
      RECT  99.5625 133.935 99.695 134.885 ;
      RECT  99.695 25.815 99.9775 133.52 ;
      RECT  99.695 133.935 99.9775 134.885 ;
      RECT  99.9775 25.815 101.8475 133.52 ;
      RECT  99.9775 133.52 101.8475 133.935 ;
      RECT  99.9775 133.935 101.8475 134.885 ;
      RECT  23.635 8.7475 23.77 20.2075 ;
      RECT  23.635 20.2075 23.77 20.6225 ;
      RECT  23.635 20.6225 23.77 130.0175 ;
      RECT  23.77 8.7475 24.185 20.2075 ;
      RECT  23.77 20.6225 24.185 130.0175 ;
      RECT  24.185 20.2075 28.3725 20.6225 ;
      RECT  24.185 20.6225 28.3725 130.0175 ;
      RECT  24.185 8.7475 27.2275 19.42 ;
      RECT  24.185 19.42 27.2275 19.835 ;
      RECT  24.185 19.835 27.2275 20.2075 ;
      RECT  27.2275 8.7475 27.6425 19.42 ;
      RECT  27.2275 19.835 27.6425 20.2075 ;
      RECT  27.6425 8.7475 28.3725 19.42 ;
      RECT  27.6425 19.42 28.3725 19.835 ;
      RECT  27.6425 19.835 28.3725 20.2075 ;
      RECT  0.56 1.85 2.285 2.715 ;
      RECT  0.56 2.715 2.285 3.13 ;
      RECT  0.56 3.13 2.285 45.94 ;
      RECT  2.285 1.85 2.7 2.715 ;
      RECT  2.285 3.13 2.7 45.94 ;
      RECT  2.7 1.85 6.1075 2.715 ;
      RECT  2.7 2.715 6.1075 3.13 ;
      RECT  2.7 3.13 6.1075 45.94 ;
      RECT  34.7925 2.33 45.8175 2.745 ;
      RECT  46.2325 2.33 84.3425 2.745 ;
      RECT  17.5975 31.795 17.6325 34.37 ;
      RECT  17.5975 34.785 17.6325 40.35 ;
      RECT  17.6325 31.795 18.0125 34.37 ;
      RECT  17.6325 34.785 18.0125 40.35 ;
      RECT  89.5125 117.7175 92.2175 118.09 ;
      RECT  89.5125 118.09 92.2175 118.505 ;
      RECT  89.5125 118.505 92.2175 120.3475 ;
      RECT  92.2175 117.7175 92.6325 118.09 ;
      RECT  92.2175 118.505 92.6325 120.3475 ;
      RECT  92.6325 117.7175 95.675 118.09 ;
      RECT  92.6325 118.09 95.675 118.505 ;
      RECT  92.6325 118.505 95.675 120.3475 ;
      RECT  101.8475 34.785 102.2625 40.35 ;
      RECT  101.8475 40.765 102.2625 43.34 ;
      RECT  17.5975 22.825 17.6325 25.4 ;
      RECT  17.5975 25.815 17.6325 31.38 ;
      RECT  17.6325 22.825 18.0125 25.4 ;
      RECT  17.6325 25.815 18.0125 31.38 ;
      RECT  84.3425 8.7475 88.3375 14.4275 ;
      RECT  84.3425 14.7775 88.3375 17.0475 ;
      RECT  88.3375 8.7475 88.37 14.4275 ;
      RECT  88.3375 14.7775 88.37 17.0475 ;
      RECT  88.37 8.7475 99.28 14.4275 ;
      RECT  88.37 14.4275 99.28 14.7775 ;
      RECT  88.37 14.7775 99.28 17.0475 ;
      RECT  28.3725 14.7775 31.5575 17.0475 ;
      RECT  31.5575 14.7775 31.9725 17.0475 ;
      RECT  31.9725 14.7775 84.3425 17.0475 ;
      RECT  12.195 2.745 16.07 38.855 ;
      RECT  12.195 38.855 16.07 39.27 ;
      RECT  12.195 39.27 16.07 40.35 ;
      RECT  16.07 39.27 16.485 40.35 ;
      RECT  16.485 2.745 17.2175 38.855 ;
      RECT  16.485 38.855 17.2175 39.27 ;
      RECT  16.485 39.27 17.2175 40.35 ;
      RECT  12.195 40.765 16.07 44.835 ;
      RECT  12.195 44.835 16.07 45.25 ;
      RECT  12.195 45.25 16.07 45.94 ;
      RECT  16.07 45.25 16.485 45.94 ;
      RECT  16.485 40.765 17.5975 44.835 ;
      RECT  16.485 44.835 17.5975 45.25 ;
      RECT  16.485 45.25 17.5975 45.94 ;
      RECT  84.3425 125.9175 84.3775 130.0175 ;
      RECT  84.3775 125.5675 88.3375 125.9175 ;
      RECT  84.3775 125.9175 88.3375 130.0175 ;
      RECT  28.3725 125.9175 31.5575 127.46 ;
      RECT  31.5575 125.9175 31.9725 127.46 ;
      RECT  31.9725 125.9175 84.3425 127.46 ;
      RECT  102.2625 20.225 103.375 20.915 ;
      RECT  102.2625 20.915 103.375 21.33 ;
      RECT  102.2625 21.33 103.375 25.4 ;
      RECT  103.375 20.225 103.79 20.915 ;
      RECT  103.79 20.225 107.86 20.915 ;
      RECT  103.79 20.915 107.86 21.33 ;
      RECT  103.79 21.33 107.86 25.4 ;
      RECT  23.635 135.3 96.7025 135.99 ;
      RECT  23.635 135.99 96.7025 136.125 ;
      RECT  96.7025 135.3 97.1175 135.99 ;
      RECT  97.1175 135.3 99.28 135.99 ;
      RECT  97.1175 135.99 99.28 136.125 ;
      RECT  102.2625 25.815 103.375 44.835 ;
      RECT  102.2625 44.835 103.375 45.25 ;
      RECT  102.2625 45.25 103.375 134.885 ;
      RECT  103.375 45.25 103.79 134.885 ;
      RECT  103.79 25.815 107.86 44.835 ;
      RECT  103.79 44.835 107.86 45.25 ;
      RECT  103.79 45.25 107.86 134.885 ;
      RECT  99.695 134.885 117.495 135.03 ;
      RECT  99.695 135.03 117.495 135.3 ;
      RECT  117.495 135.03 117.91 135.3 ;
      RECT  117.91 134.885 120.055 135.03 ;
      RECT  117.91 135.03 120.055 135.3 ;
      RECT  108.275 133.925 117.495 134.615 ;
      RECT  108.275 134.615 117.495 134.885 ;
      RECT  117.495 133.925 117.91 134.615 ;
      RECT  117.91 133.925 119.635 134.615 ;
      RECT  117.91 134.615 119.635 134.885 ;
      RECT  23.635 0.14 25.7975 0.275 ;
      RECT  23.635 0.275 25.7975 0.965 ;
      RECT  25.7975 0.275 26.2125 0.965 ;
      RECT  26.2125 0.275 120.055 0.965 ;
      RECT  88.3375 120.6975 88.37 122.9675 ;
      RECT  88.3375 123.3175 88.37 130.0175 ;
      RECT  88.37 120.6975 89.5125 122.9675 ;
      RECT  88.37 122.9675 89.5125 123.3175 ;
      RECT  88.37 123.3175 89.5125 130.0175 ;
      RECT  84.3425 120.6975 84.3775 122.9675 ;
      RECT  84.3425 123.3175 84.3775 125.5675 ;
      RECT  84.3775 120.6975 88.3375 122.9675 ;
      RECT  84.3775 123.3175 88.3375 125.5675 ;
      RECT  28.3725 120.6975 31.5575 122.9675 ;
      RECT  28.3725 123.3175 31.5575 125.5675 ;
      RECT  31.5575 120.6975 31.9725 122.9675 ;
      RECT  31.5575 123.3175 31.9725 125.5675 ;
      RECT  31.9725 120.6975 84.3425 122.9675 ;
      RECT  31.9725 123.3175 84.3425 125.5675 ;
      RECT  49.0925 0.14 120.055 0.275 ;
      RECT  26.2125 0.14 37.2375 0.275 ;
      RECT  37.6525 0.14 48.6775 0.275 ;
      RECT  28.3725 8.7475 31.5575 10.4475 ;
      RECT  28.3725 10.7975 31.5575 14.4275 ;
      RECT  31.5575 8.7475 31.9725 10.4475 ;
      RECT  31.5575 10.7975 31.9725 14.4275 ;
      RECT  31.9725 8.7475 84.3425 10.4475 ;
      RECT  31.9725 10.7975 84.3425 14.4275 ;
      RECT  16.07 30.3 16.485 32.875 ;
      RECT  103.375 42.26 103.79 44.835 ;
      RECT  103.375 21.33 103.79 23.905 ;
      RECT  103.375 24.32 103.79 25.4 ;
      RECT  16.07 27.31 16.485 29.885 ;
      RECT  103.375 39.27 103.79 41.845 ;
      RECT  16.07 33.29 16.485 35.865 ;
      RECT  16.07 36.28 16.485 38.855 ;
      RECT  103.375 25.815 103.79 26.895 ;
      RECT  20.0775 0.275 20.4925 0.965 ;
      RECT  20.4925 0.14 23.22 0.275 ;
      RECT  20.4925 0.275 23.22 0.965 ;
      RECT  103.375 27.31 103.79 29.885 ;
      RECT  0.14 0.14 2.285 0.245 ;
      RECT  0.14 0.245 2.285 0.275 ;
      RECT  2.285 0.14 2.7 0.245 ;
      RECT  2.7 0.14 20.0775 0.245 ;
      RECT  2.7 0.245 20.0775 0.275 ;
      RECT  0.14 0.275 2.285 0.66 ;
      RECT  0.14 0.66 2.285 0.965 ;
      RECT  2.285 0.66 2.7 0.965 ;
      RECT  2.7 0.275 20.0775 0.66 ;
      RECT  2.7 0.66 20.0775 0.965 ;
      RECT  103.375 30.3 103.79 32.875 ;
      RECT  16.07 40.765 16.485 41.845 ;
      RECT  16.07 42.26 16.485 44.835 ;
      RECT  103.375 33.29 103.79 35.865 ;
      RECT  103.375 36.28 103.79 38.855 ;
      RECT  16.07 24.32 16.485 26.895 ;
      RECT  16.07 2.745 16.485 20.915 ;
      RECT  16.07 21.33 16.485 23.905 ;
   LAYER  metal4 ;
      RECT  92.075 0.14 92.775 20.7725 ;
      RECT  92.075 117.1525 92.775 136.125 ;
      RECT  119.0875 20.7725 119.7875 102.3625 ;
      RECT  119.7875 20.7725 120.055 102.3625 ;
      RECT  119.7875 102.3625 120.055 117.1525 ;
      RECT  119.0875 125.325 119.7875 136.125 ;
      RECT  119.7875 117.1525 120.055 125.325 ;
      RECT  119.7875 125.325 120.055 136.125 ;
      RECT  21.165 0.14 21.865 4.565 ;
      RECT  21.865 0.14 92.075 4.565 ;
      RECT  21.865 4.565 92.075 15.145 ;
      RECT  0.14 44.6925 11.355 60.2125 ;
      RECT  0.14 60.2125 11.355 117.1525 ;
      RECT  11.355 20.7725 12.055 44.6925 ;
      RECT  11.355 60.2125 12.055 117.1525 ;
      RECT  92.775 117.2225 96.15 125.325 ;
      RECT  96.15 117.2225 96.85 125.325 ;
      RECT  0.14 120.0725 90.995 136.125 ;
      RECT  90.995 120.0725 91.695 136.125 ;
      RECT  91.695 117.1525 92.075 120.0725 ;
      RECT  91.695 120.0725 92.075 136.125 ;
      RECT  21.865 15.145 90.995 17.6025 ;
      RECT  90.995 15.145 91.695 17.6025 ;
      RECT  91.695 15.145 92.075 17.6025 ;
      RECT  91.695 17.6025 92.075 20.7725 ;
      RECT  91.695 20.7725 92.075 44.6925 ;
      RECT  91.695 44.6925 92.075 60.2125 ;
      RECT  91.695 60.2125 92.075 117.1525 ;
      RECT  105.28 132.7025 105.98 136.125 ;
      RECT  96.85 117.2225 105.28 122.1225 ;
      RECT  105.28 117.2225 105.98 122.1225 ;
      RECT  92.775 125.325 97.995 132.7025 ;
      RECT  92.775 132.7025 97.995 133.18 ;
      RECT  92.775 133.18 97.995 136.125 ;
      RECT  97.995 133.18 98.695 136.125 ;
      RECT  96.85 122.1225 97.995 122.6 ;
      RECT  96.85 122.6 97.995 125.325 ;
      RECT  97.995 122.1225 98.695 122.6 ;
      RECT  27.785 20.7725 28.165 44.6925 ;
      RECT  27.785 44.6925 28.165 60.2125 ;
      RECT  27.785 60.2125 28.165 117.1525 ;
      RECT  0.14 4.565 0.4075 9.95 ;
      RECT  0.14 9.95 0.4075 15.145 ;
      RECT  0.4075 4.565 1.1075 9.95 ;
      RECT  0.14 15.145 0.4075 20.7725 ;
      RECT  0.14 20.7725 0.4075 32.9125 ;
      RECT  0.14 32.9125 0.4075 44.6925 ;
      RECT  0.4075 32.9125 1.1075 44.6925 ;
      RECT  108.0 0.14 108.7 5.9525 ;
      RECT  108.7 0.14 120.055 5.9525 ;
      RECT  108.7 5.9525 120.055 20.7725 ;
      RECT  108.0 21.4725 108.7 102.3625 ;
      RECT  108.7 20.7725 119.0875 21.4725 ;
      RECT  14.075 0.14 14.775 2.5725 ;
      RECT  14.775 0.14 21.165 2.5725 ;
      RECT  14.075 18.0925 14.775 20.7725 ;
      RECT  0.14 117.2225 23.01 120.0725 ;
      RECT  23.01 117.2225 23.71 120.0725 ;
      RECT  23.71 117.2225 28.165 120.0725 ;
      RECT  92.775 20.7725 95.59 102.3625 ;
      RECT  92.775 102.3625 95.59 117.1525 ;
      RECT  92.775 117.1525 95.59 117.185 ;
      RECT  92.775 117.185 95.59 117.2225 ;
      RECT  95.59 117.185 96.15 117.2225 ;
      RECT  92.775 5.9525 95.59 20.74 ;
      RECT  92.775 20.74 95.59 20.7725 ;
      RECT  95.59 5.9525 96.29 20.74 ;
      RECT  1.1075 20.7725 2.47 32.9125 ;
      RECT  3.17 20.7725 11.355 32.9125 ;
      RECT  1.1075 32.9125 2.47 32.945 ;
      RECT  1.1075 32.945 2.47 44.6925 ;
      RECT  2.47 32.945 3.17 44.6925 ;
      RECT  3.17 32.9125 11.355 32.945 ;
      RECT  3.17 32.945 11.355 44.6925 ;
      RECT  1.1075 9.95 2.47 9.9825 ;
      RECT  1.1075 9.9825 2.47 15.145 ;
      RECT  2.47 9.95 3.17 9.9825 ;
      RECT  1.1075 15.145 2.47 18.0925 ;
      RECT  1.1075 18.0925 2.47 20.7725 ;
      RECT  3.17 18.0925 14.075 20.7725 ;
      RECT  0.14 0.14 5.825 2.5725 ;
      RECT  6.525 0.14 14.075 2.5725 ;
      RECT  0.14 2.5725 5.825 4.565 ;
      RECT  6.525 2.5725 14.075 4.565 ;
      RECT  1.1075 4.565 5.825 9.95 ;
      RECT  6.525 4.565 14.075 9.95 ;
      RECT  3.17 9.95 5.825 9.9825 ;
      RECT  6.525 9.95 14.075 9.9825 ;
      RECT  3.17 9.9825 5.825 15.145 ;
      RECT  6.525 9.9825 14.075 15.145 ;
      RECT  3.17 15.145 5.825 15.6225 ;
      RECT  3.17 15.6225 5.825 18.0925 ;
      RECT  5.825 15.6225 6.525 18.0925 ;
      RECT  6.525 15.145 14.075 15.6225 ;
      RECT  6.525 15.6225 14.075 18.0925 ;
      RECT  12.055 20.7725 14.215 44.6275 ;
      RECT  12.055 44.6275 14.215 44.6925 ;
      RECT  14.215 20.7725 14.915 44.6275 ;
      RECT  12.055 44.6925 14.215 60.2125 ;
      RECT  12.055 60.2125 14.215 60.2775 ;
      RECT  12.055 60.2775 14.215 117.1525 ;
      RECT  14.215 60.2775 14.915 117.1525 ;
      RECT  92.775 0.14 105.14 5.8875 ;
      RECT  92.775 5.8875 105.14 5.9525 ;
      RECT  105.14 0.14 105.84 5.8875 ;
      RECT  105.84 0.14 108.0 5.8875 ;
      RECT  105.84 5.8875 108.0 5.9525 ;
      RECT  105.84 20.7725 108.0 21.4725 ;
      RECT  105.14 21.5375 105.84 102.3625 ;
      RECT  105.84 21.4725 108.0 21.5375 ;
      RECT  105.84 21.5375 108.0 102.3625 ;
      RECT  96.29 5.9525 105.14 20.74 ;
      RECT  105.84 5.9525 108.0 20.74 ;
      RECT  105.84 20.74 108.0 20.7725 ;
      RECT  96.85 102.3625 98.085 117.1525 ;
      RECT  96.85 117.1525 98.085 117.2225 ;
      RECT  96.85 20.7725 98.085 21.4725 ;
      RECT  98.785 20.7725 105.14 21.4725 ;
      RECT  96.85 21.4725 98.085 21.5375 ;
      RECT  98.785 21.4725 105.14 21.5375 ;
      RECT  96.85 21.5375 98.085 102.3625 ;
      RECT  98.785 21.5375 105.14 102.3625 ;
      RECT  96.29 20.74 98.085 20.7725 ;
      RECT  98.785 20.74 105.14 20.7725 ;
      RECT  21.165 15.145 21.775 20.74 ;
      RECT  21.775 15.145 21.865 20.74 ;
      RECT  21.775 20.74 21.865 20.7725 ;
      RECT  14.775 18.0925 21.075 20.74 ;
      RECT  14.775 20.74 21.075 20.7725 ;
      RECT  21.075 18.0925 21.165 20.74 ;
      RECT  0.14 117.1525 21.075 117.2225 ;
      RECT  21.775 117.1525 23.01 117.2225 ;
      RECT  14.915 20.7725 21.075 44.6275 ;
      RECT  21.775 20.7725 23.01 44.6275 ;
      RECT  14.915 44.6275 21.075 44.6925 ;
      RECT  21.775 44.6275 23.01 44.6925 ;
      RECT  14.915 44.6925 21.075 60.2125 ;
      RECT  21.775 44.6925 23.01 60.2125 ;
      RECT  14.915 60.2125 21.075 60.2775 ;
      RECT  21.775 60.2125 23.01 60.2775 ;
      RECT  14.915 60.2775 21.075 117.1525 ;
      RECT  21.775 60.2775 23.01 117.1525 ;
      RECT  98.695 125.325 99.6575 132.7025 ;
      RECT  100.3575 125.325 105.28 132.7025 ;
      RECT  98.695 132.7025 99.6575 133.18 ;
      RECT  100.3575 132.7025 105.28 133.18 ;
      RECT  98.695 133.18 99.6575 133.2475 ;
      RECT  98.695 133.2475 99.6575 136.125 ;
      RECT  99.6575 133.2475 100.3575 136.125 ;
      RECT  100.3575 133.18 105.28 133.2475 ;
      RECT  100.3575 133.2475 105.28 136.125 ;
      RECT  98.695 122.1225 99.6575 122.5325 ;
      RECT  98.695 122.5325 99.6575 122.6 ;
      RECT  99.6575 122.1225 100.3575 122.5325 ;
      RECT  100.3575 122.1225 105.28 122.5325 ;
      RECT  100.3575 122.5325 105.28 122.6 ;
      RECT  98.695 122.6 99.6575 125.325 ;
      RECT  100.3575 122.6 105.28 125.325 ;
      RECT  29.325 117.1525 90.535 120.0725 ;
      RECT  29.325 17.6025 90.535 20.7725 ;
      RECT  29.325 20.7725 90.535 44.6925 ;
      RECT  29.325 44.6925 90.535 60.2125 ;
      RECT  29.325 60.2125 90.535 117.1525 ;
      RECT  21.865 17.6025 23.57 20.74 ;
      RECT  21.865 20.74 23.57 20.7725 ;
      RECT  23.57 17.6025 24.27 20.74 ;
      RECT  24.27 17.6025 28.165 20.74 ;
      RECT  24.27 20.74 28.165 20.7725 ;
      RECT  24.27 20.7725 27.085 44.6925 ;
      RECT  24.27 44.6925 27.085 60.2125 ;
      RECT  24.27 60.2125 27.085 117.1525 ;
      RECT  23.71 117.185 24.27 117.2225 ;
      RECT  24.27 117.1525 28.165 117.185 ;
      RECT  24.27 117.185 28.165 117.2225 ;
      RECT  14.775 2.5725 19.5025 4.4975 ;
      RECT  14.775 4.4975 19.5025 4.565 ;
      RECT  19.5025 2.5725 20.2025 4.4975 ;
      RECT  20.2025 2.5725 21.165 4.4975 ;
      RECT  20.2025 4.4975 21.165 4.565 ;
      RECT  14.775 4.565 19.5025 9.95 ;
      RECT  20.2025 4.565 21.165 9.95 ;
      RECT  14.775 9.95 19.5025 15.145 ;
      RECT  20.2025 9.95 21.165 15.145 ;
      RECT  14.775 15.145 19.5025 15.2125 ;
      RECT  14.775 15.2125 19.5025 18.0925 ;
      RECT  19.5025 15.2125 20.2025 18.0925 ;
      RECT  20.2025 15.145 21.165 15.2125 ;
      RECT  20.2025 15.2125 21.165 18.0925 ;
      RECT  117.725 117.2225 119.0875 122.1225 ;
      RECT  117.025 125.2925 117.725 125.325 ;
      RECT  117.725 122.1225 119.0875 125.2925 ;
      RECT  117.725 125.2925 119.0875 125.325 ;
      RECT  108.7 21.4725 117.025 102.33 ;
      RECT  108.7 102.33 117.025 102.3625 ;
      RECT  117.025 21.4725 117.725 102.33 ;
      RECT  117.725 21.4725 119.0875 102.33 ;
      RECT  117.725 102.33 119.0875 102.3625 ;
      RECT  98.785 102.3625 117.025 117.1525 ;
      RECT  117.725 102.3625 119.0875 117.1525 ;
      RECT  98.785 117.1525 117.025 117.2225 ;
      RECT  117.725 117.1525 119.0875 117.2225 ;
      RECT  105.98 125.325 113.53 132.7025 ;
      RECT  114.23 125.325 119.0875 132.7025 ;
      RECT  105.98 132.7025 113.53 135.1725 ;
      RECT  105.98 135.1725 113.53 136.125 ;
      RECT  113.53 135.1725 114.23 136.125 ;
      RECT  114.23 132.7025 119.0875 135.1725 ;
      RECT  114.23 135.1725 119.0875 136.125 ;
      RECT  105.98 117.2225 113.53 119.6525 ;
      RECT  105.98 119.6525 113.53 122.1225 ;
      RECT  113.53 117.2225 114.23 119.6525 ;
      RECT  114.23 117.2225 117.025 119.6525 ;
      RECT  114.23 119.6525 117.025 122.1225 ;
      RECT  105.98 122.1225 113.53 125.2925 ;
      RECT  114.23 122.1225 117.025 125.2925 ;
      RECT  105.98 125.2925 113.53 125.325 ;
      RECT  114.23 125.2925 117.025 125.325 ;
   END
END    freepdk45_sram_1w1r_12x256
END    LIBRARY
