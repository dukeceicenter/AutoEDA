../macros/freepdk45_sram_1w1r_16x72/freepdk45_sram_1w1r_16x72.lef