../macros/freepdk45_sram_1rw0r_20x64/freepdk45_sram_1rw0r_20x64.lef