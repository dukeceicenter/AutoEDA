../macros/freepdk45_sram_1rw0r_64x512/freepdk45_sram_1rw0r_64x512.lef