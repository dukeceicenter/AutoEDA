../macros/freepdk45_sram_1rw0r_22x64/freepdk45_sram_1rw0r_22x64.lef