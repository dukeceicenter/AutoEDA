VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_48x32_32
   CLASS BLOCK ;
   SIZE 112.245 BY 110.59 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.94 1.1075 21.075 1.2425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.8 1.1075 23.935 1.2425 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.66 1.1075 26.795 1.2425 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.52 1.1075 29.655 1.2425 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.38 1.1075 32.515 1.2425 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.24 1.1075 35.375 1.2425 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.1 1.1075 38.235 1.2425 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.96 1.1075 41.095 1.2425 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.82 1.1075 43.955 1.2425 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.68 1.1075 46.815 1.2425 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.54 1.1075 49.675 1.2425 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.4 1.1075 52.535 1.2425 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.26 1.1075 55.395 1.2425 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.12 1.1075 58.255 1.2425 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.98 1.1075 61.115 1.2425 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.84 1.1075 63.975 1.2425 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.7 1.1075 66.835 1.2425 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.56 1.1075 69.695 1.2425 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.42 1.1075 72.555 1.2425 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.28 1.1075 75.415 1.2425 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.14 1.1075 78.275 1.2425 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.0 1.1075 81.135 1.2425 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.86 1.1075 83.995 1.2425 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.72 1.1075 86.855 1.2425 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.58 1.1075 89.715 1.2425 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.44 1.1075 92.575 1.2425 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.3 1.1075 95.435 1.2425 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.16 1.1075 98.295 1.2425 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.02 1.1075 101.155 1.2425 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.88 1.1075 104.015 1.2425 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.74 1.1075 106.875 1.2425 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.6 1.1075 109.735 1.2425 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 45.6975 15.355 45.8325 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 48.4275 15.355 48.5625 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 50.6375 15.355 50.7725 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 53.3675 15.355 53.5025 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 55.5775 15.355 55.7125 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  15.22 58.3075 15.355 58.4425 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.85 19.5675 90.985 19.7025 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.85 16.8375 90.985 16.9725 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.85 14.6275 90.985 14.7625 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.85 11.8975 90.985 12.0325 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.85 9.6875 90.985 9.8225 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.85 6.9575 90.985 7.0925 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1075 0.42 1.2425 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.925 109.3475 106.06 109.4825 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1925 6.3825 1.3275 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.8225 109.2625 99.9575 109.3975 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.1725 102.64 34.3075 102.775 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.3475 102.64 35.4825 102.775 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.5225 102.64 36.6575 102.775 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.6975 102.64 37.8325 102.775 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.8725 102.64 39.0075 102.775 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.0475 102.64 40.1825 102.775 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.2225 102.64 41.3575 102.775 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.3975 102.64 42.5325 102.775 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.5725 102.64 43.7075 102.775 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.7475 102.64 44.8825 102.775 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.9225 102.64 46.0575 102.775 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.0975 102.64 47.2325 102.775 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.2725 102.64 48.4075 102.775 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.4475 102.64 49.5825 102.775 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.6225 102.64 50.7575 102.775 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.7975 102.64 51.9325 102.775 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.9725 102.64 53.1075 102.775 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.1475 102.64 54.2825 102.775 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.3225 102.64 55.4575 102.775 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.4975 102.64 56.6325 102.775 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.6725 102.64 57.8075 102.775 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.8475 102.64 58.9825 102.775 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.0225 102.64 60.1575 102.775 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.1975 102.64 61.3325 102.775 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.3725 102.64 62.5075 102.775 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.5475 102.64 63.6825 102.775 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.7225 102.64 64.8575 102.775 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.8975 102.64 66.0325 102.775 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.0725 102.64 67.2075 102.775 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.2475 102.64 68.3825 102.775 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.4225 102.64 69.5575 102.775 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.5975 102.64 70.7325 102.775 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  29.8425 19.1775 29.9775 19.3125 ;
         LAYER metal3 ;
         RECT  84.8375 31.1375 84.9725 31.2725 ;
         LAYER metal3 ;
         RECT  27.21 19.965 27.345 20.1 ;
         LAYER metal4 ;
         RECT  29.84 20.67 29.98 92.57 ;
         LAYER metal4 ;
         RECT  88.41 98.1 88.55 108.12 ;
         LAYER metal4 ;
         RECT  76.03 20.67 76.17 92.57 ;
         LAYER metal4 ;
         RECT  79.28 20.67 79.42 92.64 ;
         LAYER metal3 ;
         RECT  21.0375 43.0975 21.1725 43.2325 ;
         LAYER metal4 ;
         RECT  105.5175 78.34 105.6575 100.7425 ;
         LAYER metal3 ;
         RECT  30.9875 96.185 73.0475 96.255 ;
         LAYER metal3 ;
         RECT  21.0375 25.1575 21.1725 25.2925 ;
         LAYER metal3 ;
         RECT  2.425 2.4725 2.56 2.6075 ;
         LAYER metal3 ;
         RECT  32.0975 2.4725 32.2325 2.6075 ;
         LAYER metal3 ;
         RECT  66.4175 2.4725 66.5525 2.6075 ;
         LAYER metal3 ;
         RECT  84.8375 25.1575 84.9725 25.2925 ;
         LAYER metal4 ;
         RECT  14.935 44.59 15.075 59.55 ;
         LAYER metal3 ;
         RECT  21.0375 34.1275 21.1725 34.2625 ;
         LAYER metal3 ;
         RECT  89.2975 2.4725 89.4325 2.6075 ;
         LAYER metal4 ;
         RECT  30.92 17.5 31.06 95.49 ;
         LAYER metal3 ;
         RECT  78.665 93.14 78.8 93.275 ;
         LAYER metal4 ;
         RECT  74.95 17.5 75.09 95.49 ;
         LAYER metal3 ;
         RECT  84.8375 43.0975 84.9725 43.2325 ;
         LAYER metal4 ;
         RECT  91.13 5.85 91.27 20.81 ;
         LAYER metal3 ;
         RECT  21.0375 31.1375 21.1725 31.2725 ;
         LAYER metal3 ;
         RECT  30.9875 16.805 71.8725 16.875 ;
         LAYER metal4 ;
         RECT  26.59 20.67 26.73 92.64 ;
         LAYER metal3 ;
         RECT  21.0375 40.1075 21.1725 40.2425 ;
         LAYER metal4 ;
         RECT  17.655 2.47 17.795 17.43 ;
         LAYER metal4 ;
         RECT  0.6875 9.8475 0.8275 32.25 ;
         LAYER metal3 ;
         RECT  54.9775 2.4725 55.1125 2.6075 ;
         LAYER metal3 ;
         RECT  84.8375 34.1275 84.9725 34.2625 ;
         LAYER metal3 ;
         RECT  21.0375 22.1675 21.1725 22.3025 ;
         LAYER metal3 ;
         RECT  30.9875 100.0825 71.4025 100.1525 ;
         LAYER metal3 ;
         RECT  103.785 107.9825 103.92 108.1175 ;
         LAYER metal3 ;
         RECT  20.6575 2.4725 20.7925 2.6075 ;
         LAYER metal3 ;
         RECT  76.0325 93.9275 76.1675 94.0625 ;
         LAYER metal3 ;
         RECT  77.8575 2.4725 77.9925 2.6075 ;
         LAYER metal3 ;
         RECT  43.5375 2.4725 43.6725 2.6075 ;
         LAYER metal3 ;
         RECT  30.9875 11.37 71.4025 11.44 ;
         LAYER metal3 ;
         RECT  100.7375 2.4725 100.8725 2.6075 ;
         LAYER metal3 ;
         RECT  84.8375 22.1675 84.9725 22.3025 ;
         LAYER metal3 ;
         RECT  84.8375 40.1075 84.9725 40.2425 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  27.15 20.6375 27.29 92.6025 ;
         LAYER metal3 ;
         RECT  19.51 26.6525 19.645 26.7875 ;
         LAYER metal3 ;
         RECT  86.365 35.6225 86.5 35.7575 ;
         LAYER metal4 ;
         RECT  2.75 9.88 2.89 32.2825 ;
         LAYER metal4 ;
         RECT  74.49 17.5 74.63 95.49 ;
         LAYER metal3 ;
         RECT  80.7175 0.0025 80.8525 0.1375 ;
         LAYER metal3 ;
         RECT  19.51 44.5925 19.645 44.7275 ;
         LAYER metal4 ;
         RECT  6.105 0.0 6.245 14.96 ;
         LAYER metal3 ;
         RECT  86.365 23.6625 86.5 23.7975 ;
         LAYER metal3 ;
         RECT  86.365 26.6525 86.5 26.7875 ;
         LAYER metal3 ;
         RECT  86.365 29.6425 86.5 29.7775 ;
         LAYER metal4 ;
         RECT  99.96 95.63 100.1 110.59 ;
         LAYER metal3 ;
         RECT  86.365 32.6325 86.5 32.7675 ;
         LAYER metal3 ;
         RECT  69.2775 0.0025 69.4125 0.1375 ;
         LAYER metal3 ;
         RECT  30.9875 98.19 71.4375 98.26 ;
         LAYER metal3 ;
         RECT  57.8375 0.0025 57.9725 0.1375 ;
         LAYER metal3 ;
         RECT  86.365 20.6725 86.5 20.8075 ;
         LAYER metal3 ;
         RECT  19.51 35.6225 19.645 35.7575 ;
         LAYER metal3 ;
         RECT  34.9575 0.0025 35.0925 0.1375 ;
         LAYER metal4 ;
         RECT  24.655 20.6375 24.795 92.64 ;
         LAYER metal3 ;
         RECT  92.1575 0.0025 92.2925 0.1375 ;
         LAYER metal3 ;
         RECT  103.785 110.4525 103.92 110.5875 ;
         LAYER metal3 ;
         RECT  86.365 41.6025 86.5 41.7375 ;
         LAYER metal3 ;
         RECT  23.5175 0.0025 23.6525 0.1375 ;
         LAYER metal3 ;
         RECT  86.365 38.6125 86.5 38.7475 ;
         LAYER metal4 ;
         RECT  31.38 17.5 31.52 95.49 ;
         LAYER metal3 ;
         RECT  19.51 32.6325 19.645 32.7675 ;
         LAYER metal3 ;
         RECT  30.9875 13.42 71.4025 13.49 ;
         LAYER metal3 ;
         RECT  86.365 44.5925 86.5 44.7275 ;
         LAYER metal3 ;
         RECT  19.51 29.6425 19.645 29.7775 ;
         LAYER metal3 ;
         RECT  19.51 20.6725 19.645 20.8075 ;
         LAYER metal3 ;
         RECT  103.5975 0.0025 103.7325 0.1375 ;
         LAYER metal3 ;
         RECT  46.3975 0.0025 46.5325 0.1375 ;
         LAYER metal3 ;
         RECT  2.425 0.0025 2.56 0.1375 ;
         LAYER metal4 ;
         RECT  103.455 78.3075 103.595 100.71 ;
         LAYER metal3 ;
         RECT  19.51 23.6625 19.645 23.7975 ;
         LAYER metal4 ;
         RECT  17.795 44.525 17.935 59.615 ;
         LAYER metal3 ;
         RECT  19.51 41.6025 19.645 41.7375 ;
         LAYER metal3 ;
         RECT  19.51 38.6125 19.645 38.7475 ;
         LAYER metal4 ;
         RECT  81.215 20.6375 81.355 92.64 ;
         LAYER metal4 ;
         RECT  88.27 5.785 88.41 20.875 ;
         LAYER metal4 ;
         RECT  78.72 20.6375 78.86 92.6025 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 112.105 110.45 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 112.105 110.45 ;
   LAYER  metal3 ;
      RECT  20.8 0.14 21.215 0.9675 ;
      RECT  21.215 0.9675 23.66 1.3825 ;
      RECT  24.075 0.9675 26.52 1.3825 ;
      RECT  26.935 0.9675 29.38 1.3825 ;
      RECT  29.795 0.9675 32.24 1.3825 ;
      RECT  32.655 0.9675 35.1 1.3825 ;
      RECT  35.515 0.9675 37.96 1.3825 ;
      RECT  38.375 0.9675 40.82 1.3825 ;
      RECT  41.235 0.9675 43.68 1.3825 ;
      RECT  44.095 0.9675 46.54 1.3825 ;
      RECT  46.955 0.9675 49.4 1.3825 ;
      RECT  49.815 0.9675 52.26 1.3825 ;
      RECT  52.675 0.9675 55.12 1.3825 ;
      RECT  55.535 0.9675 57.98 1.3825 ;
      RECT  58.395 0.9675 60.84 1.3825 ;
      RECT  61.255 0.9675 63.7 1.3825 ;
      RECT  64.115 0.9675 66.56 1.3825 ;
      RECT  66.975 0.9675 69.42 1.3825 ;
      RECT  69.835 0.9675 72.28 1.3825 ;
      RECT  72.695 0.9675 75.14 1.3825 ;
      RECT  75.555 0.9675 78.0 1.3825 ;
      RECT  78.415 0.9675 80.86 1.3825 ;
      RECT  81.275 0.9675 83.72 1.3825 ;
      RECT  84.135 0.9675 86.58 1.3825 ;
      RECT  86.995 0.9675 89.44 1.3825 ;
      RECT  89.855 0.9675 92.3 1.3825 ;
      RECT  92.715 0.9675 95.16 1.3825 ;
      RECT  95.575 0.9675 98.02 1.3825 ;
      RECT  98.435 0.9675 100.88 1.3825 ;
      RECT  101.295 0.9675 103.74 1.3825 ;
      RECT  104.155 0.9675 106.6 1.3825 ;
      RECT  107.015 0.9675 109.46 1.3825 ;
      RECT  109.875 0.9675 112.105 1.3825 ;
      RECT  0.14 45.5575 15.08 45.9725 ;
      RECT  0.14 45.9725 15.08 110.45 ;
      RECT  15.08 1.3825 15.495 45.5575 ;
      RECT  15.495 45.5575 20.8 45.9725 ;
      RECT  15.495 45.9725 20.8 110.45 ;
      RECT  15.08 45.9725 15.495 48.2875 ;
      RECT  15.08 48.7025 15.495 50.4975 ;
      RECT  15.08 50.9125 15.495 53.2275 ;
      RECT  15.08 53.6425 15.495 55.4375 ;
      RECT  15.08 55.8525 15.495 58.1675 ;
      RECT  15.08 58.5825 15.495 110.45 ;
      RECT  90.71 19.8425 91.125 110.45 ;
      RECT  91.125 19.4275 112.105 19.8425 ;
      RECT  90.71 17.1125 91.125 19.4275 ;
      RECT  90.71 14.9025 91.125 16.6975 ;
      RECT  90.71 12.1725 91.125 14.4875 ;
      RECT  90.71 9.9625 91.125 11.7575 ;
      RECT  90.71 1.3825 91.125 6.8175 ;
      RECT  90.71 7.2325 91.125 9.5475 ;
      RECT  0.14 0.9675 0.145 1.3825 ;
      RECT  105.785 19.8425 106.2 109.2075 ;
      RECT  105.785 109.6225 106.2 110.45 ;
      RECT  106.2 19.8425 112.105 109.2075 ;
      RECT  106.2 109.2075 112.105 109.6225 ;
      RECT  106.2 109.6225 112.105 110.45 ;
      RECT  0.14 1.3825 6.1075 1.4675 ;
      RECT  6.1075 1.4675 6.5225 45.5575 ;
      RECT  6.5225 1.3825 15.08 1.4675 ;
      RECT  6.5225 1.4675 15.08 45.5575 ;
      RECT  0.56 0.9675 6.1075 1.0525 ;
      RECT  0.56 1.0525 6.1075 1.3825 ;
      RECT  6.1075 0.9675 6.5225 1.0525 ;
      RECT  6.5225 0.9675 20.8 1.0525 ;
      RECT  6.5225 1.0525 20.8 1.3825 ;
      RECT  91.125 19.8425 99.6825 109.1225 ;
      RECT  91.125 109.1225 99.6825 109.2075 ;
      RECT  99.6825 19.8425 100.0975 109.1225 ;
      RECT  100.0975 109.1225 105.785 109.2075 ;
      RECT  91.125 109.2075 99.6825 109.5375 ;
      RECT  91.125 109.5375 99.6825 109.6225 ;
      RECT  99.6825 109.5375 100.0975 109.6225 ;
      RECT  100.0975 109.2075 105.785 109.5375 ;
      RECT  100.0975 109.5375 105.785 109.6225 ;
      RECT  21.215 102.5 34.0325 102.915 ;
      RECT  21.215 102.915 34.0325 110.45 ;
      RECT  34.0325 102.915 34.4475 110.45 ;
      RECT  34.4475 102.915 90.71 110.45 ;
      RECT  34.4475 102.5 35.2075 102.915 ;
      RECT  35.6225 102.5 36.3825 102.915 ;
      RECT  36.7975 102.5 37.5575 102.915 ;
      RECT  37.9725 102.5 38.7325 102.915 ;
      RECT  39.1475 102.5 39.9075 102.915 ;
      RECT  40.3225 102.5 41.0825 102.915 ;
      RECT  41.4975 102.5 42.2575 102.915 ;
      RECT  42.6725 102.5 43.4325 102.915 ;
      RECT  43.8475 102.5 44.6075 102.915 ;
      RECT  45.0225 102.5 45.7825 102.915 ;
      RECT  46.1975 102.5 46.9575 102.915 ;
      RECT  47.3725 102.5 48.1325 102.915 ;
      RECT  48.5475 102.5 49.3075 102.915 ;
      RECT  49.7225 102.5 50.4825 102.915 ;
      RECT  50.8975 102.5 51.6575 102.915 ;
      RECT  52.0725 102.5 52.8325 102.915 ;
      RECT  53.2475 102.5 54.0075 102.915 ;
      RECT  54.4225 102.5 55.1825 102.915 ;
      RECT  55.5975 102.5 56.3575 102.915 ;
      RECT  56.7725 102.5 57.5325 102.915 ;
      RECT  57.9475 102.5 58.7075 102.915 ;
      RECT  59.1225 102.5 59.8825 102.915 ;
      RECT  60.2975 102.5 61.0575 102.915 ;
      RECT  61.4725 102.5 62.2325 102.915 ;
      RECT  62.6475 102.5 63.4075 102.915 ;
      RECT  63.8225 102.5 64.5825 102.915 ;
      RECT  64.9975 102.5 65.7575 102.915 ;
      RECT  66.1725 102.5 66.9325 102.915 ;
      RECT  67.3475 102.5 68.1075 102.915 ;
      RECT  68.5225 102.5 69.2825 102.915 ;
      RECT  69.6975 102.5 70.4575 102.915 ;
      RECT  70.8725 102.5 90.71 102.915 ;
      RECT  21.215 1.3825 29.7025 19.0375 ;
      RECT  21.215 19.0375 29.7025 19.4275 ;
      RECT  29.7025 1.3825 30.1175 19.0375 ;
      RECT  30.1175 19.0375 90.71 19.4275 ;
      RECT  21.215 19.4275 29.7025 19.4525 ;
      RECT  29.7025 19.4525 30.1175 19.8425 ;
      RECT  30.1175 19.4275 90.71 19.4525 ;
      RECT  30.1175 19.4525 90.71 19.8425 ;
      RECT  34.4475 19.8425 84.6975 30.9975 ;
      RECT  34.4475 30.9975 84.6975 31.4125 ;
      RECT  85.1125 30.9975 90.71 31.4125 ;
      RECT  21.215 19.8425 27.07 20.24 ;
      RECT  27.07 20.24 27.485 102.5 ;
      RECT  27.485 19.8425 34.0325 20.24 ;
      RECT  21.215 19.4525 27.07 19.825 ;
      RECT  21.215 19.825 27.07 19.8425 ;
      RECT  27.07 19.4525 27.485 19.825 ;
      RECT  27.485 19.4525 29.7025 19.825 ;
      RECT  27.485 19.825 29.7025 19.8425 ;
      RECT  20.8 42.9575 20.8975 43.3725 ;
      RECT  20.8 43.3725 20.8975 110.45 ;
      RECT  20.8975 43.3725 21.215 110.45 ;
      RECT  21.215 43.3725 21.3125 102.5 ;
      RECT  21.3125 20.24 27.07 42.9575 ;
      RECT  21.3125 42.9575 27.07 43.3725 ;
      RECT  21.3125 43.3725 27.07 102.5 ;
      RECT  34.0325 19.8425 34.4475 96.045 ;
      RECT  34.4475 31.4125 73.1875 96.045 ;
      RECT  73.1875 96.045 84.6975 96.395 ;
      RECT  73.1875 96.395 84.6975 102.5 ;
      RECT  27.485 20.24 30.8475 96.045 ;
      RECT  27.485 96.045 30.8475 96.395 ;
      RECT  27.485 96.395 30.8475 102.5 ;
      RECT  30.8475 20.24 34.0325 96.045 ;
      RECT  0.14 1.4675 2.285 2.3325 ;
      RECT  0.14 2.3325 2.285 2.7475 ;
      RECT  0.14 2.7475 2.285 45.5575 ;
      RECT  2.285 1.4675 2.7 2.3325 ;
      RECT  2.285 2.7475 2.7 45.5575 ;
      RECT  2.7 1.4675 6.1075 2.3325 ;
      RECT  2.7 2.3325 6.1075 2.7475 ;
      RECT  2.7 2.7475 6.1075 45.5575 ;
      RECT  30.1175 1.3825 31.9575 2.3325 ;
      RECT  30.1175 2.3325 31.9575 2.7475 ;
      RECT  31.9575 1.3825 32.3725 2.3325 ;
      RECT  32.3725 1.3825 90.71 2.3325 ;
      RECT  84.6975 25.4325 85.1125 30.9975 ;
      RECT  89.5725 2.3325 90.71 2.7475 ;
      RECT  73.1875 31.4125 78.525 93.0 ;
      RECT  73.1875 93.0 78.525 93.415 ;
      RECT  78.525 31.4125 78.94 93.0 ;
      RECT  78.525 93.415 78.94 96.045 ;
      RECT  78.94 31.4125 84.6975 93.0 ;
      RECT  78.94 93.0 84.6975 93.415 ;
      RECT  78.94 93.415 84.6975 96.045 ;
      RECT  84.6975 43.3725 85.1125 102.5 ;
      RECT  20.8975 25.4325 21.215 30.9975 ;
      RECT  20.8975 31.4125 21.215 33.9875 ;
      RECT  21.215 25.4325 21.3125 30.9975 ;
      RECT  21.215 31.4125 21.3125 33.9875 ;
      RECT  30.1175 2.7475 30.8475 16.665 ;
      RECT  30.1175 16.665 30.8475 17.015 ;
      RECT  30.1175 17.015 30.8475 19.0375 ;
      RECT  30.8475 17.015 31.9575 19.0375 ;
      RECT  31.9575 17.015 32.3725 19.0375 ;
      RECT  32.3725 17.015 72.0125 19.0375 ;
      RECT  72.0125 2.7475 90.71 16.665 ;
      RECT  72.0125 16.665 90.71 17.015 ;
      RECT  72.0125 17.015 90.71 19.0375 ;
      RECT  20.8975 34.4025 21.215 39.9675 ;
      RECT  20.8975 40.3825 21.215 42.9575 ;
      RECT  21.215 34.4025 21.3125 39.9675 ;
      RECT  21.215 40.3825 21.3125 42.9575 ;
      RECT  55.2525 2.3325 66.2775 2.7475 ;
      RECT  84.6975 31.4125 85.1125 33.9875 ;
      RECT  20.8975 22.4425 21.215 25.0175 ;
      RECT  21.215 20.24 21.3125 22.0275 ;
      RECT  21.215 22.4425 21.3125 25.0175 ;
      RECT  34.0325 100.2925 34.4475 102.5 ;
      RECT  34.4475 100.2925 71.5425 102.5 ;
      RECT  71.5425 99.9425 73.1875 100.2925 ;
      RECT  71.5425 100.2925 73.1875 102.5 ;
      RECT  30.8475 100.2925 34.0325 102.5 ;
      RECT  100.0975 19.8425 103.645 107.8425 ;
      RECT  100.0975 107.8425 103.645 108.2575 ;
      RECT  100.0975 108.2575 103.645 109.1225 ;
      RECT  103.645 19.8425 104.06 107.8425 ;
      RECT  103.645 108.2575 104.06 109.1225 ;
      RECT  104.06 19.8425 105.785 107.8425 ;
      RECT  104.06 107.8425 105.785 108.2575 ;
      RECT  104.06 108.2575 105.785 109.1225 ;
      RECT  15.495 1.3825 20.5175 2.3325 ;
      RECT  15.495 2.3325 20.5175 2.7475 ;
      RECT  20.5175 1.3825 20.8 2.3325 ;
      RECT  20.5175 2.7475 20.8 45.5575 ;
      RECT  20.8 1.3825 20.8975 2.3325 ;
      RECT  20.8 2.7475 20.8975 42.9575 ;
      RECT  20.8975 1.3825 20.9325 2.3325 ;
      RECT  20.8975 2.7475 20.9325 22.0275 ;
      RECT  20.9325 1.3825 21.215 2.3325 ;
      RECT  20.9325 2.3325 21.215 2.7475 ;
      RECT  20.9325 2.7475 21.215 22.0275 ;
      RECT  73.1875 93.415 75.8925 93.7875 ;
      RECT  73.1875 93.7875 75.8925 94.2025 ;
      RECT  73.1875 94.2025 75.8925 96.045 ;
      RECT  75.8925 93.415 76.3075 93.7875 ;
      RECT  75.8925 94.2025 76.3075 96.045 ;
      RECT  76.3075 93.415 78.525 93.7875 ;
      RECT  76.3075 93.7875 78.525 94.2025 ;
      RECT  76.3075 94.2025 78.525 96.045 ;
      RECT  66.6925 2.3325 77.7175 2.7475 ;
      RECT  78.1325 2.3325 89.1575 2.7475 ;
      RECT  32.3725 2.3325 43.3975 2.7475 ;
      RECT  43.8125 2.3325 54.8375 2.7475 ;
      RECT  30.8475 2.7475 31.9575 11.23 ;
      RECT  31.9575 2.7475 32.3725 11.23 ;
      RECT  32.3725 2.7475 71.5425 11.23 ;
      RECT  71.5425 2.7475 72.0125 11.23 ;
      RECT  71.5425 11.23 72.0125 11.58 ;
      RECT  71.5425 11.58 72.0125 16.665 ;
      RECT  91.125 1.3825 100.5975 2.3325 ;
      RECT  91.125 2.3325 100.5975 2.7475 ;
      RECT  91.125 2.7475 100.5975 19.4275 ;
      RECT  100.5975 1.3825 101.0125 2.3325 ;
      RECT  100.5975 2.7475 101.0125 19.4275 ;
      RECT  101.0125 1.3825 112.105 2.3325 ;
      RECT  101.0125 2.3325 112.105 2.7475 ;
      RECT  101.0125 2.7475 112.105 19.4275 ;
      RECT  84.6975 19.8425 85.1125 22.0275 ;
      RECT  84.6975 22.4425 85.1125 25.0175 ;
      RECT  84.6975 34.4025 85.1125 39.9675 ;
      RECT  84.6975 40.3825 85.1125 42.9575 ;
      RECT  15.495 2.7475 19.37 26.5125 ;
      RECT  15.495 26.5125 19.37 26.9275 ;
      RECT  15.495 26.9275 19.37 45.5575 ;
      RECT  19.785 2.7475 20.5175 26.5125 ;
      RECT  19.785 26.5125 20.5175 26.9275 ;
      RECT  19.785 26.9275 20.5175 45.5575 ;
      RECT  85.1125 31.4125 86.225 35.4825 ;
      RECT  85.1125 35.4825 86.225 35.8975 ;
      RECT  85.1125 35.8975 86.225 102.5 ;
      RECT  86.64 31.4125 90.71 35.4825 ;
      RECT  86.64 35.4825 90.71 35.8975 ;
      RECT  86.64 35.8975 90.71 102.5 ;
      RECT  21.215 0.2775 80.5775 0.9675 ;
      RECT  80.5775 0.2775 80.9925 0.9675 ;
      RECT  80.9925 0.2775 112.105 0.9675 ;
      RECT  19.37 44.8675 19.785 45.5575 ;
      RECT  85.1125 19.8425 86.225 23.5225 ;
      RECT  85.1125 23.5225 86.225 23.9375 ;
      RECT  85.1125 23.9375 86.225 30.9975 ;
      RECT  86.64 19.8425 90.71 23.5225 ;
      RECT  86.64 23.5225 90.71 23.9375 ;
      RECT  86.64 23.9375 90.71 30.9975 ;
      RECT  86.225 23.9375 86.64 26.5125 ;
      RECT  86.225 26.9275 86.64 29.5025 ;
      RECT  86.225 29.9175 86.64 30.9975 ;
      RECT  86.225 31.4125 86.64 32.4925 ;
      RECT  86.225 32.9075 86.64 35.4825 ;
      RECT  69.5525 0.14 80.5775 0.2775 ;
      RECT  34.0325 96.395 34.4475 98.05 ;
      RECT  34.0325 98.4 34.4475 99.9425 ;
      RECT  34.4475 96.395 71.5425 98.05 ;
      RECT  34.4475 98.4 71.5425 99.9425 ;
      RECT  71.5425 96.395 71.5775 98.05 ;
      RECT  71.5425 98.4 71.5775 99.9425 ;
      RECT  71.5775 96.395 73.1875 98.05 ;
      RECT  71.5775 98.05 73.1875 98.4 ;
      RECT  71.5775 98.4 73.1875 99.9425 ;
      RECT  30.8475 96.395 34.0325 98.05 ;
      RECT  30.8475 98.4 34.0325 99.9425 ;
      RECT  58.1125 0.14 69.1375 0.2775 ;
      RECT  86.225 19.8425 86.64 20.5325 ;
      RECT  86.225 20.9475 86.64 23.5225 ;
      RECT  80.9925 0.14 92.0175 0.2775 ;
      RECT  91.125 109.6225 103.645 110.3125 ;
      RECT  91.125 110.3125 103.645 110.45 ;
      RECT  103.645 109.6225 104.06 110.3125 ;
      RECT  104.06 109.6225 105.785 110.3125 ;
      RECT  104.06 110.3125 105.785 110.45 ;
      RECT  21.215 0.14 23.3775 0.2775 ;
      RECT  23.7925 0.14 34.8175 0.2775 ;
      RECT  86.225 35.8975 86.64 38.4725 ;
      RECT  86.225 38.8875 86.64 41.4625 ;
      RECT  19.37 32.9075 19.785 35.4825 ;
      RECT  30.8475 11.58 31.9575 13.28 ;
      RECT  30.8475 13.63 31.9575 16.665 ;
      RECT  31.9575 11.58 32.3725 13.28 ;
      RECT  31.9575 13.63 32.3725 16.665 ;
      RECT  32.3725 11.58 71.5425 13.28 ;
      RECT  32.3725 13.63 71.5425 16.665 ;
      RECT  86.225 41.8775 86.64 44.4525 ;
      RECT  86.225 44.8675 86.64 102.5 ;
      RECT  19.37 26.9275 19.785 29.5025 ;
      RECT  19.37 29.9175 19.785 32.4925 ;
      RECT  19.37 2.7475 19.785 20.5325 ;
      RECT  92.4325 0.14 103.4575 0.2775 ;
      RECT  103.8725 0.14 112.105 0.2775 ;
      RECT  35.2325 0.14 46.2575 0.2775 ;
      RECT  46.6725 0.14 57.6975 0.2775 ;
      RECT  0.14 0.14 2.285 0.2775 ;
      RECT  0.14 0.2775 2.285 0.9675 ;
      RECT  2.285 0.2775 2.7 0.9675 ;
      RECT  2.7 0.14 20.8 0.2775 ;
      RECT  2.7 0.2775 20.8 0.9675 ;
      RECT  19.37 20.9475 19.785 23.5225 ;
      RECT  19.37 23.9375 19.785 26.5125 ;
      RECT  19.37 41.8775 19.785 44.4525 ;
      RECT  19.37 35.8975 19.785 38.4725 ;
      RECT  19.37 38.8875 19.785 41.4625 ;
   LAYER  metal4 ;
      RECT  29.56 0.14 30.26 20.39 ;
      RECT  29.56 92.85 30.26 110.45 ;
      RECT  30.26 97.82 88.13 108.4 ;
      RECT  30.26 108.4 88.13 110.45 ;
      RECT  88.13 92.85 88.83 97.82 ;
      RECT  88.13 108.4 88.83 110.45 ;
      RECT  79.0 92.92 79.7 97.82 ;
      RECT  79.7 92.92 88.13 97.82 ;
      RECT  105.9375 92.85 112.105 97.82 ;
      RECT  105.2375 101.0225 105.9375 108.4 ;
      RECT  105.9375 97.82 112.105 101.0225 ;
      RECT  105.9375 101.0225 112.105 108.4 ;
      RECT  105.2375 20.39 105.9375 78.06 ;
      RECT  105.9375 20.39 112.105 78.06 ;
      RECT  105.9375 78.06 112.105 92.85 ;
      RECT  0.14 44.31 14.655 59.83 ;
      RECT  0.14 59.83 14.655 92.85 ;
      RECT  14.655 20.39 15.355 44.31 ;
      RECT  14.655 59.83 15.355 92.85 ;
      RECT  30.26 0.14 30.64 17.22 ;
      RECT  30.26 17.22 30.64 20.39 ;
      RECT  30.64 0.14 31.34 17.22 ;
      RECT  30.26 20.39 30.64 92.85 ;
      RECT  30.26 92.85 30.64 92.92 ;
      RECT  30.26 92.92 30.64 95.77 ;
      RECT  30.26 95.77 30.64 97.82 ;
      RECT  30.64 95.77 31.34 97.82 ;
      RECT  31.34 95.77 79.0 97.82 ;
      RECT  75.37 20.39 75.75 92.85 ;
      RECT  75.37 92.92 79.0 95.77 ;
      RECT  90.85 21.09 91.55 78.06 ;
      RECT  91.55 20.39 105.2375 21.09 ;
      RECT  90.85 0.14 91.55 5.57 ;
      RECT  91.55 0.14 112.105 5.57 ;
      RECT  91.55 5.57 112.105 17.22 ;
      RECT  91.55 17.22 112.105 20.39 ;
      RECT  0.14 92.92 26.31 110.45 ;
      RECT  26.31 92.92 27.01 110.45 ;
      RECT  27.01 92.92 29.56 110.45 ;
      RECT  17.375 0.14 18.075 2.19 ;
      RECT  17.375 17.71 18.075 20.39 ;
      RECT  18.075 0.14 29.56 2.19 ;
      RECT  18.075 2.19 29.56 17.71 ;
      RECT  0.14 20.39 0.4075 32.53 ;
      RECT  0.14 32.53 0.4075 44.31 ;
      RECT  0.4075 32.53 1.1075 44.31 ;
      RECT  0.14 2.19 0.4075 9.5675 ;
      RECT  0.14 9.5675 0.4075 17.71 ;
      RECT  0.4075 2.19 1.1075 9.5675 ;
      RECT  0.14 17.71 0.4075 20.39 ;
      RECT  27.01 92.8825 27.57 92.92 ;
      RECT  27.57 92.85 29.56 92.8825 ;
      RECT  27.57 92.8825 29.56 92.92 ;
      RECT  27.57 20.39 29.56 44.31 ;
      RECT  27.57 44.31 29.56 59.83 ;
      RECT  27.57 59.83 29.56 92.85 ;
      RECT  18.075 17.71 26.87 20.3575 ;
      RECT  26.87 17.71 27.57 20.3575 ;
      RECT  27.57 17.71 29.56 20.3575 ;
      RECT  27.57 20.3575 29.56 20.39 ;
      RECT  1.1075 20.39 2.47 32.53 ;
      RECT  3.17 20.39 14.655 32.53 ;
      RECT  1.1075 32.53 2.47 32.5625 ;
      RECT  1.1075 32.5625 2.47 44.31 ;
      RECT  2.47 32.5625 3.17 44.31 ;
      RECT  3.17 32.53 14.655 32.5625 ;
      RECT  3.17 32.5625 14.655 44.31 ;
      RECT  1.1075 9.5675 2.47 9.6 ;
      RECT  1.1075 9.6 2.47 17.71 ;
      RECT  2.47 9.5675 3.17 9.6 ;
      RECT  1.1075 17.71 2.47 20.39 ;
      RECT  3.17 17.71 17.375 20.39 ;
      RECT  0.14 0.14 5.825 2.19 ;
      RECT  6.525 0.14 17.375 2.19 ;
      RECT  1.1075 2.19 5.825 9.5675 ;
      RECT  6.525 2.19 17.375 9.5675 ;
      RECT  3.17 9.5675 5.825 9.6 ;
      RECT  6.525 9.5675 17.375 9.6 ;
      RECT  3.17 9.6 5.825 15.24 ;
      RECT  3.17 15.24 5.825 17.71 ;
      RECT  5.825 15.24 6.525 17.71 ;
      RECT  6.525 9.6 17.375 15.24 ;
      RECT  6.525 15.24 17.375 17.71 ;
      RECT  88.83 108.4 99.68 110.45 ;
      RECT  100.38 108.4 112.105 110.45 ;
      RECT  88.83 92.85 99.68 95.35 ;
      RECT  88.83 95.35 99.68 97.82 ;
      RECT  99.68 92.85 100.38 95.35 ;
      RECT  88.83 97.82 99.68 101.0225 ;
      RECT  88.83 101.0225 99.68 108.4 ;
      RECT  100.38 101.0225 105.2375 108.4 ;
      RECT  0.14 92.85 24.375 92.92 ;
      RECT  25.075 92.85 26.31 92.92 ;
      RECT  25.075 20.39 26.31 44.31 ;
      RECT  25.075 44.31 26.31 59.83 ;
      RECT  25.075 59.83 26.31 92.85 ;
      RECT  18.075 20.3575 24.375 20.39 ;
      RECT  25.075 20.3575 26.87 20.39 ;
      RECT  31.8 17.22 74.21 20.39 ;
      RECT  31.8 20.39 74.21 92.85 ;
      RECT  31.8 92.85 74.21 92.92 ;
      RECT  31.8 92.92 74.21 95.77 ;
      RECT  103.875 78.06 105.2375 92.85 ;
      RECT  91.55 21.09 103.175 78.0275 ;
      RECT  91.55 78.0275 103.175 78.06 ;
      RECT  103.175 21.09 103.875 78.0275 ;
      RECT  103.875 21.09 105.2375 78.0275 ;
      RECT  103.875 78.0275 105.2375 78.06 ;
      RECT  100.38 92.85 103.175 95.35 ;
      RECT  103.875 92.85 105.2375 95.35 ;
      RECT  100.38 95.35 103.175 97.82 ;
      RECT  103.875 95.35 105.2375 97.82 ;
      RECT  100.38 97.82 103.175 100.99 ;
      RECT  100.38 100.99 103.175 101.0225 ;
      RECT  103.175 100.99 103.875 101.0225 ;
      RECT  103.875 97.82 105.2375 100.99 ;
      RECT  103.875 100.99 105.2375 101.0225 ;
      RECT  15.355 20.39 17.515 44.245 ;
      RECT  15.355 44.245 17.515 44.31 ;
      RECT  17.515 20.39 18.215 44.245 ;
      RECT  18.215 20.39 24.375 44.245 ;
      RECT  18.215 44.245 24.375 44.31 ;
      RECT  15.355 44.31 17.515 59.83 ;
      RECT  18.215 44.31 24.375 59.83 ;
      RECT  15.355 59.83 17.515 59.895 ;
      RECT  15.355 59.895 17.515 92.85 ;
      RECT  17.515 59.895 18.215 92.85 ;
      RECT  18.215 59.83 24.375 59.895 ;
      RECT  18.215 59.895 24.375 92.85 ;
      RECT  79.7 92.85 80.935 92.92 ;
      RECT  81.635 92.85 88.13 92.92 ;
      RECT  79.7 20.39 80.935 21.09 ;
      RECT  79.7 21.09 80.935 78.06 ;
      RECT  75.37 17.22 80.935 20.3575 ;
      RECT  80.935 17.22 81.635 20.3575 ;
      RECT  79.7 78.06 80.935 92.85 ;
      RECT  81.635 78.06 103.175 92.85 ;
      RECT  31.34 0.14 87.99 5.505 ;
      RECT  31.34 5.505 87.99 5.57 ;
      RECT  87.99 0.14 88.69 5.505 ;
      RECT  88.69 0.14 90.85 5.505 ;
      RECT  88.69 5.505 90.85 5.57 ;
      RECT  31.34 5.57 87.99 17.22 ;
      RECT  88.69 5.57 90.85 17.22 ;
      RECT  81.635 20.39 87.99 21.09 ;
      RECT  88.69 20.39 90.85 21.09 ;
      RECT  81.635 21.09 87.99 21.155 ;
      RECT  81.635 21.155 87.99 78.06 ;
      RECT  87.99 21.155 88.69 78.06 ;
      RECT  88.69 21.09 90.85 21.155 ;
      RECT  88.69 21.155 90.85 78.06 ;
      RECT  81.635 17.22 87.99 20.3575 ;
      RECT  88.69 17.22 90.85 20.3575 ;
      RECT  81.635 20.3575 87.99 20.39 ;
      RECT  88.69 20.3575 90.85 20.39 ;
      RECT  76.45 20.39 78.44 92.85 ;
      RECT  75.37 92.85 78.44 92.8825 ;
      RECT  75.37 92.8825 78.44 92.92 ;
      RECT  78.44 92.8825 79.0 92.92 ;
      RECT  75.37 20.3575 78.44 20.39 ;
      RECT  79.14 20.3575 80.935 20.39 ;
   END
END    freepdk45_sram_1w1r_48x32_32
END    LIBRARY
