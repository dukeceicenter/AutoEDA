../macros/freepdk45_sram_1w1r_32x240/freepdk45_sram_1w1r_32x240.lef