../macros/freepdk45_sram_1rw0r_64x160_20/freepdk45_sram_1rw0r_64x160_20.lef