../macros/freepdk45_sram_1w1r_32x120/freepdk45_sram_1w1r_32x120.lef