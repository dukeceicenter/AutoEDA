../macros/freepdk45_sram_1w1r_38x96_32/freepdk45_sram_1w1r_38x96_32.lef