VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_16x120
   CLASS BLOCK ;
   SIZE 383.725 BY 73.3525 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.74 1.105 40.875 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.6 1.105 43.735 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.46 1.105 46.595 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.32 1.105 49.455 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.18 1.105 52.315 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.04 1.105 55.175 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.9 1.105 58.035 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.76 1.105 60.895 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.62 1.105 63.755 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.48 1.105 66.615 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.34 1.105 69.475 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.2 1.105 72.335 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.06 1.105 75.195 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.92 1.105 78.055 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.78 1.105 80.915 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.64 1.105 83.775 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.5 1.105 86.635 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.36 1.105 89.495 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.22 1.105 92.355 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.08 1.105 95.215 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.94 1.105 98.075 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.8 1.105 100.935 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.66 1.105 103.795 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.52 1.105 106.655 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.38 1.105 109.515 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.24 1.105 112.375 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.1 1.105 115.235 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.96 1.105 118.095 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.82 1.105 120.955 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.68 1.105 123.815 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.54 1.105 126.675 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.4 1.105 129.535 1.24 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.26 1.105 132.395 1.24 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.12 1.105 135.255 1.24 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.98 1.105 138.115 1.24 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.84 1.105 140.975 1.24 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.7 1.105 143.835 1.24 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.56 1.105 146.695 1.24 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.42 1.105 149.555 1.24 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.28 1.105 152.415 1.24 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.14 1.105 155.275 1.24 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.0 1.105 158.135 1.24 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.86 1.105 160.995 1.24 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.72 1.105 163.855 1.24 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.58 1.105 166.715 1.24 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.44 1.105 169.575 1.24 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.3 1.105 172.435 1.24 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.16 1.105 175.295 1.24 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.02 1.105 178.155 1.24 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.88 1.105 181.015 1.24 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.74 1.105 183.875 1.24 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.6 1.105 186.735 1.24 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.46 1.105 189.595 1.24 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.32 1.105 192.455 1.24 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.18 1.105 195.315 1.24 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.04 1.105 198.175 1.24 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.9 1.105 201.035 1.24 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.76 1.105 203.895 1.24 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.62 1.105 206.755 1.24 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.48 1.105 209.615 1.24 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.34 1.105 212.475 1.24 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.2 1.105 215.335 1.24 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.06 1.105 218.195 1.24 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.92 1.105 221.055 1.24 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.78 1.105 223.915 1.24 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.64 1.105 226.775 1.24 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.5 1.105 229.635 1.24 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.36 1.105 232.495 1.24 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.22 1.105 235.355 1.24 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.08 1.105 238.215 1.24 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.94 1.105 241.075 1.24 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.8 1.105 243.935 1.24 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.66 1.105 246.795 1.24 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.52 1.105 249.655 1.24 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.38 1.105 252.515 1.24 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.24 1.105 255.375 1.24 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.1 1.105 258.235 1.24 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.96 1.105 261.095 1.24 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.82 1.105 263.955 1.24 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.68 1.105 266.815 1.24 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.54 1.105 269.675 1.24 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.4 1.105 272.535 1.24 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.26 1.105 275.395 1.24 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.12 1.105 278.255 1.24 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.98 1.105 281.115 1.24 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.84 1.105 283.975 1.24 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.7 1.105 286.835 1.24 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.56 1.105 289.695 1.24 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.42 1.105 292.555 1.24 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.28 1.105 295.415 1.24 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.14 1.105 298.275 1.24 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.0 1.105 301.135 1.24 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.86 1.105 303.995 1.24 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.72 1.105 306.855 1.24 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.58 1.105 309.715 1.24 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.44 1.105 312.575 1.24 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.3 1.105 315.435 1.24 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.16 1.105 318.295 1.24 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.02 1.105 321.155 1.24 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.88 1.105 324.015 1.24 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.74 1.105 326.875 1.24 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.6 1.105 329.735 1.24 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.46 1.105 332.595 1.24 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.32 1.105 335.455 1.24 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.18 1.105 338.315 1.24 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.04 1.105 341.175 1.24 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.9 1.105 344.035 1.24 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.76 1.105 346.895 1.24 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.62 1.105 349.755 1.24 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.48 1.105 352.615 1.24 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.34 1.105 355.475 1.24 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.2 1.105 358.335 1.24 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.06 1.105 361.195 1.24 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.92 1.105 364.055 1.24 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.78 1.105 366.915 1.24 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.64 1.105 369.775 1.24 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.5 1.105 372.635 1.24 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.36 1.105 375.495 1.24 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.22 1.105 378.355 1.24 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.08 1.105 381.215 1.24 ;
      END
   END din0[119]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.02 47.33 35.155 47.465 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.02 50.06 35.155 50.195 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.02 52.27 35.155 52.405 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.02 55.0 35.155 55.135 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.38 30.17 219.515 30.305 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.38 27.44 219.515 27.575 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.38 25.23 219.515 25.365 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.38 22.5 219.515 22.635 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 11.71 0.42 11.845 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.255 72.11 254.39 72.245 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 11.795 6.3825 11.93 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.1525 72.025 248.2875 72.16 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.6375 65.4025 56.7725 65.5375 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.8125 65.4025 57.9475 65.5375 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.9875 65.4025 59.1225 65.5375 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.1625 65.4025 60.2975 65.5375 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.3375 65.4025 61.4725 65.5375 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.5125 65.4025 62.6475 65.5375 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.6875 65.4025 63.8225 65.5375 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.8625 65.4025 64.9975 65.5375 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.0375 65.4025 66.1725 65.5375 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.2125 65.4025 67.3475 65.5375 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.3875 65.4025 68.5225 65.5375 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.5625 65.4025 69.6975 65.5375 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.7375 65.4025 70.8725 65.5375 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.9125 65.4025 72.0475 65.5375 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.0875 65.4025 73.2225 65.5375 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.2625 65.4025 74.3975 65.5375 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.4375 65.4025 75.5725 65.5375 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.6125 65.4025 76.7475 65.5375 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.7875 65.4025 77.9225 65.5375 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.9625 65.4025 79.0975 65.5375 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.1375 65.4025 80.2725 65.5375 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.3125 65.4025 81.4475 65.5375 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.4875 65.4025 82.6225 65.5375 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.6625 65.4025 83.7975 65.5375 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.8375 65.4025 84.9725 65.5375 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.0125 65.4025 86.1475 65.5375 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.1875 65.4025 87.3225 65.5375 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.3625 65.4025 88.4975 65.5375 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.5375 65.4025 89.6725 65.5375 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.7125 65.4025 90.8475 65.5375 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.8875 65.4025 92.0225 65.5375 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.0625 65.4025 93.1975 65.5375 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.2375 65.4025 94.3725 65.5375 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.4125 65.4025 95.5475 65.5375 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.5875 65.4025 96.7225 65.5375 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.7625 65.4025 97.8975 65.5375 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.9375 65.4025 99.0725 65.5375 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.1125 65.4025 100.2475 65.5375 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.2875 65.4025 101.4225 65.5375 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.4625 65.4025 102.5975 65.5375 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.6375 65.4025 103.7725 65.5375 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.8125 65.4025 104.9475 65.5375 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.9875 65.4025 106.1225 65.5375 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.1625 65.4025 107.2975 65.5375 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.3375 65.4025 108.4725 65.5375 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.5125 65.4025 109.6475 65.5375 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.6875 65.4025 110.8225 65.5375 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.8625 65.4025 111.9975 65.5375 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.0375 65.4025 113.1725 65.5375 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.2125 65.4025 114.3475 65.5375 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.3875 65.4025 115.5225 65.5375 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.5625 65.4025 116.6975 65.5375 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.7375 65.4025 117.8725 65.5375 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.9125 65.4025 119.0475 65.5375 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.0875 65.4025 120.2225 65.5375 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.2625 65.4025 121.3975 65.5375 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.4375 65.4025 122.5725 65.5375 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.6125 65.4025 123.7475 65.5375 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.7875 65.4025 124.9225 65.5375 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.9625 65.4025 126.0975 65.5375 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.1375 65.4025 127.2725 65.5375 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.3125 65.4025 128.4475 65.5375 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.4875 65.4025 129.6225 65.5375 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.6625 65.4025 130.7975 65.5375 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.8375 65.4025 131.9725 65.5375 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.0125 65.4025 133.1475 65.5375 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.1875 65.4025 134.3225 65.5375 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.3625 65.4025 135.4975 65.5375 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.5375 65.4025 136.6725 65.5375 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.7125 65.4025 137.8475 65.5375 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.8875 65.4025 139.0225 65.5375 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.0625 65.4025 140.1975 65.5375 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.2375 65.4025 141.3725 65.5375 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.4125 65.4025 142.5475 65.5375 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.5875 65.4025 143.7225 65.5375 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.7625 65.4025 144.8975 65.5375 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.9375 65.4025 146.0725 65.5375 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.1125 65.4025 147.2475 65.5375 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.2875 65.4025 148.4225 65.5375 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.4625 65.4025 149.5975 65.5375 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.6375 65.4025 150.7725 65.5375 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.8125 65.4025 151.9475 65.5375 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.9875 65.4025 153.1225 65.5375 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.1625 65.4025 154.2975 65.5375 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.3375 65.4025 155.4725 65.5375 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.5125 65.4025 156.6475 65.5375 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.6875 65.4025 157.8225 65.5375 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.8625 65.4025 158.9975 65.5375 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.0375 65.4025 160.1725 65.5375 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.2125 65.4025 161.3475 65.5375 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.3875 65.4025 162.5225 65.5375 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.5625 65.4025 163.6975 65.5375 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.7375 65.4025 164.8725 65.5375 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.9125 65.4025 166.0475 65.5375 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.0875 65.4025 167.2225 65.5375 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.2625 65.4025 168.3975 65.5375 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.4375 65.4025 169.5725 65.5375 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.6125 65.4025 170.7475 65.5375 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.7875 65.4025 171.9225 65.5375 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.9625 65.4025 173.0975 65.5375 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.1375 65.4025 174.2725 65.5375 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.3125 65.4025 175.4475 65.5375 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.4875 65.4025 176.6225 65.5375 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.6625 65.4025 177.7975 65.5375 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.8375 65.4025 178.9725 65.5375 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.0125 65.4025 180.1475 65.5375 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.1875 65.4025 181.3225 65.5375 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.3625 65.4025 182.4975 65.5375 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.5375 65.4025 183.6725 65.5375 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.7125 65.4025 184.8475 65.5375 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.8875 65.4025 186.0225 65.5375 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.0625 65.4025 187.1975 65.5375 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.2375 65.4025 188.3725 65.5375 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.4125 65.4025 189.5475 65.5375 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.5875 65.4025 190.7225 65.5375 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.7625 65.4025 191.8975 65.5375 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.9375 65.4025 193.0725 65.5375 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.1125 65.4025 194.2475 65.5375 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.2875 65.4025 195.4225 65.5375 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.4625 65.4025 196.5975 65.5375 ;
      END
   END dout1[119]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  40.5575 32.77 40.6925 32.905 ;
         LAYER metal4 ;
         RECT  53.385 28.1025 53.525 58.2525 ;
         LAYER metal4 ;
         RECT  253.8475 41.1025 253.9875 63.505 ;
         LAYER metal3 ;
         RECT  166.2975 2.47 166.4325 2.605 ;
         LAYER metal4 ;
         RECT  200.815 28.1025 200.955 58.2525 ;
         LAYER metal3 ;
         RECT  213.6475 41.74 213.7825 41.875 ;
         LAYER metal3 ;
         RECT  45.825 30.5675 45.96 30.7025 ;
         LAYER metal3 ;
         RECT  97.6575 2.47 97.7925 2.605 ;
         LAYER metal3 ;
         RECT  252.115 70.745 252.25 70.88 ;
         LAYER metal4 ;
         RECT  0.6875 20.45 0.8275 42.8525 ;
         LAYER metal3 ;
         RECT  86.2175 2.47 86.3525 2.605 ;
         LAYER metal3 ;
         RECT  213.6475 32.77 213.7825 32.905 ;
         LAYER metal3 ;
         RECT  246.3775 2.47 246.5125 2.605 ;
         LAYER metal4 ;
         RECT  34.735 46.2225 34.875 56.2425 ;
         LAYER metal3 ;
         RECT  223.4975 2.47 223.6325 2.605 ;
         LAYER metal3 ;
         RECT  212.0575 2.47 212.1925 2.605 ;
         LAYER metal3 ;
         RECT  120.5375 2.47 120.6725 2.605 ;
         LAYER metal3 ;
         RECT  53.4525 21.9725 197.2675 22.0425 ;
         LAYER metal3 ;
         RECT  2.425 13.075 2.56 13.21 ;
         LAYER metal3 ;
         RECT  269.2575 2.47 269.3925 2.605 ;
         LAYER metal3 ;
         RECT  177.7375 2.47 177.8725 2.605 ;
         LAYER metal3 ;
         RECT  131.9775 2.47 132.1125 2.605 ;
         LAYER metal3 ;
         RECT  303.5775 2.47 303.7125 2.605 ;
         LAYER metal4 ;
         RECT  52.305 31.2725 52.445 55.3325 ;
         LAYER metal3 ;
         RECT  257.8175 2.47 257.9525 2.605 ;
         LAYER metal3 ;
         RECT  201.8975 56.69 202.0325 56.825 ;
         LAYER metal3 ;
         RECT  234.9375 2.47 235.0725 2.605 ;
         LAYER metal3 ;
         RECT  74.7775 2.47 74.9125 2.605 ;
         LAYER metal3 ;
         RECT  326.4575 2.47 326.5925 2.605 ;
         LAYER metal3 ;
         RECT  53.4525 62.845 197.2675 62.915 ;
         LAYER metal4 ;
         RECT  219.66 21.3925 219.8 31.4125 ;
         LAYER metal3 ;
         RECT  200.6175 2.47 200.7525 2.605 ;
         LAYER metal3 ;
         RECT  208.38 55.9025 208.515 56.0375 ;
         LAYER metal4 ;
         RECT  45.205 31.2725 45.345 55.4025 ;
         LAYER metal4 ;
         RECT  216.94 60.8625 217.08 70.8825 ;
         LAYER metal3 ;
         RECT  154.8575 2.47 154.9925 2.605 ;
         LAYER metal3 ;
         RECT  53.4525 27.4075 197.7375 27.4775 ;
         LAYER metal3 ;
         RECT  63.3375 2.47 63.4725 2.605 ;
         LAYER metal4 ;
         RECT  208.995 31.2725 209.135 55.4025 ;
         LAYER metal3 ;
         RECT  51.8975 2.47 52.0325 2.605 ;
         LAYER metal3 ;
         RECT  52.3075 29.78 52.4425 29.915 ;
         LAYER metal3 ;
         RECT  40.5575 35.76 40.6925 35.895 ;
         LAYER metal4 ;
         RECT  201.895 31.2725 202.035 55.3325 ;
         LAYER metal3 ;
         RECT  292.1375 2.47 292.2725 2.605 ;
         LAYER metal3 ;
         RECT  109.0975 2.47 109.2325 2.605 ;
         LAYER metal3 ;
         RECT  143.4175 2.47 143.5525 2.605 ;
         LAYER metal3 ;
         RECT  213.6475 44.73 213.7825 44.865 ;
         LAYER metal3 ;
         RECT  40.4575 2.47 40.5925 2.605 ;
         LAYER metal3 ;
         RECT  213.6475 35.76 213.7825 35.895 ;
         LAYER metal3 ;
         RECT  53.4525 58.9475 198.9125 59.0175 ;
         LAYER metal3 ;
         RECT  372.2175 2.47 372.3525 2.605 ;
         LAYER metal4 ;
         RECT  37.455 13.0725 37.595 28.0325 ;
         LAYER metal3 ;
         RECT  280.6975 2.47 280.8325 2.605 ;
         LAYER metal3 ;
         RECT  315.0175 2.47 315.1525 2.605 ;
         LAYER metal3 ;
         RECT  189.1775 2.47 189.3125 2.605 ;
         LAYER metal3 ;
         RECT  40.5575 44.73 40.6925 44.865 ;
         LAYER metal3 ;
         RECT  349.3375 2.47 349.4725 2.605 ;
         LAYER metal3 ;
         RECT  337.8975 2.47 338.0325 2.605 ;
         LAYER metal3 ;
         RECT  40.5575 41.74 40.6925 41.875 ;
         LAYER metal3 ;
         RECT  360.7775 2.47 360.9125 2.605 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  2.75 20.4825 2.89 42.885 ;
         LAYER metal3 ;
         RECT  363.6375 0.0 363.7725 0.135 ;
         LAYER metal4 ;
         RECT  6.105 10.6025 6.245 25.5625 ;
         LAYER metal3 ;
         RECT  39.03 37.255 39.165 37.39 ;
         LAYER metal4 ;
         RECT  248.29 58.3925 248.43 73.3525 ;
         LAYER metal3 ;
         RECT  272.1175 0.0 272.2525 0.135 ;
         LAYER metal3 ;
         RECT  39.03 40.245 39.165 40.38 ;
         LAYER metal3 ;
         RECT  340.7575 0.0 340.8925 0.135 ;
         LAYER metal3 ;
         RECT  306.4375 0.0 306.5725 0.135 ;
         LAYER metal3 ;
         RECT  66.1975 0.0 66.3325 0.135 ;
         LAYER metal3 ;
         RECT  39.03 31.275 39.165 31.41 ;
         LAYER metal3 ;
         RECT  252.115 73.215 252.25 73.35 ;
         LAYER metal3 ;
         RECT  375.0775 0.0 375.2125 0.135 ;
         LAYER metal3 ;
         RECT  54.7575 0.0 54.8925 0.135 ;
         LAYER metal3 ;
         RECT  317.8775 0.0 318.0125 0.135 ;
         LAYER metal3 ;
         RECT  157.7175 0.0 157.8525 0.135 ;
         LAYER metal3 ;
         RECT  180.5975 0.0 180.7325 0.135 ;
         LAYER metal3 ;
         RECT  294.9975 0.0 295.1325 0.135 ;
         LAYER metal3 ;
         RECT  2.425 10.605 2.56 10.74 ;
         LAYER metal3 ;
         RECT  134.8375 0.0 134.9725 0.135 ;
         LAYER metal3 ;
         RECT  111.9575 0.0 112.0925 0.135 ;
         LAYER metal3 ;
         RECT  53.4525 24.0225 197.2675 24.0925 ;
         LAYER metal4 ;
         RECT  251.785 41.07 251.925 63.4725 ;
         LAYER metal4 ;
         RECT  45.765 31.24 45.905 55.365 ;
         LAYER metal3 ;
         RECT  215.175 37.255 215.31 37.39 ;
         LAYER metal4 ;
         RECT  37.595 46.1575 37.735 56.3075 ;
         LAYER metal4 ;
         RECT  200.355 28.1025 200.495 58.2525 ;
         LAYER metal3 ;
         RECT  249.2375 0.0 249.3725 0.135 ;
         LAYER metal3 ;
         RECT  192.0375 0.0 192.1725 0.135 ;
         LAYER metal3 ;
         RECT  329.3175 0.0 329.4525 0.135 ;
         LAYER metal4 ;
         RECT  216.8 21.3275 216.94 31.4775 ;
         LAYER metal4 ;
         RECT  208.435 31.24 208.575 55.365 ;
         LAYER metal3 ;
         RECT  123.3975 0.0 123.5325 0.135 ;
         LAYER metal3 ;
         RECT  283.5575 0.0 283.6925 0.135 ;
         LAYER metal3 ;
         RECT  100.5175 0.0 100.6525 0.135 ;
         LAYER metal3 ;
         RECT  39.03 34.265 39.165 34.4 ;
         LAYER metal3 ;
         RECT  260.6775 0.0 260.8125 0.135 ;
         LAYER metal3 ;
         RECT  169.1575 0.0 169.2925 0.135 ;
         LAYER metal3 ;
         RECT  215.175 43.235 215.31 43.37 ;
         LAYER metal3 ;
         RECT  214.9175 0.0 215.0525 0.135 ;
         LAYER metal4 ;
         RECT  53.845 28.1025 53.985 58.2525 ;
         LAYER metal3 ;
         RECT  39.03 46.225 39.165 46.36 ;
         LAYER metal4 ;
         RECT  43.615 31.24 43.755 55.4025 ;
         LAYER metal3 ;
         RECT  89.0775 0.0 89.2125 0.135 ;
         LAYER metal3 ;
         RECT  215.175 40.245 215.31 40.38 ;
         LAYER metal3 ;
         RECT  53.4525 60.9525 197.3025 61.0225 ;
         LAYER metal3 ;
         RECT  215.175 31.275 215.31 31.41 ;
         LAYER metal3 ;
         RECT  237.7975 0.0 237.9325 0.135 ;
         LAYER metal3 ;
         RECT  146.2775 0.0 146.4125 0.135 ;
         LAYER metal3 ;
         RECT  226.3575 0.0 226.4925 0.135 ;
         LAYER metal3 ;
         RECT  352.1975 0.0 352.3325 0.135 ;
         LAYER metal3 ;
         RECT  215.175 34.265 215.31 34.4 ;
         LAYER metal3 ;
         RECT  215.175 46.225 215.31 46.36 ;
         LAYER metal3 ;
         RECT  43.3175 0.0 43.4525 0.135 ;
         LAYER metal3 ;
         RECT  203.4775 0.0 203.6125 0.135 ;
         LAYER metal3 ;
         RECT  77.6375 0.0 77.7725 0.135 ;
         LAYER metal4 ;
         RECT  210.585 31.24 210.725 55.4025 ;
         LAYER metal3 ;
         RECT  39.03 43.235 39.165 43.37 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 383.585 73.2125 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 383.585 73.2125 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 40.6 0.965 ;
      RECT  0.14 0.965 40.6 1.38 ;
      RECT  40.6 0.14 41.015 0.965 ;
      RECT  41.015 0.965 43.46 1.38 ;
      RECT  43.875 0.965 46.32 1.38 ;
      RECT  46.735 0.965 49.18 1.38 ;
      RECT  49.595 0.965 52.04 1.38 ;
      RECT  52.455 0.965 54.9 1.38 ;
      RECT  55.315 0.965 57.76 1.38 ;
      RECT  58.175 0.965 60.62 1.38 ;
      RECT  61.035 0.965 63.48 1.38 ;
      RECT  63.895 0.965 66.34 1.38 ;
      RECT  66.755 0.965 69.2 1.38 ;
      RECT  69.615 0.965 72.06 1.38 ;
      RECT  72.475 0.965 74.92 1.38 ;
      RECT  75.335 0.965 77.78 1.38 ;
      RECT  78.195 0.965 80.64 1.38 ;
      RECT  81.055 0.965 83.5 1.38 ;
      RECT  83.915 0.965 86.36 1.38 ;
      RECT  86.775 0.965 89.22 1.38 ;
      RECT  89.635 0.965 92.08 1.38 ;
      RECT  92.495 0.965 94.94 1.38 ;
      RECT  95.355 0.965 97.8 1.38 ;
      RECT  98.215 0.965 100.66 1.38 ;
      RECT  101.075 0.965 103.52 1.38 ;
      RECT  103.935 0.965 106.38 1.38 ;
      RECT  106.795 0.965 109.24 1.38 ;
      RECT  109.655 0.965 112.1 1.38 ;
      RECT  112.515 0.965 114.96 1.38 ;
      RECT  115.375 0.965 117.82 1.38 ;
      RECT  118.235 0.965 120.68 1.38 ;
      RECT  121.095 0.965 123.54 1.38 ;
      RECT  123.955 0.965 126.4 1.38 ;
      RECT  126.815 0.965 129.26 1.38 ;
      RECT  129.675 0.965 132.12 1.38 ;
      RECT  132.535 0.965 134.98 1.38 ;
      RECT  135.395 0.965 137.84 1.38 ;
      RECT  138.255 0.965 140.7 1.38 ;
      RECT  141.115 0.965 143.56 1.38 ;
      RECT  143.975 0.965 146.42 1.38 ;
      RECT  146.835 0.965 149.28 1.38 ;
      RECT  149.695 0.965 152.14 1.38 ;
      RECT  152.555 0.965 155.0 1.38 ;
      RECT  155.415 0.965 157.86 1.38 ;
      RECT  158.275 0.965 160.72 1.38 ;
      RECT  161.135 0.965 163.58 1.38 ;
      RECT  163.995 0.965 166.44 1.38 ;
      RECT  166.855 0.965 169.3 1.38 ;
      RECT  169.715 0.965 172.16 1.38 ;
      RECT  172.575 0.965 175.02 1.38 ;
      RECT  175.435 0.965 177.88 1.38 ;
      RECT  178.295 0.965 180.74 1.38 ;
      RECT  181.155 0.965 183.6 1.38 ;
      RECT  184.015 0.965 186.46 1.38 ;
      RECT  186.875 0.965 189.32 1.38 ;
      RECT  189.735 0.965 192.18 1.38 ;
      RECT  192.595 0.965 195.04 1.38 ;
      RECT  195.455 0.965 197.9 1.38 ;
      RECT  198.315 0.965 200.76 1.38 ;
      RECT  201.175 0.965 203.62 1.38 ;
      RECT  204.035 0.965 206.48 1.38 ;
      RECT  206.895 0.965 209.34 1.38 ;
      RECT  209.755 0.965 212.2 1.38 ;
      RECT  212.615 0.965 215.06 1.38 ;
      RECT  215.475 0.965 217.92 1.38 ;
      RECT  218.335 0.965 220.78 1.38 ;
      RECT  221.195 0.965 223.64 1.38 ;
      RECT  224.055 0.965 226.5 1.38 ;
      RECT  226.915 0.965 229.36 1.38 ;
      RECT  229.775 0.965 232.22 1.38 ;
      RECT  232.635 0.965 235.08 1.38 ;
      RECT  235.495 0.965 237.94 1.38 ;
      RECT  238.355 0.965 240.8 1.38 ;
      RECT  241.215 0.965 243.66 1.38 ;
      RECT  244.075 0.965 246.52 1.38 ;
      RECT  246.935 0.965 249.38 1.38 ;
      RECT  249.795 0.965 252.24 1.38 ;
      RECT  252.655 0.965 255.1 1.38 ;
      RECT  255.515 0.965 257.96 1.38 ;
      RECT  258.375 0.965 260.82 1.38 ;
      RECT  261.235 0.965 263.68 1.38 ;
      RECT  264.095 0.965 266.54 1.38 ;
      RECT  266.955 0.965 269.4 1.38 ;
      RECT  269.815 0.965 272.26 1.38 ;
      RECT  272.675 0.965 275.12 1.38 ;
      RECT  275.535 0.965 277.98 1.38 ;
      RECT  278.395 0.965 280.84 1.38 ;
      RECT  281.255 0.965 283.7 1.38 ;
      RECT  284.115 0.965 286.56 1.38 ;
      RECT  286.975 0.965 289.42 1.38 ;
      RECT  289.835 0.965 292.28 1.38 ;
      RECT  292.695 0.965 295.14 1.38 ;
      RECT  295.555 0.965 298.0 1.38 ;
      RECT  298.415 0.965 300.86 1.38 ;
      RECT  301.275 0.965 303.72 1.38 ;
      RECT  304.135 0.965 306.58 1.38 ;
      RECT  306.995 0.965 309.44 1.38 ;
      RECT  309.855 0.965 312.3 1.38 ;
      RECT  312.715 0.965 315.16 1.38 ;
      RECT  315.575 0.965 318.02 1.38 ;
      RECT  318.435 0.965 320.88 1.38 ;
      RECT  321.295 0.965 323.74 1.38 ;
      RECT  324.155 0.965 326.6 1.38 ;
      RECT  327.015 0.965 329.46 1.38 ;
      RECT  329.875 0.965 332.32 1.38 ;
      RECT  332.735 0.965 335.18 1.38 ;
      RECT  335.595 0.965 338.04 1.38 ;
      RECT  338.455 0.965 340.9 1.38 ;
      RECT  341.315 0.965 343.76 1.38 ;
      RECT  344.175 0.965 346.62 1.38 ;
      RECT  347.035 0.965 349.48 1.38 ;
      RECT  349.895 0.965 352.34 1.38 ;
      RECT  352.755 0.965 355.2 1.38 ;
      RECT  355.615 0.965 358.06 1.38 ;
      RECT  358.475 0.965 360.92 1.38 ;
      RECT  361.335 0.965 363.78 1.38 ;
      RECT  364.195 0.965 366.64 1.38 ;
      RECT  367.055 0.965 369.5 1.38 ;
      RECT  369.915 0.965 372.36 1.38 ;
      RECT  372.775 0.965 375.22 1.38 ;
      RECT  375.635 0.965 378.08 1.38 ;
      RECT  378.495 0.965 380.94 1.38 ;
      RECT  381.355 0.965 383.585 1.38 ;
      RECT  0.14 47.19 34.88 47.605 ;
      RECT  0.14 47.605 34.88 73.2125 ;
      RECT  34.88 1.38 35.295 47.19 ;
      RECT  35.295 47.19 40.6 47.605 ;
      RECT  35.295 47.605 40.6 73.2125 ;
      RECT  34.88 47.605 35.295 49.92 ;
      RECT  34.88 50.335 35.295 52.13 ;
      RECT  34.88 52.545 35.295 54.86 ;
      RECT  34.88 55.275 35.295 73.2125 ;
      RECT  219.24 30.445 219.655 73.2125 ;
      RECT  219.655 30.03 383.585 30.445 ;
      RECT  219.24 27.715 219.655 30.03 ;
      RECT  219.24 25.505 219.655 27.3 ;
      RECT  219.24 1.38 219.655 22.36 ;
      RECT  219.24 22.775 219.655 25.09 ;
      RECT  0.14 1.38 0.145 11.57 ;
      RECT  0.14 11.57 0.145 11.985 ;
      RECT  0.14 11.985 0.145 47.19 ;
      RECT  0.145 1.38 0.56 11.57 ;
      RECT  0.145 11.985 0.56 47.19 ;
      RECT  254.115 30.445 254.53 71.97 ;
      RECT  254.115 72.385 254.53 73.2125 ;
      RECT  254.53 30.445 383.585 71.97 ;
      RECT  254.53 71.97 383.585 72.385 ;
      RECT  254.53 72.385 383.585 73.2125 ;
      RECT  0.56 11.57 6.1075 11.655 ;
      RECT  0.56 11.655 6.1075 11.985 ;
      RECT  6.1075 11.57 6.5225 11.655 ;
      RECT  6.5225 11.57 34.88 11.655 ;
      RECT  6.5225 11.655 34.88 11.985 ;
      RECT  0.56 11.985 6.1075 12.07 ;
      RECT  6.1075 12.07 6.5225 47.19 ;
      RECT  6.5225 11.985 34.88 12.07 ;
      RECT  6.5225 12.07 34.88 47.19 ;
      RECT  219.655 30.445 248.0125 71.885 ;
      RECT  219.655 71.885 248.0125 71.97 ;
      RECT  248.0125 30.445 248.4275 71.885 ;
      RECT  248.4275 71.885 254.115 71.97 ;
      RECT  219.655 71.97 248.0125 72.3 ;
      RECT  219.655 72.3 248.0125 72.385 ;
      RECT  248.0125 72.3 248.4275 72.385 ;
      RECT  248.4275 71.97 254.115 72.3 ;
      RECT  248.4275 72.3 254.115 72.385 ;
      RECT  41.015 65.2625 56.4975 65.6775 ;
      RECT  41.015 65.6775 56.4975 73.2125 ;
      RECT  56.4975 65.6775 56.9125 73.2125 ;
      RECT  56.9125 65.6775 219.24 73.2125 ;
      RECT  56.9125 65.2625 57.6725 65.6775 ;
      RECT  58.0875 65.2625 58.8475 65.6775 ;
      RECT  59.2625 65.2625 60.0225 65.6775 ;
      RECT  60.4375 65.2625 61.1975 65.6775 ;
      RECT  61.6125 65.2625 62.3725 65.6775 ;
      RECT  62.7875 65.2625 63.5475 65.6775 ;
      RECT  63.9625 65.2625 64.7225 65.6775 ;
      RECT  65.1375 65.2625 65.8975 65.6775 ;
      RECT  66.3125 65.2625 67.0725 65.6775 ;
      RECT  67.4875 65.2625 68.2475 65.6775 ;
      RECT  68.6625 65.2625 69.4225 65.6775 ;
      RECT  69.8375 65.2625 70.5975 65.6775 ;
      RECT  71.0125 65.2625 71.7725 65.6775 ;
      RECT  72.1875 65.2625 72.9475 65.6775 ;
      RECT  73.3625 65.2625 74.1225 65.6775 ;
      RECT  74.5375 65.2625 75.2975 65.6775 ;
      RECT  75.7125 65.2625 76.4725 65.6775 ;
      RECT  76.8875 65.2625 77.6475 65.6775 ;
      RECT  78.0625 65.2625 78.8225 65.6775 ;
      RECT  79.2375 65.2625 79.9975 65.6775 ;
      RECT  80.4125 65.2625 81.1725 65.6775 ;
      RECT  81.5875 65.2625 82.3475 65.6775 ;
      RECT  82.7625 65.2625 83.5225 65.6775 ;
      RECT  83.9375 65.2625 84.6975 65.6775 ;
      RECT  85.1125 65.2625 85.8725 65.6775 ;
      RECT  86.2875 65.2625 87.0475 65.6775 ;
      RECT  87.4625 65.2625 88.2225 65.6775 ;
      RECT  88.6375 65.2625 89.3975 65.6775 ;
      RECT  89.8125 65.2625 90.5725 65.6775 ;
      RECT  90.9875 65.2625 91.7475 65.6775 ;
      RECT  92.1625 65.2625 92.9225 65.6775 ;
      RECT  93.3375 65.2625 94.0975 65.6775 ;
      RECT  94.5125 65.2625 95.2725 65.6775 ;
      RECT  95.6875 65.2625 96.4475 65.6775 ;
      RECT  96.8625 65.2625 97.6225 65.6775 ;
      RECT  98.0375 65.2625 98.7975 65.6775 ;
      RECT  99.2125 65.2625 99.9725 65.6775 ;
      RECT  100.3875 65.2625 101.1475 65.6775 ;
      RECT  101.5625 65.2625 102.3225 65.6775 ;
      RECT  102.7375 65.2625 103.4975 65.6775 ;
      RECT  103.9125 65.2625 104.6725 65.6775 ;
      RECT  105.0875 65.2625 105.8475 65.6775 ;
      RECT  106.2625 65.2625 107.0225 65.6775 ;
      RECT  107.4375 65.2625 108.1975 65.6775 ;
      RECT  108.6125 65.2625 109.3725 65.6775 ;
      RECT  109.7875 65.2625 110.5475 65.6775 ;
      RECT  110.9625 65.2625 111.7225 65.6775 ;
      RECT  112.1375 65.2625 112.8975 65.6775 ;
      RECT  113.3125 65.2625 114.0725 65.6775 ;
      RECT  114.4875 65.2625 115.2475 65.6775 ;
      RECT  115.6625 65.2625 116.4225 65.6775 ;
      RECT  116.8375 65.2625 117.5975 65.6775 ;
      RECT  118.0125 65.2625 118.7725 65.6775 ;
      RECT  119.1875 65.2625 119.9475 65.6775 ;
      RECT  120.3625 65.2625 121.1225 65.6775 ;
      RECT  121.5375 65.2625 122.2975 65.6775 ;
      RECT  122.7125 65.2625 123.4725 65.6775 ;
      RECT  123.8875 65.2625 124.6475 65.6775 ;
      RECT  125.0625 65.2625 125.8225 65.6775 ;
      RECT  126.2375 65.2625 126.9975 65.6775 ;
      RECT  127.4125 65.2625 128.1725 65.6775 ;
      RECT  128.5875 65.2625 129.3475 65.6775 ;
      RECT  129.7625 65.2625 130.5225 65.6775 ;
      RECT  130.9375 65.2625 131.6975 65.6775 ;
      RECT  132.1125 65.2625 132.8725 65.6775 ;
      RECT  133.2875 65.2625 134.0475 65.6775 ;
      RECT  134.4625 65.2625 135.2225 65.6775 ;
      RECT  135.6375 65.2625 136.3975 65.6775 ;
      RECT  136.8125 65.2625 137.5725 65.6775 ;
      RECT  137.9875 65.2625 138.7475 65.6775 ;
      RECT  139.1625 65.2625 139.9225 65.6775 ;
      RECT  140.3375 65.2625 141.0975 65.6775 ;
      RECT  141.5125 65.2625 142.2725 65.6775 ;
      RECT  142.6875 65.2625 143.4475 65.6775 ;
      RECT  143.8625 65.2625 144.6225 65.6775 ;
      RECT  145.0375 65.2625 145.7975 65.6775 ;
      RECT  146.2125 65.2625 146.9725 65.6775 ;
      RECT  147.3875 65.2625 148.1475 65.6775 ;
      RECT  148.5625 65.2625 149.3225 65.6775 ;
      RECT  149.7375 65.2625 150.4975 65.6775 ;
      RECT  150.9125 65.2625 151.6725 65.6775 ;
      RECT  152.0875 65.2625 152.8475 65.6775 ;
      RECT  153.2625 65.2625 154.0225 65.6775 ;
      RECT  154.4375 65.2625 155.1975 65.6775 ;
      RECT  155.6125 65.2625 156.3725 65.6775 ;
      RECT  156.7875 65.2625 157.5475 65.6775 ;
      RECT  157.9625 65.2625 158.7225 65.6775 ;
      RECT  159.1375 65.2625 159.8975 65.6775 ;
      RECT  160.3125 65.2625 161.0725 65.6775 ;
      RECT  161.4875 65.2625 162.2475 65.6775 ;
      RECT  162.6625 65.2625 163.4225 65.6775 ;
      RECT  163.8375 65.2625 164.5975 65.6775 ;
      RECT  165.0125 65.2625 165.7725 65.6775 ;
      RECT  166.1875 65.2625 166.9475 65.6775 ;
      RECT  167.3625 65.2625 168.1225 65.6775 ;
      RECT  168.5375 65.2625 169.2975 65.6775 ;
      RECT  169.7125 65.2625 170.4725 65.6775 ;
      RECT  170.8875 65.2625 171.6475 65.6775 ;
      RECT  172.0625 65.2625 172.8225 65.6775 ;
      RECT  173.2375 65.2625 173.9975 65.6775 ;
      RECT  174.4125 65.2625 175.1725 65.6775 ;
      RECT  175.5875 65.2625 176.3475 65.6775 ;
      RECT  176.7625 65.2625 177.5225 65.6775 ;
      RECT  177.9375 65.2625 178.6975 65.6775 ;
      RECT  179.1125 65.2625 179.8725 65.6775 ;
      RECT  180.2875 65.2625 181.0475 65.6775 ;
      RECT  181.4625 65.2625 182.2225 65.6775 ;
      RECT  182.6375 65.2625 183.3975 65.6775 ;
      RECT  183.8125 65.2625 184.5725 65.6775 ;
      RECT  184.9875 65.2625 185.7475 65.6775 ;
      RECT  186.1625 65.2625 186.9225 65.6775 ;
      RECT  187.3375 65.2625 188.0975 65.6775 ;
      RECT  188.5125 65.2625 189.2725 65.6775 ;
      RECT  189.6875 65.2625 190.4475 65.6775 ;
      RECT  190.8625 65.2625 191.6225 65.6775 ;
      RECT  192.0375 65.2625 192.7975 65.6775 ;
      RECT  193.2125 65.2625 193.9725 65.6775 ;
      RECT  194.3875 65.2625 195.1475 65.6775 ;
      RECT  195.5625 65.2625 196.3225 65.6775 ;
      RECT  196.7375 65.2625 219.24 65.6775 ;
      RECT  40.8325 1.38 41.015 32.63 ;
      RECT  40.8325 32.63 41.015 33.045 ;
      RECT  40.8325 33.045 41.015 73.2125 ;
      RECT  35.295 32.63 40.4175 33.045 ;
      RECT  41.015 1.38 166.1575 2.33 ;
      RECT  166.1575 1.38 166.5725 2.33 ;
      RECT  166.5725 1.38 219.24 2.33 ;
      RECT  56.9125 30.445 213.5075 41.6 ;
      RECT  56.9125 41.6 213.5075 42.015 ;
      RECT  213.9225 41.6 219.24 42.015 ;
      RECT  41.015 30.03 45.685 30.4275 ;
      RECT  41.015 30.4275 45.685 30.445 ;
      RECT  45.685 30.03 46.1 30.4275 ;
      RECT  46.1 30.4275 219.24 30.445 ;
      RECT  41.015 30.445 45.685 30.8425 ;
      RECT  41.015 30.8425 45.685 65.2625 ;
      RECT  45.685 30.8425 46.1 65.2625 ;
      RECT  46.1 30.445 56.4975 30.8425 ;
      RECT  248.4275 30.445 251.975 70.605 ;
      RECT  248.4275 70.605 251.975 71.02 ;
      RECT  248.4275 71.02 251.975 71.885 ;
      RECT  251.975 30.445 252.39 70.605 ;
      RECT  251.975 71.02 252.39 71.885 ;
      RECT  252.39 30.445 254.115 70.605 ;
      RECT  252.39 70.605 254.115 71.02 ;
      RECT  252.39 71.02 254.115 71.885 ;
      RECT  86.4925 2.33 97.5175 2.745 ;
      RECT  213.5075 30.445 213.9225 32.63 ;
      RECT  219.655 1.38 246.2375 2.33 ;
      RECT  219.655 2.745 246.2375 30.03 ;
      RECT  246.2375 1.38 246.6525 2.33 ;
      RECT  246.2375 2.745 246.6525 30.03 ;
      RECT  246.6525 1.38 383.585 2.33 ;
      RECT  246.6525 2.745 383.585 30.03 ;
      RECT  219.655 2.33 223.3575 2.745 ;
      RECT  212.3325 2.33 219.24 2.745 ;
      RECT  41.015 2.745 53.3125 21.8325 ;
      RECT  41.015 21.8325 53.3125 22.1825 ;
      RECT  53.3125 2.745 166.1575 21.8325 ;
      RECT  166.1575 2.745 166.5725 21.8325 ;
      RECT  166.5725 2.745 197.4075 21.8325 ;
      RECT  197.4075 2.745 219.24 21.8325 ;
      RECT  197.4075 21.8325 219.24 22.1825 ;
      RECT  0.56 12.07 2.285 12.935 ;
      RECT  0.56 12.935 2.285 13.35 ;
      RECT  0.56 13.35 2.285 47.19 ;
      RECT  2.285 12.07 2.7 12.935 ;
      RECT  2.285 13.35 2.7 47.19 ;
      RECT  2.7 12.07 6.1075 12.935 ;
      RECT  2.7 12.935 6.1075 13.35 ;
      RECT  2.7 13.35 6.1075 47.19 ;
      RECT  166.5725 2.33 177.5975 2.745 ;
      RECT  120.8125 2.33 131.8375 2.745 ;
      RECT  246.6525 2.33 257.6775 2.745 ;
      RECT  258.0925 2.33 269.1175 2.745 ;
      RECT  56.9125 42.015 201.7575 56.55 ;
      RECT  56.9125 56.55 201.7575 56.965 ;
      RECT  201.7575 42.015 202.1725 56.55 ;
      RECT  201.7575 56.965 202.1725 65.2625 ;
      RECT  202.1725 56.55 213.5075 56.965 ;
      RECT  202.1725 56.965 213.5075 65.2625 ;
      RECT  223.7725 2.33 234.7975 2.745 ;
      RECT  235.2125 2.33 246.2375 2.745 ;
      RECT  75.0525 2.33 86.0775 2.745 ;
      RECT  56.4975 63.055 56.9125 65.2625 ;
      RECT  46.1 30.8425 53.3125 62.705 ;
      RECT  46.1 62.705 53.3125 63.055 ;
      RECT  46.1 63.055 53.3125 65.2625 ;
      RECT  53.3125 63.055 56.4975 65.2625 ;
      RECT  56.9125 63.055 197.4075 65.2625 ;
      RECT  197.4075 62.705 201.7575 63.055 ;
      RECT  197.4075 63.055 201.7575 65.2625 ;
      RECT  200.8925 2.33 211.9175 2.745 ;
      RECT  202.1725 42.015 208.24 55.7625 ;
      RECT  202.1725 55.7625 208.24 56.1775 ;
      RECT  202.1725 56.1775 208.24 56.55 ;
      RECT  208.24 42.015 208.655 55.7625 ;
      RECT  208.24 56.1775 208.655 56.55 ;
      RECT  208.655 42.015 213.5075 55.7625 ;
      RECT  208.655 55.7625 213.5075 56.1775 ;
      RECT  208.655 56.1775 213.5075 56.55 ;
      RECT  155.1325 2.33 166.1575 2.745 ;
      RECT  53.3125 27.6175 166.1575 30.03 ;
      RECT  166.1575 27.6175 166.5725 30.03 ;
      RECT  166.5725 27.6175 197.4075 30.03 ;
      RECT  197.4075 22.1825 197.8775 27.2675 ;
      RECT  197.4075 27.6175 197.8775 30.03 ;
      RECT  197.8775 22.1825 219.24 27.2675 ;
      RECT  197.8775 27.2675 219.24 27.6175 ;
      RECT  197.8775 27.6175 219.24 30.03 ;
      RECT  63.6125 2.33 74.6375 2.745 ;
      RECT  41.015 2.33 51.7575 2.745 ;
      RECT  52.1725 2.33 63.1975 2.745 ;
      RECT  46.1 30.03 52.1675 30.055 ;
      RECT  46.1 30.055 52.1675 30.4275 ;
      RECT  52.1675 30.055 52.5825 30.4275 ;
      RECT  52.5825 30.03 219.24 30.055 ;
      RECT  52.5825 30.055 219.24 30.4275 ;
      RECT  41.015 22.1825 52.1675 29.64 ;
      RECT  41.015 29.64 52.1675 30.03 ;
      RECT  52.1675 22.1825 52.5825 29.64 ;
      RECT  52.5825 22.1825 53.3125 29.64 ;
      RECT  52.5825 29.64 53.3125 30.03 ;
      RECT  40.6 33.045 40.8325 35.62 ;
      RECT  40.4175 33.045 40.6 35.62 ;
      RECT  292.4125 2.33 303.4375 2.745 ;
      RECT  97.9325 2.33 108.9575 2.745 ;
      RECT  109.3725 2.33 120.3975 2.745 ;
      RECT  132.2525 2.33 143.2775 2.745 ;
      RECT  143.6925 2.33 154.7175 2.745 ;
      RECT  213.5075 42.015 213.9225 44.59 ;
      RECT  213.5075 45.005 213.9225 65.2625 ;
      RECT  40.6 1.38 40.7325 2.33 ;
      RECT  40.6 2.745 40.7325 32.63 ;
      RECT  40.7325 1.38 40.8325 2.33 ;
      RECT  40.7325 2.33 40.8325 2.745 ;
      RECT  40.7325 2.745 40.8325 32.63 ;
      RECT  35.295 1.38 40.3175 2.33 ;
      RECT  35.295 2.33 40.3175 2.745 ;
      RECT  40.3175 1.38 40.4175 2.33 ;
      RECT  40.3175 2.745 40.4175 32.63 ;
      RECT  40.4175 1.38 40.6 2.33 ;
      RECT  40.4175 2.745 40.6 32.63 ;
      RECT  213.5075 33.045 213.9225 35.62 ;
      RECT  213.5075 36.035 213.9225 41.6 ;
      RECT  56.4975 30.445 56.9125 58.8075 ;
      RECT  53.3125 30.8425 56.4975 58.8075 ;
      RECT  56.9125 56.965 197.4075 58.8075 ;
      RECT  197.4075 56.965 199.0525 58.8075 ;
      RECT  199.0525 56.965 201.7575 58.8075 ;
      RECT  199.0525 58.8075 201.7575 59.1575 ;
      RECT  199.0525 59.1575 201.7575 62.705 ;
      RECT  372.4925 2.33 383.585 2.745 ;
      RECT  269.5325 2.33 280.5575 2.745 ;
      RECT  280.9725 2.33 291.9975 2.745 ;
      RECT  303.8525 2.33 314.8775 2.745 ;
      RECT  315.2925 2.33 326.3175 2.745 ;
      RECT  178.0125 2.33 189.0375 2.745 ;
      RECT  189.4525 2.33 200.4775 2.745 ;
      RECT  40.6 45.005 40.8325 73.2125 ;
      RECT  40.4175 45.005 40.6 47.19 ;
      RECT  326.7325 2.33 337.7575 2.745 ;
      RECT  338.1725 2.33 349.1975 2.745 ;
      RECT  40.6 36.035 40.8325 41.6 ;
      RECT  40.6 42.015 40.8325 44.59 ;
      RECT  40.4175 36.035 40.6 41.6 ;
      RECT  40.4175 42.015 40.6 44.59 ;
      RECT  349.6125 2.33 360.6375 2.745 ;
      RECT  361.0525 2.33 372.0775 2.745 ;
      RECT  41.015 0.275 363.4975 0.965 ;
      RECT  363.4975 0.275 363.9125 0.965 ;
      RECT  363.9125 0.275 383.585 0.965 ;
      RECT  35.295 33.045 38.89 37.115 ;
      RECT  35.295 37.115 38.89 37.53 ;
      RECT  35.295 37.53 38.89 47.19 ;
      RECT  39.305 33.045 40.4175 37.115 ;
      RECT  39.305 37.115 40.4175 37.53 ;
      RECT  39.305 37.53 40.4175 47.19 ;
      RECT  38.89 37.53 39.305 40.105 ;
      RECT  35.295 2.745 38.89 31.135 ;
      RECT  35.295 31.135 38.89 31.55 ;
      RECT  35.295 31.55 38.89 32.63 ;
      RECT  38.89 2.745 39.305 31.135 ;
      RECT  38.89 31.55 39.305 32.63 ;
      RECT  39.305 2.745 40.3175 31.135 ;
      RECT  39.305 31.135 40.3175 31.55 ;
      RECT  39.305 31.55 40.3175 32.63 ;
      RECT  219.655 72.385 251.975 73.075 ;
      RECT  219.655 73.075 251.975 73.2125 ;
      RECT  251.975 72.385 252.39 73.075 ;
      RECT  252.39 72.385 254.115 73.075 ;
      RECT  252.39 73.075 254.115 73.2125 ;
      RECT  363.9125 0.14 374.9375 0.275 ;
      RECT  375.3525 0.14 383.585 0.275 ;
      RECT  55.0325 0.14 66.0575 0.275 ;
      RECT  306.7125 0.14 317.7375 0.275 ;
      RECT  295.2725 0.14 306.2975 0.275 ;
      RECT  0.56 1.38 2.285 10.465 ;
      RECT  0.56 10.465 2.285 10.88 ;
      RECT  0.56 10.88 2.285 11.57 ;
      RECT  2.285 1.38 2.7 10.465 ;
      RECT  2.285 10.88 2.7 11.57 ;
      RECT  2.7 1.38 34.88 10.465 ;
      RECT  2.7 10.465 34.88 10.88 ;
      RECT  2.7 10.88 34.88 11.57 ;
      RECT  53.3125 22.1825 166.1575 23.8825 ;
      RECT  53.3125 24.2325 166.1575 27.2675 ;
      RECT  166.1575 22.1825 166.5725 23.8825 ;
      RECT  166.1575 24.2325 166.5725 27.2675 ;
      RECT  166.5725 22.1825 197.4075 23.8825 ;
      RECT  166.5725 24.2325 197.4075 27.2675 ;
      RECT  213.9225 30.445 215.035 37.115 ;
      RECT  213.9225 37.115 215.035 37.53 ;
      RECT  213.9225 37.53 215.035 41.6 ;
      RECT  215.45 30.445 219.24 37.115 ;
      RECT  215.45 37.115 219.24 37.53 ;
      RECT  215.45 37.53 219.24 41.6 ;
      RECT  180.8725 0.14 191.8975 0.275 ;
      RECT  318.1525 0.14 329.1775 0.275 ;
      RECT  329.5925 0.14 340.6175 0.275 ;
      RECT  112.2325 0.14 123.2575 0.275 ;
      RECT  123.6725 0.14 134.6975 0.275 ;
      RECT  272.3925 0.14 283.4175 0.275 ;
      RECT  283.8325 0.14 294.8575 0.275 ;
      RECT  100.7925 0.14 111.8175 0.275 ;
      RECT  38.89 33.045 39.305 34.125 ;
      RECT  38.89 34.54 39.305 37.115 ;
      RECT  249.5125 0.14 260.5375 0.275 ;
      RECT  260.9525 0.14 271.9775 0.275 ;
      RECT  157.9925 0.14 169.0175 0.275 ;
      RECT  169.4325 0.14 180.4575 0.275 ;
      RECT  213.9225 42.015 215.035 43.095 ;
      RECT  213.9225 43.095 215.035 43.51 ;
      RECT  213.9225 43.51 215.035 65.2625 ;
      RECT  215.035 42.015 215.45 43.095 ;
      RECT  215.45 42.015 219.24 43.095 ;
      RECT  215.45 43.095 219.24 43.51 ;
      RECT  215.45 43.51 219.24 65.2625 ;
      RECT  38.89 46.5 39.305 47.19 ;
      RECT  89.3525 0.14 100.3775 0.275 ;
      RECT  215.035 37.53 215.45 40.105 ;
      RECT  215.035 40.52 215.45 41.6 ;
      RECT  56.4975 59.1575 56.9125 60.8125 ;
      RECT  56.4975 61.1625 56.9125 62.705 ;
      RECT  53.3125 59.1575 56.4975 60.8125 ;
      RECT  53.3125 61.1625 56.4975 62.705 ;
      RECT  56.9125 59.1575 197.4075 60.8125 ;
      RECT  56.9125 61.1625 197.4075 62.705 ;
      RECT  197.4075 59.1575 197.4425 60.8125 ;
      RECT  197.4075 61.1625 197.4425 62.705 ;
      RECT  197.4425 59.1575 199.0525 60.8125 ;
      RECT  197.4425 60.8125 199.0525 61.1625 ;
      RECT  197.4425 61.1625 199.0525 62.705 ;
      RECT  215.035 30.445 215.45 31.135 ;
      RECT  238.0725 0.14 249.0975 0.275 ;
      RECT  135.1125 0.14 146.1375 0.275 ;
      RECT  146.5525 0.14 157.5775 0.275 ;
      RECT  215.1925 0.14 226.2175 0.275 ;
      RECT  226.6325 0.14 237.6575 0.275 ;
      RECT  341.0325 0.14 352.0575 0.275 ;
      RECT  352.4725 0.14 363.4975 0.275 ;
      RECT  215.035 31.55 215.45 34.125 ;
      RECT  215.035 34.54 215.45 37.115 ;
      RECT  215.035 43.51 215.45 46.085 ;
      RECT  215.035 46.5 215.45 65.2625 ;
      RECT  41.015 0.14 43.1775 0.275 ;
      RECT  43.5925 0.14 54.6175 0.275 ;
      RECT  192.3125 0.14 203.3375 0.275 ;
      RECT  203.7525 0.14 214.7775 0.275 ;
      RECT  66.4725 0.14 77.4975 0.275 ;
      RECT  77.9125 0.14 88.9375 0.275 ;
      RECT  38.89 40.52 39.305 43.095 ;
      RECT  38.89 43.51 39.305 46.085 ;
   LAYER  metal4 ;
      RECT  0.14 58.5325 53.105 73.2125 ;
      RECT  53.105 0.14 53.805 27.8225 ;
      RECT  53.105 58.5325 53.805 73.2125 ;
      RECT  253.5675 27.8225 254.2675 40.8225 ;
      RECT  254.2675 27.8225 383.585 40.8225 ;
      RECT  254.2675 40.8225 383.585 58.5325 ;
      RECT  253.5675 63.785 254.2675 73.2125 ;
      RECT  254.2675 58.5325 383.585 63.785 ;
      RECT  254.2675 63.785 383.585 73.2125 ;
      RECT  0.14 0.14 0.4075 20.17 ;
      RECT  0.14 20.17 0.4075 27.8225 ;
      RECT  0.4075 0.14 1.1075 20.17 ;
      RECT  0.14 27.8225 0.4075 43.1325 ;
      RECT  0.14 43.1325 0.4075 58.5325 ;
      RECT  0.4075 43.1325 1.1075 58.5325 ;
      RECT  1.1075 45.9425 34.455 56.5225 ;
      RECT  1.1075 56.5225 34.455 58.5325 ;
      RECT  34.455 43.1325 35.155 45.9425 ;
      RECT  34.455 56.5225 35.155 58.5325 ;
      RECT  52.025 27.8225 52.725 30.9925 ;
      RECT  52.725 27.8225 53.105 30.9925 ;
      RECT  52.725 30.9925 53.105 43.1325 ;
      RECT  52.725 43.1325 53.105 45.9425 ;
      RECT  52.025 55.6125 52.725 56.5225 ;
      RECT  52.725 45.9425 53.105 55.6125 ;
      RECT  52.725 55.6125 53.105 56.5225 ;
      RECT  219.38 0.14 220.08 21.1125 ;
      RECT  220.08 0.14 383.585 21.1125 ;
      RECT  220.08 21.1125 383.585 27.8225 ;
      RECT  219.38 31.6925 220.08 40.8225 ;
      RECT  220.08 27.8225 253.5675 31.6925 ;
      RECT  44.925 55.6825 45.625 56.5225 ;
      RECT  45.625 55.6825 52.025 56.5225 ;
      RECT  53.805 58.5325 216.66 60.5825 ;
      RECT  53.805 60.5825 216.66 63.785 ;
      RECT  216.66 58.5325 217.36 60.5825 ;
      RECT  53.805 63.785 216.66 71.1625 ;
      RECT  53.805 71.1625 216.66 73.2125 ;
      RECT  216.66 71.1625 217.36 73.2125 ;
      RECT  201.235 55.6825 208.715 58.5325 ;
      RECT  208.715 55.6825 209.415 58.5325 ;
      RECT  201.235 40.8225 201.615 55.6125 ;
      RECT  201.235 55.6125 201.615 55.6825 ;
      RECT  201.615 55.6125 202.315 55.6825 ;
      RECT  201.235 30.9925 201.615 31.6925 ;
      RECT  201.235 31.6925 201.615 40.8225 ;
      RECT  37.175 0.14 37.875 12.7925 ;
      RECT  37.875 0.14 53.105 12.7925 ;
      RECT  37.875 12.7925 53.105 20.17 ;
      RECT  37.875 20.17 53.105 27.8225 ;
      RECT  37.175 28.3125 37.875 30.9925 ;
      RECT  37.875 27.8225 52.025 28.3125 ;
      RECT  1.1075 43.1325 2.47 43.165 ;
      RECT  1.1075 43.165 2.47 45.9425 ;
      RECT  2.47 43.165 3.17 45.9425 ;
      RECT  3.17 43.1325 34.455 43.165 ;
      RECT  3.17 43.165 34.455 45.9425 ;
      RECT  1.1075 30.9925 2.47 43.1325 ;
      RECT  1.1075 20.17 2.47 20.2025 ;
      RECT  1.1075 20.2025 2.47 27.8225 ;
      RECT  2.47 20.17 3.17 20.2025 ;
      RECT  1.1075 27.8225 2.47 28.3125 ;
      RECT  3.17 27.8225 37.175 28.3125 ;
      RECT  1.1075 28.3125 2.47 30.9925 ;
      RECT  3.17 28.3125 37.175 30.9925 ;
      RECT  1.1075 0.14 5.825 10.3225 ;
      RECT  1.1075 10.3225 5.825 12.7925 ;
      RECT  5.825 0.14 6.525 10.3225 ;
      RECT  6.525 0.14 37.175 10.3225 ;
      RECT  6.525 10.3225 37.175 12.7925 ;
      RECT  1.1075 12.7925 5.825 20.17 ;
      RECT  6.525 12.7925 37.175 20.17 ;
      RECT  3.17 20.17 5.825 20.2025 ;
      RECT  6.525 20.17 37.175 20.2025 ;
      RECT  3.17 20.2025 5.825 25.8425 ;
      RECT  3.17 25.8425 5.825 27.8225 ;
      RECT  5.825 25.8425 6.525 27.8225 ;
      RECT  6.525 20.2025 37.175 25.8425 ;
      RECT  6.525 25.8425 37.175 27.8225 ;
      RECT  217.36 58.5325 248.01 60.5825 ;
      RECT  217.36 60.5825 248.01 63.785 ;
      RECT  217.36 63.785 248.01 71.1625 ;
      RECT  248.71 63.785 253.5675 71.1625 ;
      RECT  217.36 71.1625 248.01 73.2125 ;
      RECT  248.71 71.1625 253.5675 73.2125 ;
      RECT  209.415 55.6825 248.01 58.1125 ;
      RECT  209.415 58.1125 248.01 58.5325 ;
      RECT  248.01 55.6825 248.71 58.1125 ;
      RECT  220.08 31.6925 251.505 40.79 ;
      RECT  220.08 40.79 251.505 40.8225 ;
      RECT  251.505 31.6925 252.205 40.79 ;
      RECT  252.205 31.6925 253.5675 40.79 ;
      RECT  252.205 40.79 253.5675 40.8225 ;
      RECT  252.205 40.8225 253.5675 55.6825 ;
      RECT  248.71 58.5325 251.505 60.5825 ;
      RECT  252.205 58.5325 253.5675 60.5825 ;
      RECT  248.71 60.5825 251.505 63.7525 ;
      RECT  248.71 63.7525 251.505 63.785 ;
      RECT  251.505 63.7525 252.205 63.785 ;
      RECT  252.205 60.5825 253.5675 63.7525 ;
      RECT  252.205 63.7525 253.5675 63.785 ;
      RECT  248.71 55.6825 251.505 58.1125 ;
      RECT  252.205 55.6825 253.5675 58.1125 ;
      RECT  248.71 58.1125 251.505 58.5325 ;
      RECT  252.205 58.1125 253.5675 58.5325 ;
      RECT  46.185 30.9925 52.025 43.1325 ;
      RECT  46.185 43.1325 52.025 45.9425 ;
      RECT  46.185 45.9425 52.025 55.6125 ;
      RECT  45.625 55.645 46.185 55.6825 ;
      RECT  46.185 55.6125 52.025 55.645 ;
      RECT  46.185 55.645 52.025 55.6825 ;
      RECT  37.875 28.3125 45.485 30.96 ;
      RECT  45.485 28.3125 46.185 30.96 ;
      RECT  46.185 28.3125 52.025 30.96 ;
      RECT  46.185 30.96 52.025 30.9925 ;
      RECT  35.155 56.5225 37.315 56.5875 ;
      RECT  35.155 56.5875 37.315 58.5325 ;
      RECT  37.315 56.5875 38.015 58.5325 ;
      RECT  38.015 56.5225 53.105 56.5875 ;
      RECT  38.015 56.5875 53.105 58.5325 ;
      RECT  35.155 43.1325 37.315 45.8775 ;
      RECT  35.155 45.8775 37.315 45.9425 ;
      RECT  37.315 43.1325 38.015 45.8775 ;
      RECT  35.155 45.9425 37.315 55.6125 ;
      RECT  35.155 55.6125 37.315 55.6825 ;
      RECT  35.155 55.6825 37.315 56.5225 ;
      RECT  38.015 55.6825 44.925 56.5225 ;
      RECT  53.805 0.14 216.52 21.0475 ;
      RECT  53.805 21.0475 216.52 21.1125 ;
      RECT  216.52 0.14 217.22 21.0475 ;
      RECT  217.22 0.14 219.38 21.0475 ;
      RECT  217.22 21.0475 219.38 21.1125 ;
      RECT  53.805 21.1125 216.52 27.8225 ;
      RECT  217.22 21.1125 219.38 27.8225 ;
      RECT  217.22 27.8225 219.38 30.9925 ;
      RECT  217.22 30.9925 219.38 31.6925 ;
      RECT  216.52 31.7575 217.22 40.8225 ;
      RECT  217.22 31.6925 219.38 31.7575 ;
      RECT  217.22 31.7575 219.38 40.8225 ;
      RECT  201.235 27.8225 208.155 30.96 ;
      RECT  201.235 30.96 208.155 30.9925 ;
      RECT  208.155 27.8225 208.715 30.96 ;
      RECT  208.715 27.8225 208.855 30.96 ;
      RECT  208.855 27.8225 209.415 30.96 ;
      RECT  208.855 30.96 209.415 30.9925 ;
      RECT  202.315 40.8225 208.155 55.6125 ;
      RECT  202.315 55.6125 208.155 55.645 ;
      RECT  202.315 55.645 208.155 55.6825 ;
      RECT  208.155 55.645 208.715 55.6825 ;
      RECT  202.315 30.9925 208.155 31.6925 ;
      RECT  202.315 31.6925 208.155 40.8225 ;
      RECT  54.265 27.8225 200.075 40.8225 ;
      RECT  54.265 40.8225 200.075 58.5325 ;
      RECT  3.17 30.9925 43.335 43.1325 ;
      RECT  44.035 30.9925 44.925 43.1325 ;
      RECT  37.875 30.96 43.335 30.9925 ;
      RECT  44.035 30.96 45.485 30.9925 ;
      RECT  38.015 43.1325 43.335 45.8775 ;
      RECT  44.035 43.1325 44.925 45.8775 ;
      RECT  38.015 45.8775 43.335 45.9425 ;
      RECT  44.035 45.8775 44.925 45.9425 ;
      RECT  38.015 45.9425 43.335 55.6125 ;
      RECT  44.035 45.9425 44.925 55.6125 ;
      RECT  38.015 55.6125 43.335 55.6825 ;
      RECT  44.035 55.6125 44.925 55.6825 ;
      RECT  209.415 40.8225 210.305 55.6825 ;
      RECT  211.005 40.8225 251.505 55.6825 ;
      RECT  209.415 27.8225 210.305 30.96 ;
      RECT  209.415 30.96 210.305 30.9925 ;
      RECT  210.305 27.8225 211.005 30.96 ;
      RECT  211.005 27.8225 216.52 30.96 ;
      RECT  211.005 30.96 216.52 30.9925 ;
      RECT  209.415 30.9925 210.305 31.6925 ;
      RECT  211.005 30.9925 216.52 31.6925 ;
      RECT  209.415 31.6925 210.305 31.7575 ;
      RECT  211.005 31.6925 216.52 31.7575 ;
      RECT  209.415 31.7575 210.305 40.8225 ;
      RECT  211.005 31.7575 216.52 40.8225 ;
   END
END    freepdk45_sram_1w1r_16x120
END    LIBRARY
