VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_1w1r_13x128
   CLASS BLOCK ;
   SIZE 126.005 BY 88.705 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  23.36 1.105 23.495 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  26.22 1.105 26.355 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.08 1.105 29.215 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.94 1.105 32.075 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.8 1.105 34.935 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.66 1.105 37.795 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.52 1.105 40.655 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.38 1.105 43.515 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.24 1.105 46.375 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.1 1.105 49.235 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.96 1.105 52.095 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.82 1.105 54.955 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.68 1.105 57.815 1.24 ;
      END
   END din0[12]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  17.64 1.105 17.775 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  20.5 1.105 20.635 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 43.37 12.055 43.505 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 46.1 12.055 46.235 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 48.31 12.055 48.445 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 51.04 12.055 51.175 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  11.92 53.25 12.055 53.385 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.23 87.465 105.365 87.6 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.37 87.465 102.505 87.6 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.81 20.23 113.945 20.365 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.81 17.5 113.945 17.635 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.81 15.29 113.945 15.425 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.81 12.56 113.945 12.695 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.81 10.35 113.945 10.485 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.77 0.42 1.905 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.585 86.09 125.72 86.225 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.855 6.3825 1.99 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.4825 86.005 119.6175 86.14 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.2525 82.5975 32.3875 82.7325 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.9525 82.5975 37.0875 82.7325 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.6525 82.5975 41.7875 82.7325 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.3525 82.5975 46.4875 82.7325 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.0525 82.5975 51.1875 82.7325 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.7525 82.5975 55.8875 82.7325 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.4525 82.5975 60.5875 82.7325 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.1525 82.5975 65.2875 82.7325 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.8525 82.5975 69.9875 82.7325 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.5525 82.5975 74.6875 82.7325 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.2525 82.5975 79.3875 82.7325 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.9525 82.5975 84.0875 82.7325 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.6525 82.5975 88.7875 82.7325 ;
      END
   END dout1[12]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  114.09 8.9175 114.23 21.4725 ;
         LAYER metal3 ;
         RECT  18.0175 34.79 18.1525 34.925 ;
         LAYER metal3 ;
         RECT  29.0675 17.4675 93.4525 17.5375 ;
         LAYER metal4 ;
         RECT  11.635 42.2625 11.775 54.8175 ;
         LAYER metal3 ;
         RECT  18.0175 37.78 18.1525 37.915 ;
         LAYER metal3 ;
         RECT  27.9225 19.84 28.0575 19.975 ;
         LAYER metal3 ;
         RECT  18.0175 31.8 18.1525 31.935 ;
         LAYER metal3 ;
         RECT  123.445 84.725 123.58 84.86 ;
         LAYER metal4 ;
         RECT  101.96 21.3325 102.1 69.3825 ;
         LAYER metal3 ;
         RECT  57.3975 2.47 57.5325 2.605 ;
         LAYER metal3 ;
         RECT  18.3625 25.82 18.4975 25.955 ;
         LAYER metal4 ;
         RECT  97.61 21.3325 97.75 69.3125 ;
         LAYER metal4 ;
         RECT  14.355 3.1325 14.495 18.0925 ;
         LAYER metal4 ;
         RECT  96.53 18.1625 96.67 72.2325 ;
         LAYER metal3 ;
         RECT  29.0675 80.04 89.4575 80.11 ;
         LAYER metal3 ;
         RECT  107.5175 34.79 107.6525 34.925 ;
         LAYER metal4 ;
         RECT  103.805 75.32 103.945 85.34 ;
         LAYER metal3 ;
         RECT  45.9575 2.47 46.0925 2.605 ;
         LAYER metal3 ;
         RECT  34.5175 2.47 34.6525 2.605 ;
         LAYER metal3 ;
         RECT  101.345 69.8825 101.48 70.0175 ;
         LAYER metal3 ;
         RECT  18.3625 22.83 18.4975 22.965 ;
         LAYER metal3 ;
         RECT  97.6125 70.67 97.7475 70.805 ;
         LAYER metal3 ;
         RECT  23.0775 2.47 23.2125 2.605 ;
         LAYER metal4 ;
         RECT  0.6875 10.51 0.8275 32.9125 ;
         LAYER metal4 ;
         RECT  23.57 21.3325 23.71 69.3825 ;
         LAYER metal4 ;
         RECT  125.1775 55.0825 125.3175 77.485 ;
         LAYER metal3 ;
         RECT  24.19 20.6275 24.325 20.7625 ;
         LAYER metal3 ;
         RECT  17.3575 2.47 17.4925 2.605 ;
         LAYER metal3 ;
         RECT  107.5175 31.8 107.6525 31.935 ;
         LAYER metal3 ;
         RECT  107.1725 25.82 107.3075 25.955 ;
         LAYER metal3 ;
         RECT  107.5175 37.78 107.6525 37.915 ;
         LAYER metal3 ;
         RECT  29.0675 72.9275 94.6275 72.9975 ;
         LAYER metal3 ;
         RECT  2.425 3.135 2.56 3.27 ;
         LAYER metal4 ;
         RECT  27.92 21.3325 28.06 69.3125 ;
         LAYER metal4 ;
         RECT  21.725 5.125 21.865 15.145 ;
         LAYER metal4 ;
         RECT  29.0 18.1625 29.14 72.2325 ;
         LAYER metal3 ;
         RECT  105.5125 86.1 105.6475 86.235 ;
         LAYER metal3 ;
         RECT  18.0175 40.77 18.1525 40.905 ;
         LAYER metal3 ;
         RECT  107.1725 22.83 107.3075 22.965 ;
         LAYER metal4 ;
         RECT  111.37 74.8425 111.51 84.8625 ;
         LAYER metal3 ;
         RECT  29.0675 8.8175 89.4575 8.8875 ;
         LAYER metal3 ;
         RECT  107.5175 40.77 107.6525 40.905 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  29.46 18.1625 29.6 72.2325 ;
         LAYER metal3 ;
         RECT  16.21 30.305 16.345 30.44 ;
         LAYER metal3 ;
         RECT  16.21 36.285 16.345 36.42 ;
         LAYER metal4 ;
         RECT  24.13 21.3 24.27 69.345 ;
         LAYER metal4 ;
         RECT  2.75 10.5425 2.89 32.945 ;
         LAYER metal3 ;
         RECT  108.7 21.335 108.835 21.47 ;
         LAYER metal4 ;
         RECT  14.495 42.1975 14.635 54.7525 ;
         LAYER metal3 ;
         RECT  123.445 87.195 123.58 87.33 ;
         LAYER metal3 ;
         RECT  16.21 42.265 16.345 42.4 ;
         LAYER metal3 ;
         RECT  29.0675 75.5475 93.485 75.6175 ;
         LAYER metal3 ;
         RECT  16.21 39.275 16.345 39.41 ;
         LAYER metal3 ;
         RECT  37.3775 0.0 37.5125 0.135 ;
         LAYER metal3 ;
         RECT  60.2575 0.0 60.3925 0.135 ;
         LAYER metal3 ;
         RECT  16.835 21.335 16.97 21.47 ;
         LAYER metal4 ;
         RECT  21.98 21.3 22.12 69.3825 ;
         LAYER metal4 ;
         RECT  6.105 0.6625 6.245 15.6225 ;
         LAYER metal4 ;
         RECT  103.55 21.3 103.69 69.3825 ;
         LAYER metal3 ;
         RECT  2.425 0.665 2.56 0.8 ;
         LAYER metal3 ;
         RECT  16.21 33.295 16.345 33.43 ;
         LAYER metal4 ;
         RECT  119.62 72.3725 119.76 87.3325 ;
         LAYER metal3 ;
         RECT  108.7 27.315 108.835 27.45 ;
         LAYER metal4 ;
         RECT  96.07 18.1625 96.21 72.2325 ;
         LAYER metal3 ;
         RECT  25.9375 0.0 26.0725 0.135 ;
         LAYER metal4 ;
         RECT  105.4675 75.2525 105.6075 85.4075 ;
         LAYER metal4 ;
         RECT  111.23 8.9825 111.37 21.5375 ;
         LAYER metal3 ;
         RECT  109.325 33.295 109.46 33.43 ;
         LAYER metal3 ;
         RECT  20.2175 0.0 20.3525 0.135 ;
         LAYER metal3 ;
         RECT  29.0675 78.1475 89.4925 78.2175 ;
         LAYER metal3 ;
         RECT  48.8175 0.0 48.9525 0.135 ;
         LAYER metal3 ;
         RECT  108.7 24.325 108.835 24.46 ;
         LAYER metal3 ;
         RECT  16.835 24.325 16.97 24.46 ;
         LAYER metal3 ;
         RECT  109.325 39.275 109.46 39.41 ;
         LAYER metal3 ;
         RECT  16.835 27.315 16.97 27.45 ;
         LAYER metal3 ;
         RECT  109.325 30.305 109.46 30.44 ;
         LAYER metal3 ;
         RECT  109.325 42.265 109.46 42.4 ;
         LAYER metal3 ;
         RECT  109.325 36.285 109.46 36.42 ;
         LAYER metal3 ;
         RECT  102.6525 88.57 102.7875 88.705 ;
         LAYER metal3 ;
         RECT  29.0675 14.8475 93.485 14.9175 ;
         LAYER metal3 ;
         RECT  29.0675 10.8675 89.4575 10.9375 ;
         LAYER metal4 ;
         RECT  20.0625 5.0575 20.2025 15.2125 ;
         LAYER metal4 ;
         RECT  123.115 55.05 123.255 77.4525 ;
         LAYER metal4 ;
         RECT  101.4 21.3 101.54 69.345 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 125.865 88.565 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 125.865 88.565 ;
   LAYER  metal3 ;
      RECT  23.22 0.14 23.635 0.965 ;
      RECT  23.635 0.965 26.08 1.38 ;
      RECT  26.495 0.965 28.94 1.38 ;
      RECT  29.355 0.965 31.8 1.38 ;
      RECT  32.215 0.965 34.66 1.38 ;
      RECT  35.075 0.965 37.52 1.38 ;
      RECT  37.935 0.965 40.38 1.38 ;
      RECT  40.795 0.965 43.24 1.38 ;
      RECT  43.655 0.965 46.1 1.38 ;
      RECT  46.515 0.965 48.96 1.38 ;
      RECT  49.375 0.965 51.82 1.38 ;
      RECT  52.235 0.965 54.68 1.38 ;
      RECT  55.095 0.965 57.54 1.38 ;
      RECT  57.955 0.965 125.865 1.38 ;
      RECT  0.14 0.965 17.5 1.38 ;
      RECT  17.915 0.965 20.36 1.38 ;
      RECT  20.775 0.965 23.22 1.38 ;
      RECT  0.14 43.23 11.78 43.645 ;
      RECT  0.14 43.645 11.78 88.565 ;
      RECT  11.78 1.38 12.195 43.23 ;
      RECT  12.195 43.23 23.22 43.645 ;
      RECT  12.195 43.645 23.22 88.565 ;
      RECT  11.78 43.645 12.195 45.96 ;
      RECT  11.78 46.375 12.195 48.17 ;
      RECT  11.78 48.585 12.195 50.9 ;
      RECT  11.78 51.315 12.195 53.11 ;
      RECT  11.78 53.525 12.195 88.565 ;
      RECT  105.09 87.74 105.505 88.565 ;
      RECT  105.505 87.74 125.865 88.565 ;
      RECT  23.635 87.325 102.23 87.74 ;
      RECT  102.645 87.325 105.09 87.74 ;
      RECT  105.505 1.38 113.67 20.09 ;
      RECT  105.505 20.09 113.67 20.505 ;
      RECT  113.67 20.505 114.085 87.325 ;
      RECT  114.085 1.38 125.865 20.09 ;
      RECT  114.085 20.09 125.865 20.505 ;
      RECT  113.67 17.775 114.085 20.09 ;
      RECT  113.67 15.565 114.085 17.36 ;
      RECT  113.67 12.835 114.085 15.15 ;
      RECT  113.67 1.38 114.085 10.21 ;
      RECT  113.67 10.625 114.085 12.42 ;
      RECT  0.14 1.38 0.145 1.63 ;
      RECT  0.14 1.63 0.145 2.045 ;
      RECT  0.14 2.045 0.145 43.23 ;
      RECT  0.145 1.38 0.56 1.63 ;
      RECT  0.145 2.045 0.56 43.23 ;
      RECT  0.56 1.38 11.78 1.63 ;
      RECT  125.445 20.505 125.86 85.95 ;
      RECT  125.445 86.365 125.86 87.325 ;
      RECT  125.86 20.505 125.865 85.95 ;
      RECT  125.86 85.95 125.865 86.365 ;
      RECT  125.86 86.365 125.865 87.325 ;
      RECT  0.56 1.63 6.1075 1.715 ;
      RECT  0.56 1.715 6.1075 2.045 ;
      RECT  6.1075 1.63 6.5225 1.715 ;
      RECT  6.5225 1.63 11.78 1.715 ;
      RECT  6.5225 1.715 11.78 2.045 ;
      RECT  0.56 2.045 6.1075 2.13 ;
      RECT  6.1075 2.13 6.5225 43.23 ;
      RECT  6.5225 2.045 11.78 2.13 ;
      RECT  6.5225 2.13 11.78 43.23 ;
      RECT  114.085 20.505 119.3425 85.865 ;
      RECT  114.085 85.865 119.3425 85.95 ;
      RECT  119.3425 20.505 119.7575 85.865 ;
      RECT  119.7575 85.865 125.445 85.95 ;
      RECT  114.085 85.95 119.3425 86.28 ;
      RECT  114.085 86.28 119.3425 86.365 ;
      RECT  119.3425 86.28 119.7575 86.365 ;
      RECT  119.7575 85.95 125.445 86.28 ;
      RECT  119.7575 86.28 125.445 86.365 ;
      RECT  23.635 82.4575 32.1125 82.8725 ;
      RECT  23.635 82.8725 32.1125 87.325 ;
      RECT  32.1125 82.8725 32.5275 87.325 ;
      RECT  32.5275 82.8725 105.09 87.325 ;
      RECT  32.5275 82.4575 36.8125 82.8725 ;
      RECT  37.2275 82.4575 41.5125 82.8725 ;
      RECT  41.9275 82.4575 46.2125 82.8725 ;
      RECT  46.6275 82.4575 50.9125 82.8725 ;
      RECT  51.3275 82.4575 55.6125 82.8725 ;
      RECT  56.0275 82.4575 60.3125 82.8725 ;
      RECT  60.7275 82.4575 65.0125 82.8725 ;
      RECT  65.4275 82.4575 69.7125 82.8725 ;
      RECT  70.1275 82.4575 74.4125 82.8725 ;
      RECT  74.8275 82.4575 79.1125 82.8725 ;
      RECT  79.5275 82.4575 83.8125 82.8725 ;
      RECT  84.2275 82.4575 88.5125 82.8725 ;
      RECT  88.9275 82.4575 105.09 82.8725 ;
      RECT  12.195 34.65 17.8775 35.065 ;
      RECT  18.2925 34.65 23.22 35.065 ;
      RECT  18.2925 35.065 23.22 43.23 ;
      RECT  23.635 1.38 28.9275 17.3275 ;
      RECT  23.635 17.3275 28.9275 17.6775 ;
      RECT  93.5925 17.3275 105.09 17.6775 ;
      RECT  17.8775 35.065 18.2925 37.64 ;
      RECT  23.635 17.6775 27.7825 19.7 ;
      RECT  23.635 19.7 27.7825 20.115 ;
      RECT  27.7825 17.6775 28.1975 19.7 ;
      RECT  27.7825 20.115 28.1975 82.4575 ;
      RECT  28.1975 17.6775 28.9275 19.7 ;
      RECT  28.1975 19.7 28.9275 20.115 ;
      RECT  28.1975 20.115 28.9275 82.4575 ;
      RECT  17.8775 32.075 18.2925 34.65 ;
      RECT  119.7575 20.505 123.305 84.585 ;
      RECT  119.7575 84.585 123.305 85.0 ;
      RECT  119.7575 85.0 123.305 85.865 ;
      RECT  123.305 20.505 123.72 84.585 ;
      RECT  123.305 85.0 123.72 85.865 ;
      RECT  123.72 20.505 125.445 84.585 ;
      RECT  123.72 84.585 125.445 85.0 ;
      RECT  123.72 85.0 125.445 85.865 ;
      RECT  32.5275 1.38 57.2575 2.33 ;
      RECT  57.2575 1.38 57.6725 2.33 ;
      RECT  57.6725 1.38 93.5925 2.33 ;
      RECT  57.6725 2.33 93.5925 2.745 ;
      RECT  18.2925 26.095 18.6375 34.65 ;
      RECT  18.6375 25.68 23.22 26.095 ;
      RECT  18.6375 26.095 23.22 34.65 ;
      RECT  17.8775 1.38 18.2225 25.68 ;
      RECT  17.8775 25.68 18.2225 26.095 ;
      RECT  17.8775 26.095 18.2225 31.66 ;
      RECT  18.2225 26.095 18.2925 31.66 ;
      RECT  28.9275 80.25 32.1125 82.4575 ;
      RECT  32.1125 80.25 32.5275 82.4575 ;
      RECT  32.5275 80.25 89.5975 82.4575 ;
      RECT  89.5975 79.9 93.5925 80.25 ;
      RECT  89.5975 80.25 93.5925 82.4575 ;
      RECT  105.505 34.65 107.3775 35.065 ;
      RECT  107.7925 34.65 113.67 35.065 ;
      RECT  46.2325 2.33 57.2575 2.745 ;
      RECT  32.5275 2.33 34.3775 2.745 ;
      RECT  34.7925 2.33 45.8175 2.745 ;
      RECT  93.5925 17.6775 101.205 69.7425 ;
      RECT  93.5925 69.7425 101.205 70.1575 ;
      RECT  101.205 17.6775 101.62 69.7425 ;
      RECT  101.205 70.1575 101.62 82.4575 ;
      RECT  101.62 17.6775 105.09 69.7425 ;
      RECT  101.62 69.7425 105.09 70.1575 ;
      RECT  101.62 70.1575 105.09 82.4575 ;
      RECT  18.2925 1.38 18.6375 22.69 ;
      RECT  18.2925 23.105 18.6375 25.68 ;
      RECT  18.2225 1.38 18.2925 22.69 ;
      RECT  18.2225 23.105 18.2925 25.68 ;
      RECT  93.5925 70.1575 97.4725 70.53 ;
      RECT  93.5925 70.53 97.4725 70.945 ;
      RECT  97.4725 70.1575 97.8875 70.53 ;
      RECT  97.4725 70.945 97.8875 82.4575 ;
      RECT  97.8875 70.1575 101.205 70.53 ;
      RECT  97.8875 70.53 101.205 70.945 ;
      RECT  97.8875 70.945 101.205 82.4575 ;
      RECT  23.22 1.38 23.3525 2.33 ;
      RECT  23.22 2.745 23.3525 88.565 ;
      RECT  23.3525 1.38 23.635 2.33 ;
      RECT  23.3525 2.33 23.635 2.745 ;
      RECT  23.3525 2.745 23.635 88.565 ;
      RECT  18.6375 1.38 22.9375 2.33 ;
      RECT  18.6375 2.33 22.9375 2.745 ;
      RECT  18.6375 2.745 22.9375 25.68 ;
      RECT  22.9375 1.38 23.22 2.33 ;
      RECT  22.9375 2.745 23.22 25.68 ;
      RECT  23.635 20.115 24.05 20.4875 ;
      RECT  23.635 20.4875 24.05 20.9025 ;
      RECT  23.635 20.9025 24.05 82.4575 ;
      RECT  24.05 20.115 24.465 20.4875 ;
      RECT  24.05 20.9025 24.465 82.4575 ;
      RECT  24.465 20.115 27.7825 20.4875 ;
      RECT  24.465 20.4875 27.7825 20.9025 ;
      RECT  24.465 20.9025 27.7825 82.4575 ;
      RECT  12.195 1.38 17.2175 2.33 ;
      RECT  12.195 2.33 17.2175 2.745 ;
      RECT  17.2175 1.38 17.6325 2.33 ;
      RECT  17.2175 2.745 17.6325 34.65 ;
      RECT  17.6325 1.38 17.8775 2.33 ;
      RECT  17.6325 2.33 17.8775 2.745 ;
      RECT  17.6325 2.745 17.8775 34.65 ;
      RECT  107.3775 32.075 107.7925 34.65 ;
      RECT  105.505 20.505 107.0325 25.68 ;
      RECT  105.505 25.68 107.0325 26.095 ;
      RECT  105.505 26.095 107.0325 34.65 ;
      RECT  107.0325 26.095 107.3775 34.65 ;
      RECT  107.3775 26.095 107.4475 31.66 ;
      RECT  107.4475 20.505 107.7925 25.68 ;
      RECT  107.4475 25.68 107.7925 26.095 ;
      RECT  107.4475 26.095 107.7925 31.66 ;
      RECT  107.3775 35.065 107.7925 37.64 ;
      RECT  28.9275 17.6775 32.1125 72.7875 ;
      RECT  32.1125 17.6775 32.5275 72.7875 ;
      RECT  32.5275 17.6775 89.5975 72.7875 ;
      RECT  89.5975 17.6775 93.5925 72.7875 ;
      RECT  93.5925 70.945 94.7675 72.7875 ;
      RECT  94.7675 70.945 97.4725 72.7875 ;
      RECT  94.7675 72.7875 97.4725 73.1375 ;
      RECT  94.7675 73.1375 97.4725 82.4575 ;
      RECT  0.56 2.13 2.285 2.995 ;
      RECT  0.56 2.995 2.285 3.41 ;
      RECT  0.56 3.41 2.285 43.23 ;
      RECT  2.285 2.13 2.7 2.995 ;
      RECT  2.285 3.41 2.7 43.23 ;
      RECT  2.7 2.13 6.1075 2.995 ;
      RECT  2.7 2.995 6.1075 3.41 ;
      RECT  2.7 3.41 6.1075 43.23 ;
      RECT  105.09 1.38 105.3725 85.96 ;
      RECT  105.09 85.96 105.3725 86.375 ;
      RECT  105.09 86.375 105.3725 87.325 ;
      RECT  105.3725 1.38 105.505 85.96 ;
      RECT  105.3725 86.375 105.505 87.325 ;
      RECT  105.505 35.065 105.7875 85.96 ;
      RECT  105.505 86.375 105.7875 87.325 ;
      RECT  105.7875 35.065 107.3775 85.96 ;
      RECT  105.7875 85.96 107.3775 86.375 ;
      RECT  105.7875 86.375 107.3775 87.325 ;
      RECT  17.8775 38.055 18.2925 40.63 ;
      RECT  17.8775 41.045 18.2925 43.23 ;
      RECT  107.0325 20.505 107.3775 22.69 ;
      RECT  107.0325 23.105 107.3775 25.68 ;
      RECT  107.3775 20.505 107.4475 22.69 ;
      RECT  107.3775 23.105 107.4475 25.68 ;
      RECT  28.9275 1.38 32.1125 8.6775 ;
      RECT  32.1125 1.38 32.5275 8.6775 ;
      RECT  32.5275 2.745 57.2575 8.6775 ;
      RECT  57.2575 2.745 57.6725 8.6775 ;
      RECT  57.6725 2.745 89.5975 8.6775 ;
      RECT  89.5975 2.745 93.5925 8.6775 ;
      RECT  89.5975 8.6775 93.5925 9.0275 ;
      RECT  107.3775 38.055 107.7925 40.63 ;
      RECT  107.3775 41.045 107.7925 87.325 ;
      RECT  12.195 2.745 16.07 30.165 ;
      RECT  12.195 30.165 16.07 30.58 ;
      RECT  12.195 30.58 16.07 34.65 ;
      RECT  16.07 2.745 16.485 30.165 ;
      RECT  16.485 30.165 17.2175 30.58 ;
      RECT  16.485 30.58 17.2175 34.65 ;
      RECT  12.195 35.065 16.07 36.145 ;
      RECT  12.195 36.145 16.07 36.56 ;
      RECT  12.195 36.56 16.07 43.23 ;
      RECT  16.07 35.065 16.485 36.145 ;
      RECT  16.485 35.065 17.8775 36.145 ;
      RECT  16.485 36.145 17.8775 36.56 ;
      RECT  16.485 36.56 17.8775 43.23 ;
      RECT  107.7925 20.505 108.56 21.195 ;
      RECT  107.7925 21.195 108.56 21.61 ;
      RECT  107.7925 21.61 108.56 34.65 ;
      RECT  108.56 20.505 108.975 21.195 ;
      RECT  108.975 20.505 113.67 21.195 ;
      RECT  108.975 21.195 113.67 21.61 ;
      RECT  105.505 87.325 123.305 87.47 ;
      RECT  105.505 87.47 123.305 87.74 ;
      RECT  123.305 87.47 123.72 87.74 ;
      RECT  123.72 87.325 125.865 87.47 ;
      RECT  123.72 87.47 125.865 87.74 ;
      RECT  114.085 86.365 123.305 87.055 ;
      RECT  114.085 87.055 123.305 87.325 ;
      RECT  123.305 86.365 123.72 87.055 ;
      RECT  123.72 86.365 125.445 87.055 ;
      RECT  123.72 87.055 125.445 87.325 ;
      RECT  16.07 42.54 16.485 43.23 ;
      RECT  28.9275 73.1375 32.1125 75.4075 ;
      RECT  32.1125 73.1375 32.5275 75.4075 ;
      RECT  32.5275 73.1375 89.5975 75.4075 ;
      RECT  89.5975 73.1375 93.5925 75.4075 ;
      RECT  93.5925 73.1375 93.625 75.4075 ;
      RECT  93.5925 75.7575 93.625 82.4575 ;
      RECT  93.625 73.1375 94.7675 75.4075 ;
      RECT  93.625 75.4075 94.7675 75.7575 ;
      RECT  93.625 75.7575 94.7675 82.4575 ;
      RECT  16.07 36.56 16.485 39.135 ;
      RECT  16.07 39.55 16.485 42.125 ;
      RECT  23.635 0.275 37.2375 0.965 ;
      RECT  37.2375 0.275 37.6525 0.965 ;
      RECT  37.6525 0.275 125.865 0.965 ;
      RECT  60.5325 0.14 125.865 0.275 ;
      RECT  16.485 2.745 16.695 21.195 ;
      RECT  16.485 21.195 16.695 21.61 ;
      RECT  16.485 21.61 16.695 30.165 ;
      RECT  16.695 2.745 17.11 21.195 ;
      RECT  17.11 2.745 17.2175 21.195 ;
      RECT  17.11 21.195 17.2175 21.61 ;
      RECT  17.11 21.61 17.2175 30.165 ;
      RECT  0.14 0.14 2.285 0.525 ;
      RECT  0.14 0.525 2.285 0.94 ;
      RECT  0.14 0.94 2.285 0.965 ;
      RECT  2.285 0.14 2.7 0.525 ;
      RECT  2.285 0.94 2.7 0.965 ;
      RECT  2.7 0.525 23.22 0.94 ;
      RECT  2.7 0.94 23.22 0.965 ;
      RECT  16.07 30.58 16.485 33.155 ;
      RECT  16.07 33.57 16.485 34.65 ;
      RECT  108.56 27.59 108.975 34.65 ;
      RECT  23.635 0.14 25.7975 0.275 ;
      RECT  26.2125 0.14 37.2375 0.275 ;
      RECT  108.975 21.61 109.185 33.155 ;
      RECT  108.975 33.155 109.185 33.57 ;
      RECT  108.975 33.57 109.185 34.65 ;
      RECT  109.185 33.57 109.6 34.65 ;
      RECT  109.6 21.61 113.67 33.155 ;
      RECT  109.6 33.155 113.67 33.57 ;
      RECT  109.6 33.57 113.67 34.65 ;
      RECT  2.7 0.14 20.0775 0.275 ;
      RECT  2.7 0.275 20.0775 0.525 ;
      RECT  20.0775 0.275 20.4925 0.525 ;
      RECT  20.4925 0.14 23.22 0.275 ;
      RECT  20.4925 0.275 23.22 0.525 ;
      RECT  28.9275 75.7575 32.1125 78.0075 ;
      RECT  28.9275 78.3575 32.1125 79.9 ;
      RECT  32.1125 75.7575 32.5275 78.0075 ;
      RECT  32.1125 78.3575 32.5275 79.9 ;
      RECT  32.5275 75.7575 89.5975 78.0075 ;
      RECT  32.5275 78.3575 89.5975 79.9 ;
      RECT  89.5975 75.7575 89.6325 78.0075 ;
      RECT  89.5975 78.3575 89.6325 79.9 ;
      RECT  89.6325 75.7575 93.5925 78.0075 ;
      RECT  89.6325 78.0075 93.5925 78.3575 ;
      RECT  89.6325 78.3575 93.5925 79.9 ;
      RECT  37.6525 0.14 48.6775 0.275 ;
      RECT  49.0925 0.14 60.1175 0.275 ;
      RECT  108.56 21.61 108.975 24.185 ;
      RECT  108.56 24.6 108.975 27.175 ;
      RECT  16.695 21.61 17.11 24.185 ;
      RECT  107.7925 35.065 109.185 39.135 ;
      RECT  107.7925 39.135 109.185 39.55 ;
      RECT  107.7925 39.55 109.185 87.325 ;
      RECT  109.6 35.065 113.67 39.135 ;
      RECT  109.6 39.135 113.67 39.55 ;
      RECT  109.6 39.55 113.67 87.325 ;
      RECT  16.695 24.6 17.11 27.175 ;
      RECT  16.695 27.59 17.11 30.165 ;
      RECT  109.185 21.61 109.6 30.165 ;
      RECT  109.185 30.58 109.6 33.155 ;
      RECT  109.185 39.55 109.6 42.125 ;
      RECT  109.185 42.54 109.6 87.325 ;
      RECT  109.185 35.065 109.6 36.145 ;
      RECT  109.185 36.56 109.6 39.135 ;
      RECT  23.635 87.74 102.5125 88.43 ;
      RECT  23.635 88.43 102.5125 88.565 ;
      RECT  102.5125 87.74 102.9275 88.43 ;
      RECT  102.9275 87.74 105.09 88.43 ;
      RECT  102.9275 88.43 105.09 88.565 ;
      RECT  93.5925 1.38 93.625 14.7075 ;
      RECT  93.5925 15.0575 93.625 17.3275 ;
      RECT  93.625 1.38 105.09 14.7075 ;
      RECT  93.625 14.7075 105.09 15.0575 ;
      RECT  93.625 15.0575 105.09 17.3275 ;
      RECT  28.9275 15.0575 32.1125 17.3275 ;
      RECT  32.1125 15.0575 32.5275 17.3275 ;
      RECT  32.5275 15.0575 57.2575 17.3275 ;
      RECT  57.2575 15.0575 57.6725 17.3275 ;
      RECT  57.6725 15.0575 89.5975 17.3275 ;
      RECT  89.5975 9.0275 93.5925 14.7075 ;
      RECT  89.5975 15.0575 93.5925 17.3275 ;
      RECT  28.9275 9.0275 32.1125 10.7275 ;
      RECT  28.9275 11.0775 32.1125 14.7075 ;
      RECT  32.1125 9.0275 32.5275 10.7275 ;
      RECT  32.1125 11.0775 32.5275 14.7075 ;
      RECT  32.5275 9.0275 57.2575 10.7275 ;
      RECT  32.5275 11.0775 57.2575 14.7075 ;
      RECT  57.2575 9.0275 57.6725 10.7275 ;
      RECT  57.2575 11.0775 57.6725 14.7075 ;
      RECT  57.6725 9.0275 89.5975 10.7275 ;
      RECT  57.6725 11.0775 89.5975 14.7075 ;
   LAYER  metal4 ;
      RECT  113.81 0.14 114.51 8.6375 ;
      RECT  113.81 21.7525 114.51 88.565 ;
      RECT  114.51 0.14 125.865 8.6375 ;
      RECT  114.51 8.6375 125.865 21.7525 ;
      RECT  0.14 41.9825 11.355 55.0975 ;
      RECT  0.14 55.0975 11.355 88.565 ;
      RECT  11.355 21.7525 12.055 41.9825 ;
      RECT  11.355 55.0975 12.055 88.565 ;
      RECT  101.68 69.6625 102.38 88.565 ;
      RECT  97.33 69.5925 98.03 69.6625 ;
      RECT  14.075 0.14 14.775 2.8525 ;
      RECT  14.775 0.14 113.81 2.8525 ;
      RECT  14.075 18.3725 14.775 21.0525 ;
      RECT  12.055 72.5125 96.25 88.565 ;
      RECT  96.25 72.5125 96.95 88.565 ;
      RECT  96.95 69.6625 101.68 72.5125 ;
      RECT  96.95 72.5125 101.68 88.565 ;
      RECT  96.95 21.0525 97.33 21.7525 ;
      RECT  96.95 21.7525 97.33 41.9825 ;
      RECT  96.95 41.9825 97.33 55.0975 ;
      RECT  96.95 55.0975 97.33 69.5925 ;
      RECT  96.95 69.5925 97.33 69.6625 ;
      RECT  96.25 8.6375 96.95 17.8825 ;
      RECT  96.95 8.6375 101.68 17.8825 ;
      RECT  96.95 17.8825 101.68 18.3725 ;
      RECT  102.38 69.6625 103.525 75.04 ;
      RECT  102.38 75.04 103.525 85.62 ;
      RECT  102.38 85.62 103.525 88.565 ;
      RECT  103.525 69.6625 104.225 75.04 ;
      RECT  103.525 85.62 104.225 88.565 ;
      RECT  0.14 21.7525 0.4075 33.1925 ;
      RECT  0.14 33.1925 0.4075 41.9825 ;
      RECT  0.4075 33.1925 1.1075 41.9825 ;
      RECT  0.14 8.6375 0.4075 10.23 ;
      RECT  0.14 10.23 0.4075 18.3725 ;
      RECT  0.4075 8.6375 1.1075 10.23 ;
      RECT  0.14 18.3725 0.4075 21.0525 ;
      RECT  0.14 21.0525 0.4075 21.7525 ;
      RECT  124.8975 21.7525 125.5975 54.8025 ;
      RECT  124.8975 77.765 125.5975 88.565 ;
      RECT  125.5975 21.7525 125.865 54.8025 ;
      RECT  125.5975 54.8025 125.865 77.765 ;
      RECT  125.5975 77.765 125.865 88.565 ;
      RECT  21.445 2.8525 22.145 4.845 ;
      RECT  22.145 2.8525 113.81 4.845 ;
      RECT  22.145 4.845 113.81 8.6375 ;
      RECT  21.445 15.425 22.145 17.8825 ;
      RECT  22.145 8.6375 96.25 15.425 ;
      RECT  22.145 15.425 96.25 17.8825 ;
      RECT  12.055 69.6625 28.72 72.5125 ;
      RECT  14.775 17.8825 28.72 18.3725 ;
      RECT  28.34 21.7525 28.72 41.9825 ;
      RECT  28.34 41.9825 28.72 55.0975 ;
      RECT  28.34 55.0975 28.72 69.5925 ;
      RECT  28.34 21.0525 28.72 21.7525 ;
      RECT  104.225 69.6625 111.09 74.5625 ;
      RECT  111.09 69.6625 111.79 74.5625 ;
      RECT  111.79 69.6625 113.81 74.5625 ;
      RECT  111.79 74.5625 113.81 75.04 ;
      RECT  111.09 85.1425 111.79 85.62 ;
      RECT  111.79 75.04 113.81 85.1425 ;
      RECT  111.79 85.1425 113.81 85.62 ;
      RECT  24.55 21.7525 27.64 41.9825 ;
      RECT  24.55 41.9825 27.64 55.0975 ;
      RECT  24.55 55.0975 27.64 69.5925 ;
      RECT  24.55 21.0525 27.64 21.7525 ;
      RECT  14.775 18.3725 23.85 21.02 ;
      RECT  23.85 18.3725 24.55 21.02 ;
      RECT  24.55 18.3725 28.72 21.02 ;
      RECT  24.55 21.02 28.72 21.0525 ;
      RECT  23.99 69.625 24.55 69.6625 ;
      RECT  24.55 69.5925 28.72 69.625 ;
      RECT  24.55 69.625 28.72 69.6625 ;
      RECT  1.1075 21.7525 2.47 33.1925 ;
      RECT  3.17 21.7525 11.355 33.1925 ;
      RECT  1.1075 33.1925 2.47 33.225 ;
      RECT  1.1075 33.225 2.47 41.9825 ;
      RECT  2.47 33.225 3.17 41.9825 ;
      RECT  3.17 33.1925 11.355 33.225 ;
      RECT  3.17 33.225 11.355 41.9825 ;
      RECT  1.1075 10.23 2.47 10.2625 ;
      RECT  1.1075 10.2625 2.47 18.3725 ;
      RECT  2.47 10.23 3.17 10.2625 ;
      RECT  1.1075 18.3725 2.47 21.0525 ;
      RECT  3.17 18.3725 14.075 21.0525 ;
      RECT  1.1075 21.0525 2.47 21.7525 ;
      RECT  12.055 21.7525 14.215 41.9175 ;
      RECT  12.055 41.9175 14.215 41.9825 ;
      RECT  14.215 21.7525 14.915 41.9175 ;
      RECT  12.055 41.9825 14.215 55.0325 ;
      RECT  12.055 55.0325 14.215 55.0975 ;
      RECT  14.215 55.0325 14.915 55.0975 ;
      RECT  12.055 55.0975 21.7 69.5925 ;
      RECT  22.4 55.0975 23.29 69.5925 ;
      RECT  12.055 69.5925 21.7 69.6625 ;
      RECT  22.4 69.5925 23.29 69.6625 ;
      RECT  14.775 21.02 21.7 21.0525 ;
      RECT  22.4 21.02 23.85 21.0525 ;
      RECT  3.17 21.0525 21.7 21.7525 ;
      RECT  22.4 21.0525 23.29 21.7525 ;
      RECT  14.915 21.7525 21.7 41.9175 ;
      RECT  22.4 21.7525 23.29 41.9175 ;
      RECT  14.915 41.9175 21.7 41.9825 ;
      RECT  22.4 41.9175 23.29 41.9825 ;
      RECT  14.915 41.9825 21.7 55.0325 ;
      RECT  22.4 41.9825 23.29 55.0325 ;
      RECT  14.915 55.0325 21.7 55.0975 ;
      RECT  22.4 55.0325 23.29 55.0975 ;
      RECT  0.14 0.14 5.825 0.3825 ;
      RECT  0.14 0.3825 5.825 2.8525 ;
      RECT  5.825 0.14 6.525 0.3825 ;
      RECT  6.525 0.14 14.075 0.3825 ;
      RECT  6.525 0.3825 14.075 2.8525 ;
      RECT  0.14 2.8525 5.825 8.6375 ;
      RECT  6.525 2.8525 14.075 8.6375 ;
      RECT  1.1075 8.6375 5.825 10.23 ;
      RECT  6.525 8.6375 14.075 10.23 ;
      RECT  3.17 10.23 5.825 10.2625 ;
      RECT  6.525 10.23 14.075 10.2625 ;
      RECT  3.17 10.2625 5.825 15.9025 ;
      RECT  3.17 15.9025 5.825 18.3725 ;
      RECT  5.825 15.9025 6.525 18.3725 ;
      RECT  6.525 10.2625 14.075 15.9025 ;
      RECT  6.525 15.9025 14.075 18.3725 ;
      RECT  102.38 8.6375 103.27 21.02 ;
      RECT  102.38 21.02 103.27 21.0525 ;
      RECT  103.27 8.6375 103.97 21.02 ;
      RECT  102.38 21.0525 103.27 21.7525 ;
      RECT  102.38 21.7525 103.27 41.9825 ;
      RECT  102.38 41.9825 103.27 55.0975 ;
      RECT  103.97 41.9825 113.81 55.0975 ;
      RECT  102.38 55.0975 103.27 69.6625 ;
      RECT  103.97 55.0975 113.81 69.6625 ;
      RECT  114.51 54.8025 119.34 72.0925 ;
      RECT  114.51 72.0925 119.34 77.765 ;
      RECT  119.34 54.8025 120.04 72.0925 ;
      RECT  114.51 77.765 119.34 87.6125 ;
      RECT  114.51 87.6125 119.34 88.565 ;
      RECT  119.34 87.6125 120.04 88.565 ;
      RECT  120.04 77.765 124.8975 87.6125 ;
      RECT  120.04 87.6125 124.8975 88.565 ;
      RECT  29.88 69.6625 95.79 72.5125 ;
      RECT  29.88 17.8825 95.79 18.3725 ;
      RECT  29.88 18.3725 95.79 21.0525 ;
      RECT  29.88 69.5925 95.79 69.6625 ;
      RECT  29.88 21.7525 95.79 41.9825 ;
      RECT  29.88 41.9825 95.79 55.0975 ;
      RECT  29.88 55.0975 95.79 69.5925 ;
      RECT  29.88 21.0525 95.79 21.7525 ;
      RECT  104.225 85.62 105.1875 85.6875 ;
      RECT  104.225 85.6875 105.1875 88.565 ;
      RECT  105.1875 85.6875 105.8875 88.565 ;
      RECT  105.8875 85.62 113.81 85.6875 ;
      RECT  105.8875 85.6875 113.81 88.565 ;
      RECT  104.225 74.5625 105.1875 74.9725 ;
      RECT  104.225 74.9725 105.1875 75.04 ;
      RECT  105.1875 74.5625 105.8875 74.9725 ;
      RECT  105.8875 74.5625 111.09 74.9725 ;
      RECT  105.8875 74.9725 111.09 75.04 ;
      RECT  104.225 75.04 105.1875 85.1425 ;
      RECT  105.8875 75.04 111.09 85.1425 ;
      RECT  104.225 85.1425 105.1875 85.62 ;
      RECT  105.8875 85.1425 111.09 85.62 ;
      RECT  103.97 8.6375 110.95 8.7025 ;
      RECT  103.97 8.7025 110.95 21.02 ;
      RECT  110.95 8.6375 111.65 8.7025 ;
      RECT  111.65 8.6375 113.81 8.7025 ;
      RECT  111.65 8.7025 113.81 21.02 ;
      RECT  103.97 21.02 110.95 21.0525 ;
      RECT  111.65 21.02 113.81 21.0525 ;
      RECT  103.97 21.0525 110.95 21.7525 ;
      RECT  111.65 21.0525 113.81 21.7525 ;
      RECT  103.97 21.7525 110.95 21.8175 ;
      RECT  103.97 21.8175 110.95 41.9825 ;
      RECT  110.95 21.8175 111.65 41.9825 ;
      RECT  111.65 21.7525 113.81 21.8175 ;
      RECT  111.65 21.8175 113.81 41.9825 ;
      RECT  14.775 2.8525 19.7825 4.7775 ;
      RECT  14.775 4.7775 19.7825 4.845 ;
      RECT  19.7825 2.8525 20.4825 4.7775 ;
      RECT  20.4825 2.8525 21.445 4.7775 ;
      RECT  20.4825 4.7775 21.445 4.845 ;
      RECT  14.775 4.845 19.7825 8.6375 ;
      RECT  20.4825 4.845 21.445 8.6375 ;
      RECT  14.775 8.6375 19.7825 15.425 ;
      RECT  20.4825 8.6375 21.445 15.425 ;
      RECT  14.775 15.425 19.7825 15.4925 ;
      RECT  14.775 15.4925 19.7825 17.8825 ;
      RECT  19.7825 15.4925 20.4825 17.8825 ;
      RECT  20.4825 15.425 21.445 15.4925 ;
      RECT  20.4825 15.4925 21.445 17.8825 ;
      RECT  114.51 21.7525 122.835 54.77 ;
      RECT  114.51 54.77 122.835 54.8025 ;
      RECT  122.835 21.7525 123.535 54.77 ;
      RECT  123.535 21.7525 124.8975 54.77 ;
      RECT  123.535 54.77 124.8975 54.8025 ;
      RECT  120.04 54.8025 122.835 72.0925 ;
      RECT  123.535 54.8025 124.8975 72.0925 ;
      RECT  120.04 72.0925 122.835 77.7325 ;
      RECT  120.04 77.7325 122.835 77.765 ;
      RECT  122.835 77.7325 123.535 77.765 ;
      RECT  123.535 72.0925 124.8975 77.7325 ;
      RECT  123.535 77.7325 124.8975 77.765 ;
      RECT  101.68 8.6375 101.82 21.02 ;
      RECT  101.82 8.6375 102.38 21.02 ;
      RECT  101.82 21.02 102.38 21.0525 ;
      RECT  98.03 21.0525 101.12 21.7525 ;
      RECT  98.03 21.7525 101.12 41.9825 ;
      RECT  98.03 41.9825 101.12 55.0975 ;
      RECT  98.03 55.0975 101.12 69.5925 ;
      RECT  98.03 69.5925 101.12 69.625 ;
      RECT  98.03 69.625 101.12 69.6625 ;
      RECT  101.12 69.625 101.68 69.6625 ;
      RECT  96.95 18.3725 101.12 21.02 ;
      RECT  96.95 21.02 101.12 21.0525 ;
      RECT  101.12 18.3725 101.68 21.02 ;
   END
END    freepdk45_sram_1w1r_13x128
END    LIBRARY
